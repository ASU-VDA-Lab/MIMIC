module fake_ibex_1789_n_6916 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_974, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_854, n_1008, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_993, n_1012, n_689, n_960, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1004, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_6916);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_974;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_689;
input n_960;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1004;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_6916;

wire n_4557;
wire n_6873;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_6616;
wire n_6848;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_6744;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_6658;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_6842;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_6760;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_1070;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_6602;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_6562;
wire n_3979;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_4854;
wire n_6732;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6674;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_1078;
wire n_4422;
wire n_5743;
wire n_6868;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_1305;
wire n_2088;
wire n_6724;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_6638;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_6878;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_1424;
wire n_2625;
wire n_2444;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_6114;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_6864;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_1042;
wire n_5252;
wire n_6209;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_6824;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_6540;
wire n_4489;
wire n_6912;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2924;
wire n_2456;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_6802;
wire n_4725;
wire n_6691;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5969;
wire n_5920;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_6855;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6711;
wire n_6124;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_6136;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6128;
wire n_2361;
wire n_6804;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_6714;
wire n_4114;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_6857;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_6859;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_6379;
wire n_6911;
wire n_6766;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6893;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6850;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_6827;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_6699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_6901;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3477;
wire n_3070;
wire n_1575;
wire n_6773;
wire n_4416;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6765;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_6704;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_6727;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_6883;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_6652;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6915;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6731;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_6902;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_6837;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_6767;
wire n_4858;
wire n_6733;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_6723;
wire n_3339;
wire n_6900;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_1517;
wire n_5973;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_6856;
wire n_5770;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_6682;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_6777;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_6185;
wire n_6706;
wire n_5342;
wire n_6884;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_6745;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_1072;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_6881;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_6816;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_6712;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_6656;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_4919;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_6863;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_6805;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_6771;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_6695;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_6673;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_6910;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_6482;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_6483;
wire n_4686;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_6800;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4962;
wire n_1082;
wire n_4797;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_6897;
wire n_2982;
wire n_2634;
wire n_3124;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6847;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_6737;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_6780;
wire n_4309;
wire n_4027;
wire n_6758;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_6176;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_1033;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_6909;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6662;
wire n_6461;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_6823;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_6725;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_6914;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4970;
wire n_4652;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_6566;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_6808;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_6747;
wire n_3856;
wire n_6496;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_6787;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_6784;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_6741;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_5319;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5543;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_6807;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_6795;
wire n_6898;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_6785;
wire n_6738;
wire n_3030;
wire n_5631;
wire n_6818;
wire n_5983;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_6021;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_6899;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_6754;
wire n_4067;
wire n_6822;
wire n_6796;
wire n_6849;
wire n_6836;
wire n_4997;
wire n_5906;
wire n_6755;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_6476;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_6669;
wire n_5357;
wire n_6717;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_1709;
wire n_6655;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_6790;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_6840;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_6748;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6676;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_6448;
wire n_3684;
wire n_6667;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2573;
wire n_1793;
wire n_2424;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_6653;
wire n_3098;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5488;
wire n_3107;
wire n_5465;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_1053;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_6560;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_3614;
wire n_2888;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6701;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_2832;
wire n_4991;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_6907;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_6661;
wire n_6730;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_1775;
wire n_6889;
wire n_6361;
wire n_6803;
wire n_2570;
wire n_4025;
wire n_6751;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_6696;
wire n_2395;
wire n_6062;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3718;
wire n_3398;
wire n_6252;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_6726;
wire n_3238;
wire n_6740;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_6799;
wire n_2463;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_1251;
wire n_6657;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_6716;
wire n_6797;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_6694;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_6647;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_1067;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_6846;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_6398;
wire n_6700;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_6853;
wire n_1294;
wire n_1351;
wire n_6679;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_1830;
wire n_6770;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_6660;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_5096;
wire n_6480;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_6693;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_6819;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5869;
wire n_5862;
wire n_1238;
wire n_3959;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_3044;
wire n_3493;
wire n_2868;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_6860;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_6833;
wire n_2159;
wire n_6865;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_6794;
wire n_3637;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_5277;
wire n_5900;
wire n_3647;
wire n_6240;
wire n_3928;
wire n_3619;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_6498;
wire n_6720;
wire n_1669;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_6854;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_6832;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_6779;
wire n_2567;
wire n_5645;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_6887;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_6769;
wire n_6903;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_6861;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_6697;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_6826;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_6380;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_6703;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6719;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_3791;
wire n_6904;
wire n_6778;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_6444;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_6749;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_6692;
wire n_6590;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_6702;
wire n_3046;
wire n_6551;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_5644;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_6820;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_5324;
wire n_6547;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_6589;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5510;
wire n_5329;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_6879;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_6310;
wire n_6852;
wire n_5061;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_6249;
wire n_3559;
wire n_5184;
wire n_6440;
wire n_5747;
wire n_6575;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_6689;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_6643;
wire n_6569;
wire n_6814;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_5464;
wire n_6895;
wire n_6548;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_6890;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_6789;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_6867;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_6764;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_6772;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_3097;
wire n_2906;
wire n_5495;
wire n_6908;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_3822;
wire n_1276;
wire n_6874;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_6736;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_6025;
wire n_6168;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_6713;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_6750;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_6675;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_6828;
wire n_5123;
wire n_6160;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_6875;
wire n_1701;
wire n_5236;
wire n_6678;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_6870;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_6715;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_6140;
wire n_5903;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_6663;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_6844;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_6843;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_6877;
wire n_2821;
wire n_6892;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_6752;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_6698;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_1628;
wire n_6810;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1395;
wire n_1115;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_6049;
wire n_2419;
wire n_6671;
wire n_6791;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_6768;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6260;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_6906;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_6834;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_6812;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_4426;
wire n_3116;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_6001;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_6687;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_6762;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_6759;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_3960;
wire n_4007;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_4163;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_6886;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_1587;
wire n_2555;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_6710;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_6776;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_6905;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_1642;
wire n_5744;
wire n_6798;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_6665;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_6888;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_6677;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_6781;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_6811;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_6685;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_1060;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_6722;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6573;
wire n_6786;
wire n_6774;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_6851;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_6729;
wire n_6882;
wire n_1168;
wire n_5500;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6167;
wire n_6189;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_6721;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_6885;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_6806;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5984;
wire n_6385;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_6793;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_6746;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_6728;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_6858;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_6841;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_6896;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_6132;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6872;
wire n_6089;
wire n_5211;
wire n_1668;
wire n_5861;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3896;
wire n_3533;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6831;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_6690;
wire n_4650;
wire n_6415;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_6688;
wire n_2876;
wire n_6670;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_6680;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_6046;
wire n_1326;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_6705;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_6913;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_6355;
wire n_4755;
wire n_6329;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_6734;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_6825;
wire n_1036;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_6743;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_6809;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_6632;
wire n_2717;
wire n_1589;
wire n_5720;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_6654;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_6871;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_6672;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_5682;
wire n_6891;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1464;
wire n_1566;
wire n_6565;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6601;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_3331;
wire n_2999;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_6821;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_6775;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_6683;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6815;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5855;
wire n_5819;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_6763;
wire n_6782;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_6839;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_6515;
wire n_6619;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_6664;
wire n_5992;
wire n_5105;
wire n_6761;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_6894;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_6099;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_3747;
wire n_1323;
wire n_6753;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_5485;
wire n_5737;
wire n_6876;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_6829;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_6830;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_5306;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_6838;
wire n_2698;
wire n_6869;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_6735;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_6866;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_6742;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_6709;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_6756;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_6250;
wire n_6718;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_1167;
wire n_3231;
wire n_6423;
wire n_6659;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6668;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_6757;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_2345;
wire n_1139;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_6880;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_6686;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_1088;
wire n_6666;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_6708;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_6801;
wire n_1547;
wire n_1542;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_1131;
wire n_6707;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_6835;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_6792;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_1161;
wire n_1103;
wire n_6739;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_4147;
wire n_3992;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_2870;
wire n_6862;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_6783;
wire n_4738;
wire n_6604;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_6788;
wire n_2668;
wire n_6684;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_6817;
wire n_1661;
wire n_6261;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_1039;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_6845;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_6572;
wire n_4544;
wire n_4595;
wire n_4418;
wire n_2770;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_6813;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5594;
wire n_5335;
wire n_3417;
wire n_2725;
wire n_6681;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_109),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_364),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_919),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_506),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_442),
.Y(n_1026)
);

CKINVDCx16_ASAP7_75t_R g1027 ( 
.A(n_105),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_616),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_57),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_999),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_726),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_965),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_36),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_926),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_929),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_887),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_975),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_68),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_10),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_377),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_265),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_880),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_222),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_537),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_584),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_440),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_292),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_475),
.Y(n_1048)
);

BUFx10_ASAP7_75t_L g1049 ( 
.A(n_1001),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_769),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_319),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_155),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_663),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_870),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_689),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_123),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_197),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_875),
.Y(n_1058)
);

BUFx10_ASAP7_75t_L g1059 ( 
.A(n_827),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_191),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_151),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_961),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_102),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_991),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_265),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_878),
.Y(n_1066)
);

BUFx8_ASAP7_75t_SL g1067 ( 
.A(n_662),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_718),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_454),
.Y(n_1069)
);

BUFx8_ASAP7_75t_SL g1070 ( 
.A(n_11),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_695),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_388),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_557),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_835),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_552),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_883),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_39),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_875),
.Y(n_1078)
);

CKINVDCx14_ASAP7_75t_R g1079 ( 
.A(n_1000),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1013),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_27),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_179),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_433),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_709),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_694),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_470),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_129),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_261),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_808),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_304),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_739),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_269),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_963),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_720),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_79),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_460),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_115),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_801),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_187),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_285),
.Y(n_1100)
);

BUFx10_ASAP7_75t_L g1101 ( 
.A(n_977),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_939),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_617),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_547),
.Y(n_1104)
);

CKINVDCx16_ASAP7_75t_R g1105 ( 
.A(n_406),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_4),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_806),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_555),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_211),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_324),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_748),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_647),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_337),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_478),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_375),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_145),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_205),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_992),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_804),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_556),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_314),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_448),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_1017),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_630),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_1020),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_129),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_918),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_969),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_707),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_230),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_967),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_291),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_948),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_663),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_522),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_832),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_403),
.Y(n_1137)
);

BUFx10_ASAP7_75t_L g1138 ( 
.A(n_1003),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1007),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_904),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_38),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_481),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_988),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_885),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_518),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_877),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_654),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_637),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_39),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_604),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_934),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_532),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_597),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_236),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_743),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_623),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_504),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_266),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_898),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_256),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_971),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_243),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_316),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_930),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_720),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_749),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_487),
.Y(n_1167)
);

BUFx10_ASAP7_75t_L g1168 ( 
.A(n_15),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_97),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1021),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_71),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_256),
.Y(n_1172)
);

BUFx8_ASAP7_75t_SL g1173 ( 
.A(n_890),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_259),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1019),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_925),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_392),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_123),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_723),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_697),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_999),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_426),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_200),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_465),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_368),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_11),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_28),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_351),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_328),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_380),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_399),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_921),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_356),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_983),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_552),
.Y(n_1195)
);

CKINVDCx14_ASAP7_75t_R g1196 ( 
.A(n_979),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_968),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_154),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_993),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_826),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_587),
.Y(n_1201)
);

BUFx10_ASAP7_75t_L g1202 ( 
.A(n_554),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1002),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_346),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1014),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_281),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_967),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_509),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_917),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_673),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_392),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_258),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_138),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_955),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_111),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_55),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_783),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_532),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_268),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_972),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_118),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_964),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_998),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_521),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_49),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_144),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_738),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_236),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_170),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_633),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_122),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_876),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_266),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1002),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_514),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_621),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_611),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_349),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_908),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_986),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_189),
.Y(n_1241)
);

BUFx5_ASAP7_75t_L g1242 ( 
.A(n_430),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_890),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_451),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_709),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_524),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_38),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_350),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_306),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_555),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_391),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_84),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_658),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_611),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_994),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_36),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_345),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_604),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1015),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_401),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_803),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_55),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_16),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_672),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_275),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_123),
.Y(n_1266)
);

BUFx5_ASAP7_75t_L g1267 ( 
.A(n_51),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_34),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_698),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_112),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_441),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_108),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_723),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_913),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_715),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_429),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_989),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_996),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_570),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1013),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_599),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_956),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_907),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_506),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_978),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_868),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_349),
.Y(n_1287)
);

CKINVDCx16_ASAP7_75t_R g1288 ( 
.A(n_970),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_906),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_746),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_960),
.Y(n_1291)
);

BUFx5_ASAP7_75t_L g1292 ( 
.A(n_945),
.Y(n_1292)
);

BUFx10_ASAP7_75t_L g1293 ( 
.A(n_303),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_6),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_523),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1004),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_987),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_880),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_353),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_888),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_169),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1008),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_815),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_881),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_95),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_796),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_149),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_127),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_950),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_588),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1018),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_113),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_267),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_889),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1012),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_964),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_976),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_376),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_258),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_975),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_31),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_142),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1005),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_737),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_923),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_831),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_330),
.Y(n_1327)
);

INVxp67_ASAP7_75t_SL g1328 ( 
.A(n_203),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_689),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_828),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_952),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_669),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_457),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_19),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_751),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_497),
.Y(n_1336)
);

CKINVDCx14_ASAP7_75t_R g1337 ( 
.A(n_990),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_699),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_981),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_601),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_809),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_458),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_629),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_534),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_957),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_946),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_997),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_41),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_892),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_756),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_910),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_937),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1012),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_924),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1011),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_530),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_389),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_210),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_857),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_933),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1004),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_693),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_974),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_277),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1010),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_984),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_678),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_849),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_57),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_225),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_953),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_24),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_413),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_4),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_932),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_239),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_822),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_149),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_771),
.Y(n_1379)
);

BUFx10_ASAP7_75t_L g1380 ( 
.A(n_575),
.Y(n_1380)
);

BUFx10_ASAP7_75t_L g1381 ( 
.A(n_396),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_767),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_323),
.Y(n_1383)
);

BUFx2_ASAP7_75t_SL g1384 ( 
.A(n_938),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_132),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_61),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_584),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_356),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_762),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_445),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_966),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_333),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_947),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_664),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_468),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_99),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_474),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_643),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_895),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_985),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_887),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_555),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_242),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_771),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_733),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_282),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_845),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_14),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_973),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_228),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_940),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_556),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_731),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_240),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_436),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_144),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_958),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_175),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_600),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1016),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_320),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_253),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_936),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_711),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_196),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_316),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_588),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_568),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_86),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_696),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_688),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_889),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_703),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_934),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_150),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_920),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_419),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_275),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_956),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_982),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_170),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_892),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_863),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_255),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_951),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_433),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_626),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_884),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_288),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_905),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_85),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_65),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_337),
.Y(n_1453)
);

CKINVDCx6p67_ASAP7_75t_R g1454 ( 
.A(n_218),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_928),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_682),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_230),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_395),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_207),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_496),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_587),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_226),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_612),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_442),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_644),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_914),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_868),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_207),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_531),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_592),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_569),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_330),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_489),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_897),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_287),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_102),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_909),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_846),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_894),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_64),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_674),
.Y(n_1481)
);

BUFx5_ASAP7_75t_L g1482 ( 
.A(n_795),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_393),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_486),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_738),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_949),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_899),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_423),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_347),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_715),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_995),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_913),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_540),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_832),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_818),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_597),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_900),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_330),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_105),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_935),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_829),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_441),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_671),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_482),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_89),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_954),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_512),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_44),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_893),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_901),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_721),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_915),
.Y(n_1512)
);

CKINVDCx6p67_ASAP7_75t_R g1513 ( 
.A(n_988),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_499),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_251),
.Y(n_1515)
);

BUFx10_ASAP7_75t_L g1516 ( 
.A(n_342),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_313),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_891),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_783),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_711),
.Y(n_1520)
);

BUFx5_ASAP7_75t_L g1521 ( 
.A(n_625),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_930),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_108),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_63),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_914),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_886),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_358),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_620),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_882),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_159),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_874),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_45),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_162),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_580),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_888),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_650),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_460),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_428),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_903),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_959),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_306),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1006),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_635),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_269),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_768),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_652),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_292),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_403),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_81),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_710),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_639),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_451),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_911),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_486),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_579),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_896),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_807),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_925),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_854),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_24),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_500),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_789),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_574),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_249),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_139),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_433),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_919),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_759),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_457),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_922),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_152),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_845),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_253),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_289),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_830),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_509),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_833),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_160),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_879),
.Y(n_1579)
);

BUFx10_ASAP7_75t_L g1580 ( 
.A(n_102),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_822),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_943),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_298),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_10),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_654),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_195),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_457),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_584),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_384),
.Y(n_1589)
);

BUFx10_ASAP7_75t_L g1590 ( 
.A(n_218),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_462),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_422),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_143),
.Y(n_1593)
);

CKINVDCx16_ASAP7_75t_R g1594 ( 
.A(n_799),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_688),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_858),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_502),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_942),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_105),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_916),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_122),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_78),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_951),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_643),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_594),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1001),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_239),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_380),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_468),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_419),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1003),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_902),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_369),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_141),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_817),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_846),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_962),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_299),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_922),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_944),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_912),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_82),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1009),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_596),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_400),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_927),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_221),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_472),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_772),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_407),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_551),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_941),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_621),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_264),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_139),
.Y(n_1635)
);

BUFx10_ASAP7_75t_L g1636 ( 
.A(n_189),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_188),
.Y(n_1637)
);

BUFx8_ASAP7_75t_SL g1638 ( 
.A(n_638),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_51),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_571),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_901),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_246),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_785),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_112),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_636),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1014),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_542),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_273),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_646),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_413),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_765),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_980),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_346),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_287),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_931),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_621),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1349),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1615),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1349),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1172),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1191),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1228),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1231),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1269),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1270),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1454),
.Y(n_1666)
);

INVxp33_ASAP7_75t_SL g1667 ( 
.A(n_1423),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1224),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1306),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1319),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1340),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1292),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1358),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1427),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1067),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1511),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1656),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1067),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1260),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1268),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1350),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1023),
.Y(n_1682)
);

INVxp33_ASAP7_75t_SL g1683 ( 
.A(n_1620),
.Y(n_1683)
);

CKINVDCx16_ASAP7_75t_R g1684 ( 
.A(n_1027),
.Y(n_1684)
);

INVxp33_ASAP7_75t_L g1685 ( 
.A(n_1447),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1476),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1488),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1039),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1032),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1043),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1140),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1047),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1053),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1056),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1070),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1286),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1077),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1081),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1085),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1091),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1092),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1292),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1112),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1116),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1117),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1119),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1070),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1124),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1129),
.Y(n_1709)
);

INVxp33_ASAP7_75t_SL g1710 ( 
.A(n_1022),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1134),
.Y(n_1711)
);

INVxp33_ASAP7_75t_SL g1712 ( 
.A(n_1025),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1156),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1023),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1167),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1638),
.Y(n_1716)
);

CKINVDCx16_ASAP7_75t_R g1717 ( 
.A(n_1105),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1169),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1638),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1171),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1059),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1174),
.Y(n_1722)
);

CKINVDCx16_ASAP7_75t_R g1723 ( 
.A(n_1543),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1143),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1183),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1188),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1059),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1200),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1206),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1323),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1221),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1466),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1225),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1229),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1079),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1059),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1235),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1143),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1237),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1292),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1241),
.Y(n_1741)
);

INVxp67_ASAP7_75t_SL g1742 ( 
.A(n_1185),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1244),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1185),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1246),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1247),
.Y(n_1746)
);

INVxp33_ASAP7_75t_L g1747 ( 
.A(n_1173),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1249),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1292),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1250),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1079),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1251),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1337),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1261),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1337),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1049),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1196),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1140),
.Y(n_1758)
);

INVxp67_ASAP7_75t_SL g1759 ( 
.A(n_1246),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1271),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1272),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1120),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1279),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1292),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1287),
.Y(n_1765)
);

INVxp33_ASAP7_75t_SL g1766 ( 
.A(n_1026),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1301),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1303),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1312),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1292),
.Y(n_1770)
);

INVxp33_ASAP7_75t_SL g1771 ( 
.A(n_1029),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1324),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1140),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1335),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_1196),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1362),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1120),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1364),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1140),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1173),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1369),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1370),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1292),
.Y(n_1783)
);

CKINVDCx16_ASAP7_75t_R g1784 ( 
.A(n_1594),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1362),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1373),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1372),
.Y(n_1787)
);

BUFx2_ASAP7_75t_L g1788 ( 
.A(n_1373),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1120),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1374),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1691),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1724),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1735),
.Y(n_1793)
);

AND2x6_ASAP7_75t_L g1794 ( 
.A(n_1721),
.B(n_1515),
.Y(n_1794)
);

INVx2_ASAP7_75t_SL g1795 ( 
.A(n_1786),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1658),
.Y(n_1796)
);

INVx6_ASAP7_75t_L g1797 ( 
.A(n_1684),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1691),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1721),
.B(n_1242),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1788),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1685),
.B(n_1163),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1682),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1691),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1738),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1714),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1727),
.Y(n_1806)
);

BUFx8_ASAP7_75t_SL g1807 ( 
.A(n_1675),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1758),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1668),
.Y(n_1809)
);

BUFx8_ASAP7_75t_L g1810 ( 
.A(n_1687),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1742),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1667),
.A2(n_1253),
.B1(n_1258),
.B2(n_1075),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1758),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1744),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1678),
.Y(n_1815)
);

BUFx12f_ASAP7_75t_L g1816 ( 
.A(n_1695),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1657),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1727),
.B(n_1031),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1756),
.B(n_1443),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1717),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1723),
.A2(n_1253),
.B1(n_1258),
.B2(n_1075),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1660),
.B(n_1291),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1777),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1661),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1659),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1672),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1702),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1784),
.A2(n_1040),
.B1(n_1041),
.B2(n_1033),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1707),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1777),
.Y(n_1830)
);

OAI21x1_ASAP7_75t_L g1831 ( 
.A1(n_1740),
.A2(n_1046),
.B(n_1028),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1749),
.Y(n_1832)
);

BUFx8_ASAP7_75t_SL g1833 ( 
.A(n_1716),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1758),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1764),
.Y(n_1835)
);

INVx5_ASAP7_75t_L g1836 ( 
.A(n_1773),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1773),
.Y(n_1837)
);

INVx5_ASAP7_75t_L g1838 ( 
.A(n_1773),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1719),
.A2(n_1552),
.B1(n_1527),
.B2(n_1051),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1745),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1710),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1770),
.Y(n_1842)
);

BUFx12f_ASAP7_75t_L g1843 ( 
.A(n_1780),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1759),
.Y(n_1844)
);

INVx5_ASAP7_75t_L g1845 ( 
.A(n_1779),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1789),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1776),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1789),
.B(n_1736),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1779),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1779),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1762),
.B(n_1646),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1783),
.Y(n_1852)
);

INVxp33_ASAP7_75t_SL g1853 ( 
.A(n_1666),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1662),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1751),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1663),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1785),
.Y(n_1857)
);

INVx5_ASAP7_75t_L g1858 ( 
.A(n_1683),
.Y(n_1858)
);

INVx6_ASAP7_75t_L g1859 ( 
.A(n_1666),
.Y(n_1859)
);

INVx6_ASAP7_75t_L g1860 ( 
.A(n_1747),
.Y(n_1860)
);

AOI22x1_ASAP7_75t_SL g1861 ( 
.A1(n_1753),
.A2(n_1552),
.B1(n_1527),
.B2(n_1071),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1755),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1664),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1665),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1669),
.Y(n_1865)
);

AOI22x1_ASAP7_75t_SL g1866 ( 
.A1(n_1757),
.A2(n_1096),
.B1(n_1097),
.B2(n_1038),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1670),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1671),
.Y(n_1868)
);

BUFx12f_ASAP7_75t_L g1869 ( 
.A(n_1775),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1689),
.B(n_1163),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1677),
.B(n_1455),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1696),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1688),
.Y(n_1873)
);

OA21x2_ASAP7_75t_L g1874 ( 
.A1(n_1790),
.A2(n_1046),
.B(n_1028),
.Y(n_1874)
);

INVx4_ASAP7_75t_L g1875 ( 
.A(n_1673),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1674),
.Y(n_1876)
);

BUFx12f_ASAP7_75t_L g1877 ( 
.A(n_1712),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1676),
.Y(n_1878)
);

INVx5_ASAP7_75t_L g1879 ( 
.A(n_1730),
.Y(n_1879)
);

BUFx6f_ASAP7_75t_L g1880 ( 
.A(n_1690),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1766),
.B(n_1044),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1771),
.B(n_1045),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1679),
.Y(n_1883)
);

INVx5_ASAP7_75t_L g1884 ( 
.A(n_1732),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1692),
.Y(n_1885)
);

AOI22x1_ASAP7_75t_R g1886 ( 
.A1(n_1680),
.A2(n_1099),
.B1(n_1109),
.B2(n_1104),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1693),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1694),
.Y(n_1888)
);

INVx5_ASAP7_75t_L g1889 ( 
.A(n_1697),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1698),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1699),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1700),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1701),
.B(n_1048),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1703),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1704),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1705),
.Y(n_1896)
);

BUFx6f_ASAP7_75t_L g1897 ( 
.A(n_1706),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1708),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1709),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1711),
.Y(n_1900)
);

BUFx6f_ASAP7_75t_L g1901 ( 
.A(n_1713),
.Y(n_1901)
);

BUFx12f_ASAP7_75t_L g1902 ( 
.A(n_1681),
.Y(n_1902)
);

INVx4_ASAP7_75t_L g1903 ( 
.A(n_1686),
.Y(n_1903)
);

CKINVDCx6p67_ASAP7_75t_R g1904 ( 
.A(n_1715),
.Y(n_1904)
);

BUFx8_ASAP7_75t_L g1905 ( 
.A(n_1718),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1720),
.B(n_1050),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1722),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1725),
.B(n_1163),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1726),
.B(n_1052),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1728),
.Y(n_1910)
);

INVxp33_ASAP7_75t_SL g1911 ( 
.A(n_1729),
.Y(n_1911)
);

AND2x6_ASAP7_75t_L g1912 ( 
.A(n_1731),
.B(n_1515),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1733),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1734),
.B(n_1168),
.Y(n_1914)
);

INVx6_ASAP7_75t_L g1915 ( 
.A(n_1737),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1739),
.B(n_1513),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1741),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1743),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1746),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1748),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1750),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1752),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1754),
.Y(n_1923)
);

OAI21x1_ASAP7_75t_L g1924 ( 
.A1(n_1760),
.A2(n_1060),
.B(n_1057),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1761),
.Y(n_1925)
);

INVxp33_ASAP7_75t_SL g1926 ( 
.A(n_1763),
.Y(n_1926)
);

OA21x2_ASAP7_75t_L g1927 ( 
.A1(n_1765),
.A2(n_1060),
.B(n_1057),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1767),
.B(n_1242),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1768),
.B(n_1061),
.Y(n_1929)
);

OA21x2_ASAP7_75t_L g1930 ( 
.A1(n_1787),
.A2(n_1149),
.B(n_1111),
.Y(n_1930)
);

INVx5_ASAP7_75t_L g1931 ( 
.A(n_1769),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1772),
.B(n_1168),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1774),
.B(n_1455),
.Y(n_1933)
);

OA21x2_ASAP7_75t_L g1934 ( 
.A1(n_1782),
.A2(n_1149),
.B(n_1111),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1778),
.B(n_1063),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1781),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1658),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1691),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1724),
.Y(n_1939)
);

BUFx6f_ASAP7_75t_L g1940 ( 
.A(n_1691),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1691),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1786),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1724),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1786),
.B(n_1065),
.Y(n_1944)
);

BUFx12f_ASAP7_75t_L g1945 ( 
.A(n_1675),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1658),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1724),
.Y(n_1947)
);

XOR2xp5_ASAP7_75t_L g1948 ( 
.A(n_1675),
.B(n_1114),
.Y(n_1948)
);

OA21x2_ASAP7_75t_L g1949 ( 
.A1(n_1672),
.A2(n_1180),
.B(n_1157),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1786),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1735),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1675),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1691),
.Y(n_1953)
);

OA21x2_ASAP7_75t_L g1954 ( 
.A1(n_1672),
.A2(n_1180),
.B(n_1157),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1724),
.Y(n_1955)
);

INVx4_ASAP7_75t_L g1956 ( 
.A(n_1786),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1691),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1786),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1724),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1724),
.Y(n_1960)
);

OAI22x1_ASAP7_75t_L g1961 ( 
.A1(n_1675),
.A2(n_1069),
.B1(n_1072),
.B2(n_1068),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1786),
.Y(n_1962)
);

BUFx8_ASAP7_75t_L g1963 ( 
.A(n_1668),
.Y(n_1963)
);

CKINVDCx20_ASAP7_75t_R g1964 ( 
.A(n_1684),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1685),
.B(n_1168),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1724),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1724),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_L g1968 ( 
.A1(n_1672),
.A2(n_1318),
.B(n_1294),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1667),
.A2(n_1082),
.B1(n_1083),
.B2(n_1073),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1724),
.Y(n_1970)
);

NAND2x1p5_ASAP7_75t_L g1971 ( 
.A(n_1721),
.B(n_1517),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_SL g1972 ( 
.A(n_1721),
.B(n_1202),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1675),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1724),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1786),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1724),
.Y(n_1976)
);

OA21x2_ASAP7_75t_L g1977 ( 
.A1(n_1672),
.A2(n_1318),
.B(n_1294),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1685),
.B(n_1202),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1691),
.Y(n_1979)
);

INVx4_ASAP7_75t_L g1980 ( 
.A(n_1786),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1667),
.A2(n_1086),
.B1(n_1087),
.B2(n_1084),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1724),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1786),
.Y(n_1983)
);

OAI21x1_ASAP7_75t_L g1984 ( 
.A1(n_1672),
.A2(n_1405),
.B(n_1332),
.Y(n_1984)
);

BUFx2_ASAP7_75t_L g1985 ( 
.A(n_1735),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1735),
.B(n_1517),
.Y(n_1986)
);

CKINVDCx20_ASAP7_75t_R g1987 ( 
.A(n_1684),
.Y(n_1987)
);

INVx5_ASAP7_75t_L g1988 ( 
.A(n_1756),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1685),
.B(n_1202),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1735),
.B(n_1076),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1735),
.B(n_1076),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1724),
.Y(n_1992)
);

BUFx3_ASAP7_75t_L g1993 ( 
.A(n_1786),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1735),
.B(n_1199),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1724),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1691),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1691),
.Y(n_1997)
);

AOI22x1_ASAP7_75t_SL g1998 ( 
.A1(n_1675),
.A2(n_1154),
.B1(n_1394),
.B2(n_1330),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1724),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1786),
.B(n_1088),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1691),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1786),
.B(n_1089),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1685),
.B(n_1215),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1724),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1735),
.B(n_1199),
.Y(n_2005)
);

INVx4_ASAP7_75t_L g2006 ( 
.A(n_1786),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1786),
.Y(n_2007)
);

INVx3_ASAP7_75t_L g2008 ( 
.A(n_1724),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1735),
.B(n_1223),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1685),
.A2(n_1094),
.B1(n_1095),
.B2(n_1090),
.Y(n_2010)
);

CKINVDCx20_ASAP7_75t_R g2011 ( 
.A(n_1684),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1691),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1691),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1685),
.B(n_1215),
.Y(n_2014)
);

INVxp67_ASAP7_75t_L g2015 ( 
.A(n_1658),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1724),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1685),
.B(n_1215),
.Y(n_2017)
);

INVxp33_ASAP7_75t_SL g2018 ( 
.A(n_1721),
.Y(n_2018)
);

BUFx6f_ASAP7_75t_L g2019 ( 
.A(n_1691),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1786),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1924),
.Y(n_2021)
);

BUFx2_ASAP7_75t_L g2022 ( 
.A(n_1904),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1873),
.B(n_1431),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1904),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1911),
.B(n_1288),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1859),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1908),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1924),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1908),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1914),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1874),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1873),
.B(n_1508),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1831),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1923),
.B(n_1910),
.Y(n_2034)
);

CKINVDCx8_ASAP7_75t_R g2035 ( 
.A(n_1820),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1914),
.Y(n_2036)
);

BUFx8_ASAP7_75t_L g2037 ( 
.A(n_1877),
.Y(n_2037)
);

INVxp33_ASAP7_75t_SL g2038 ( 
.A(n_1841),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_2018),
.Y(n_2039)
);

OA21x2_ASAP7_75t_L g2040 ( 
.A1(n_1831),
.A2(n_1395),
.B(n_1386),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1923),
.B(n_1242),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1927),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2015),
.B(n_1293),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1854),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1864),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1930),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1934),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1968),
.Y(n_2048)
);

INVx3_ASAP7_75t_L g2049 ( 
.A(n_1864),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1846),
.B(n_1328),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1867),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1921),
.B(n_1242),
.Y(n_2052)
);

INVx4_ASAP7_75t_L g2053 ( 
.A(n_1830),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1949),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1856),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1954),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1977),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1898),
.B(n_1242),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1968),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1867),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1878),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1926),
.B(n_1293),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1863),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1801),
.B(n_1293),
.Y(n_2064)
);

CKINVDCx16_ASAP7_75t_R g2065 ( 
.A(n_1972),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1984),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1796),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1984),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1880),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1868),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1880),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1890),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1900),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1865),
.Y(n_2074)
);

INVx5_ASAP7_75t_L g2075 ( 
.A(n_1912),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1876),
.Y(n_2076)
);

BUFx8_ASAP7_75t_L g2077 ( 
.A(n_1816),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1932),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1937),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1993),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1817),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1890),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1825),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1848),
.B(n_1098),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1891),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1891),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_1946),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1892),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_1853),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1801),
.B(n_1380),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1893),
.B(n_1242),
.Y(n_2091)
);

NAND2xp33_ASAP7_75t_L g2092 ( 
.A(n_1912),
.B(n_1242),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1846),
.B(n_1343),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1806),
.B(n_1035),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1906),
.B(n_1267),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1909),
.B(n_1267),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_1912),
.Y(n_2097)
);

AND2x4_ASAP7_75t_L g2098 ( 
.A(n_1823),
.B(n_1036),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_1804),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1892),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1988),
.B(n_1054),
.Y(n_2101)
);

NAND2x1_ASAP7_75t_L g2102 ( 
.A(n_1794),
.B(n_1332),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1894),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1894),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1897),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1897),
.Y(n_2106)
);

INVx6_ASAP7_75t_L g2107 ( 
.A(n_1860),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1901),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_1965),
.B(n_1380),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1971),
.B(n_1818),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1901),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1907),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_SL g2113 ( 
.A(n_1965),
.B(n_1380),
.Y(n_2113)
);

HB1xp67_ASAP7_75t_L g2114 ( 
.A(n_1809),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1907),
.Y(n_2115)
);

BUFx2_ASAP7_75t_L g2116 ( 
.A(n_1872),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1919),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1919),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1792),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1929),
.B(n_1267),
.Y(n_2120)
);

INVx3_ASAP7_75t_L g2121 ( 
.A(n_1947),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1939),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1943),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1807),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1794),
.Y(n_2125)
);

AND2x4_ASAP7_75t_L g2126 ( 
.A(n_1988),
.B(n_1058),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1935),
.B(n_1267),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1915),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1933),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1802),
.B(n_1267),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1955),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1805),
.B(n_1267),
.Y(n_2132)
);

NAND2xp33_ASAP7_75t_SL g2133 ( 
.A(n_1978),
.B(n_1100),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1811),
.Y(n_2134)
);

CKINVDCx8_ASAP7_75t_R g2135 ( 
.A(n_1815),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1959),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1814),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_1978),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1840),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1844),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1794),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1847),
.Y(n_2142)
);

BUFx3_ASAP7_75t_L g2143 ( 
.A(n_1797),
.Y(n_2143)
);

CKINVDCx16_ASAP7_75t_R g2144 ( 
.A(n_1964),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1960),
.Y(n_2145)
);

INVx3_ASAP7_75t_L g2146 ( 
.A(n_1966),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1857),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1967),
.Y(n_2148)
);

BUFx6f_ASAP7_75t_L g2149 ( 
.A(n_1974),
.Y(n_2149)
);

NAND2xp33_ASAP7_75t_L g2150 ( 
.A(n_2003),
.B(n_1267),
.Y(n_2150)
);

AND2x4_ASAP7_75t_L g2151 ( 
.A(n_1986),
.B(n_1074),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2003),
.B(n_1078),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_2008),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1824),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1895),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_1903),
.B(n_1103),
.Y(n_2156)
);

CKINVDCx20_ASAP7_75t_R g2157 ( 
.A(n_1810),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1899),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2017),
.B(n_1482),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1970),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1913),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2017),
.B(n_1482),
.Y(n_2162)
);

INVx6_ASAP7_75t_L g2163 ( 
.A(n_1902),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1918),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1920),
.Y(n_2165)
);

BUFx8_ASAP7_75t_L g2166 ( 
.A(n_1945),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1989),
.B(n_1381),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1936),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2014),
.B(n_1381),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1885),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_1851),
.B(n_1080),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1887),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1888),
.B(n_1482),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1896),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1917),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1976),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1922),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1793),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1925),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1982),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1992),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1995),
.Y(n_2182)
);

INVx3_ASAP7_75t_L g2183 ( 
.A(n_1875),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_1883),
.B(n_1870),
.Y(n_2184)
);

INVx4_ASAP7_75t_L g2185 ( 
.A(n_1858),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1999),
.Y(n_2186)
);

INVx4_ASAP7_75t_L g2187 ( 
.A(n_1858),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2004),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_1819),
.B(n_1102),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2016),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1871),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1889),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1889),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1944),
.B(n_1482),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2000),
.B(n_2002),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1951),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1852),
.Y(n_2197)
);

AND2x6_ASAP7_75t_L g2198 ( 
.A(n_1916),
.B(n_1405),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1931),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1852),
.Y(n_2200)
);

INVxp67_ASAP7_75t_L g2201 ( 
.A(n_1963),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1985),
.B(n_1381),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1826),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1931),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1827),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1832),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1990),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1991),
.Y(n_2208)
);

BUFx2_ASAP7_75t_L g2209 ( 
.A(n_1956),
.Y(n_2209)
);

INVxp67_ASAP7_75t_L g2210 ( 
.A(n_1881),
.Y(n_2210)
);

BUFx3_ASAP7_75t_L g2211 ( 
.A(n_1869),
.Y(n_2211)
);

INVx3_ASAP7_75t_L g2212 ( 
.A(n_1980),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1994),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1795),
.B(n_1482),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2005),
.Y(n_2215)
);

BUFx3_ASAP7_75t_L g2216 ( 
.A(n_1843),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2009),
.Y(n_2217)
);

INVx3_ASAP7_75t_L g2218 ( 
.A(n_2006),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1795),
.B(n_1482),
.Y(n_2219)
);

BUFx6f_ASAP7_75t_L g2220 ( 
.A(n_1855),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1882),
.B(n_1482),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_1800),
.B(n_1106),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1822),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1905),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1969),
.B(n_1516),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1862),
.Y(n_2226)
);

CKINVDCx5p33_ASAP7_75t_R g2227 ( 
.A(n_1833),
.Y(n_2227)
);

BUFx3_ASAP7_75t_L g2228 ( 
.A(n_1829),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1942),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1950),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1879),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1958),
.Y(n_2232)
);

INVx3_ASAP7_75t_L g2233 ( 
.A(n_1879),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_1987),
.Y(n_2234)
);

INVx5_ASAP7_75t_L g2235 ( 
.A(n_1791),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_L g2236 ( 
.A(n_1962),
.B(n_1107),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_2011),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1975),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1983),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1835),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2007),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2020),
.Y(n_2242)
);

XNOR2x2_ASAP7_75t_R g2243 ( 
.A(n_1948),
.B(n_0),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1842),
.Y(n_2244)
);

NOR2x1_ASAP7_75t_L g2245 ( 
.A(n_2010),
.B(n_1398),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_1884),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1799),
.B(n_1521),
.Y(n_2247)
);

INVx3_ASAP7_75t_L g2248 ( 
.A(n_1884),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1928),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1836),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1981),
.B(n_1521),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_1828),
.A2(n_1110),
.B1(n_1113),
.B2(n_1108),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1791),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_1952),
.B(n_1128),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1961),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1961),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1836),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1838),
.Y(n_2258)
);

OA21x2_ASAP7_75t_L g2259 ( 
.A1(n_1812),
.A2(n_1413),
.B(n_1412),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_1798),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_1973),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1838),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_1839),
.B(n_1516),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1845),
.Y(n_2264)
);

INVx3_ASAP7_75t_L g2265 ( 
.A(n_1845),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1798),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1803),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1803),
.Y(n_2268)
);

CKINVDCx11_ASAP7_75t_R g2269 ( 
.A(n_1886),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1808),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_1808),
.B(n_1131),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1813),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1821),
.B(n_1516),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1813),
.Y(n_2274)
);

XNOR2xp5_ASAP7_75t_L g2275 ( 
.A(n_1861),
.B(n_1402),
.Y(n_2275)
);

NOR2x1_ASAP7_75t_L g2276 ( 
.A(n_1834),
.B(n_1421),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1834),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1837),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1837),
.Y(n_2279)
);

INVx5_ASAP7_75t_L g2280 ( 
.A(n_1849),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_1849),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1850),
.B(n_1521),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2019),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1850),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_1866),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1938),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2019),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1938),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1940),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2013),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1940),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1941),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_1941),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1953),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_1953),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1957),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1957),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2013),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1979),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1979),
.Y(n_2300)
);

BUFx6f_ASAP7_75t_L g2301 ( 
.A(n_1996),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1996),
.Y(n_2302)
);

INVxp67_ASAP7_75t_SL g2303 ( 
.A(n_1997),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_1998),
.B(n_1580),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_1997),
.B(n_1580),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2001),
.B(n_1521),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2001),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2012),
.B(n_1580),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2012),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2015),
.B(n_1590),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_1859),
.Y(n_2311)
);

BUFx3_ASAP7_75t_L g2312 ( 
.A(n_1859),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_1904),
.Y(n_2313)
);

INVx3_ASAP7_75t_L g2314 ( 
.A(n_1859),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1904),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_1908),
.B(n_1181),
.Y(n_2316)
);

INVx3_ASAP7_75t_L g2317 ( 
.A(n_1859),
.Y(n_2317)
);

BUFx6f_ASAP7_75t_L g2318 ( 
.A(n_1904),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1873),
.B(n_1521),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1873),
.B(n_1521),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_2018),
.Y(n_2321)
);

BUFx3_ASAP7_75t_L g2322 ( 
.A(n_1859),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1904),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_1859),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1924),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1904),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2015),
.B(n_1590),
.Y(n_2327)
);

AO22x2_ASAP7_75t_L g2328 ( 
.A1(n_2053),
.A2(n_1384),
.B1(n_1152),
.B2(n_1198),
.Y(n_2328)
);

BUFx4f_ASAP7_75t_L g2329 ( 
.A(n_2313),
.Y(n_2329)
);

BUFx3_ASAP7_75t_L g2330 ( 
.A(n_2037),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2174),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2195),
.B(n_1115),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2174),
.Y(n_2333)
);

BUFx3_ASAP7_75t_L g2334 ( 
.A(n_2037),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2316),
.B(n_1121),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2027),
.Y(n_2336)
);

INVx3_ASAP7_75t_L g2337 ( 
.A(n_2313),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2029),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2030),
.Y(n_2339)
);

INVx2_ASAP7_75t_SL g2340 ( 
.A(n_2178),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2036),
.Y(n_2341)
);

NAND2xp33_ASAP7_75t_SL g2342 ( 
.A(n_2318),
.B(n_1410),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2031),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_2318),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2042),
.Y(n_2345)
);

INVxp67_ASAP7_75t_SL g2346 ( 
.A(n_2067),
.Y(n_2346)
);

AOI22xp33_ASAP7_75t_L g2347 ( 
.A1(n_2245),
.A2(n_1636),
.B1(n_1590),
.B2(n_1438),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2316),
.B(n_1122),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2046),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2047),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2054),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2134),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2056),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2137),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2057),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2021),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2028),
.Y(n_2357)
);

INVxp33_ASAP7_75t_L g2358 ( 
.A(n_2079),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2087),
.B(n_1419),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2325),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2170),
.Y(n_2361)
);

OAI22xp5_ASAP7_75t_L g2362 ( 
.A1(n_2078),
.A2(n_1461),
.B1(n_1470),
.B2(n_1444),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_2033),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2172),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2077),
.Y(n_2365)
);

AO22x2_ASAP7_75t_L g2366 ( 
.A1(n_2255),
.A2(n_1179),
.B1(n_1264),
.B2(n_1233),
.Y(n_2366)
);

AOI22xp33_ASAP7_75t_L g2367 ( 
.A1(n_2223),
.A2(n_1636),
.B1(n_1485),
.B2(n_1514),
.Y(n_2367)
);

INVxp67_ASAP7_75t_L g2368 ( 
.A(n_2114),
.Y(n_2368)
);

AND2x6_ASAP7_75t_L g2369 ( 
.A(n_2097),
.B(n_1425),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_2077),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_2113),
.B(n_1126),
.Y(n_2371)
);

AND2x6_ASAP7_75t_L g2372 ( 
.A(n_2097),
.B(n_2024),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2210),
.B(n_1130),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2139),
.Y(n_2374)
);

BUFx3_ASAP7_75t_L g2375 ( 
.A(n_2166),
.Y(n_2375)
);

AND3x2_ASAP7_75t_L g2376 ( 
.A(n_2201),
.B(n_1523),
.C(n_1483),
.Y(n_2376)
);

BUFx2_ASAP7_75t_L g2377 ( 
.A(n_2178),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2140),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2271),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2050),
.B(n_1132),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2271),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2119),
.Y(n_2382)
);

NAND3xp33_ASAP7_75t_L g2383 ( 
.A(n_2025),
.B(n_1136),
.C(n_1135),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2122),
.Y(n_2384)
);

INVx5_ASAP7_75t_L g2385 ( 
.A(n_2022),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2050),
.B(n_1137),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2123),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2075),
.B(n_2022),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_2196),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2131),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_2033),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2142),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2147),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2136),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2145),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2175),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2148),
.Y(n_2397)
);

INVxp33_ASAP7_75t_L g2398 ( 
.A(n_2196),
.Y(n_2398)
);

INVx2_ASAP7_75t_SL g2399 ( 
.A(n_2312),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2177),
.Y(n_2400)
);

NAND2xp33_ASAP7_75t_L g2401 ( 
.A(n_2075),
.B(n_1521),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2093),
.B(n_1141),
.Y(n_2402)
);

BUFx6f_ASAP7_75t_L g2403 ( 
.A(n_2059),
.Y(n_2403)
);

AOI22x1_ASAP7_75t_L g2404 ( 
.A1(n_2066),
.A2(n_1449),
.B1(n_1471),
.B2(n_1425),
.Y(n_2404)
);

NAND3xp33_ASAP7_75t_L g2405 ( 
.A(n_2084),
.B(n_1145),
.C(n_1142),
.Y(n_2405)
);

INVx3_ASAP7_75t_L g2406 ( 
.A(n_2045),
.Y(n_2406)
);

NOR2x1p5_ASAP7_75t_L g2407 ( 
.A(n_2224),
.B(n_1147),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_2049),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2093),
.B(n_1148),
.Y(n_2409)
);

INVx3_ASAP7_75t_L g2410 ( 
.A(n_2051),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2160),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2176),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2179),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2155),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2173),
.Y(n_2415)
);

INVx3_ASAP7_75t_L g2416 ( 
.A(n_2060),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2158),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2064),
.B(n_1150),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_2138),
.B(n_1583),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2090),
.B(n_1153),
.Y(n_2420)
);

INVx1_ASAP7_75t_SL g2421 ( 
.A(n_2116),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_2157),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_2075),
.B(n_2315),
.Y(n_2423)
);

NAND3xp33_ASAP7_75t_L g2424 ( 
.A(n_2156),
.B(n_1158),
.C(n_1155),
.Y(n_2424)
);

INVx4_ASAP7_75t_L g2425 ( 
.A(n_2220),
.Y(n_2425)
);

OAI22xp33_ASAP7_75t_L g2426 ( 
.A1(n_2039),
.A2(n_1614),
.B1(n_1637),
.B2(n_1605),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2074),
.Y(n_2427)
);

AOI21x1_ASAP7_75t_L g2428 ( 
.A1(n_2048),
.A2(n_1428),
.B(n_1424),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2076),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2044),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2161),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2164),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2055),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2321),
.B(n_1636),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2165),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_2038),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2168),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2109),
.B(n_1160),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_2323),
.B(n_1162),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2023),
.B(n_1165),
.Y(n_2440)
);

OAI22xp33_ASAP7_75t_SL g2441 ( 
.A1(n_2065),
.A2(n_1177),
.B1(n_1178),
.B2(n_1166),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2032),
.B(n_1182),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2061),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2081),
.Y(n_2444)
);

AOI22xp33_ASAP7_75t_L g2445 ( 
.A1(n_2152),
.A2(n_1186),
.B1(n_1187),
.B2(n_1184),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2167),
.B(n_1189),
.Y(n_2446)
);

NAND3xp33_ASAP7_75t_L g2447 ( 
.A(n_2222),
.B(n_1193),
.C(n_1190),
.Y(n_2447)
);

AND3x2_ASAP7_75t_L g2448 ( 
.A(n_2285),
.B(n_2116),
.C(n_2243),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2083),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_2089),
.Y(n_2450)
);

INVx1_ASAP7_75t_SL g2451 ( 
.A(n_2322),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2130),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2132),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2068),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2043),
.B(n_1195),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_2166),
.Y(n_2456)
);

INVx2_ASAP7_75t_SL g2457 ( 
.A(n_2324),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2149),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2169),
.B(n_1201),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2310),
.B(n_2327),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2034),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2073),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2202),
.B(n_1049),
.Y(n_2463)
);

NOR2xp33_ASAP7_75t_L g2464 ( 
.A(n_2152),
.B(n_1204),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2048),
.Y(n_2465)
);

AOI22xp33_ASAP7_75t_L g2466 ( 
.A1(n_2259),
.A2(n_1211),
.B1(n_1212),
.B2(n_1210),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2229),
.Y(n_2467)
);

BUFx10_ASAP7_75t_L g2468 ( 
.A(n_2163),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2184),
.B(n_1213),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_2149),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_2102),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2230),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_2234),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_SL g2474 ( 
.A(n_2326),
.B(n_2125),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2203),
.Y(n_2475)
);

INVx2_ASAP7_75t_SL g2476 ( 
.A(n_2220),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_2059),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2205),
.Y(n_2478)
);

INVxp33_ASAP7_75t_L g2479 ( 
.A(n_2226),
.Y(n_2479)
);

INVx1_ASAP7_75t_SL g2480 ( 
.A(n_2209),
.Y(n_2480)
);

OR2x6_ASAP7_75t_L g2481 ( 
.A(n_2163),
.B(n_1223),
.Y(n_2481)
);

OR2x6_ASAP7_75t_L g2482 ( 
.A(n_2216),
.B(n_1311),
.Y(n_2482)
);

XOR2xp5_ASAP7_75t_L g2483 ( 
.A(n_2237),
.B(n_1066),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2159),
.B(n_1216),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2232),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2238),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2162),
.B(n_1217),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2094),
.B(n_1218),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2239),
.Y(n_2489)
);

INVx2_ASAP7_75t_SL g2490 ( 
.A(n_2226),
.Y(n_2490)
);

INVxp33_ASAP7_75t_L g2491 ( 
.A(n_2080),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2206),
.Y(n_2492)
);

NOR2x1p5_ASAP7_75t_L g2493 ( 
.A(n_2211),
.B(n_1219),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2240),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2094),
.B(n_1226),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2244),
.Y(n_2496)
);

AOI22xp5_ASAP7_75t_L g2497 ( 
.A1(n_2133),
.A2(n_1230),
.B1(n_1236),
.B2(n_1227),
.Y(n_2497)
);

BUFx2_ASAP7_75t_L g2498 ( 
.A(n_2209),
.Y(n_2498)
);

NAND2xp33_ASAP7_75t_L g2499 ( 
.A(n_2125),
.B(n_1238),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2141),
.B(n_2184),
.Y(n_2500)
);

AND2x2_ASAP7_75t_SL g2501 ( 
.A(n_2144),
.B(n_1192),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2040),
.Y(n_2502)
);

INVx2_ASAP7_75t_SL g2503 ( 
.A(n_2107),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2040),
.Y(n_2504)
);

INVxp67_ASAP7_75t_L g2505 ( 
.A(n_2080),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2180),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2124),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2098),
.B(n_1245),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2241),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2242),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2052),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2102),
.Y(n_2512)
);

INVxp67_ASAP7_75t_L g2513 ( 
.A(n_2098),
.Y(n_2513)
);

OR2x6_ASAP7_75t_L g2514 ( 
.A(n_2143),
.B(n_1311),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2062),
.B(n_1248),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2181),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2182),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2186),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2107),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2251),
.B(n_1252),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2214),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2188),
.Y(n_2522)
);

BUFx6f_ASAP7_75t_L g2523 ( 
.A(n_2260),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2225),
.B(n_1257),
.Y(n_2524)
);

INVx2_ASAP7_75t_SL g2525 ( 
.A(n_2026),
.Y(n_2525)
);

NAND3xp33_ASAP7_75t_L g2526 ( 
.A(n_2236),
.B(n_2252),
.C(n_2150),
.Y(n_2526)
);

INVx3_ASAP7_75t_L g2527 ( 
.A(n_2069),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2190),
.Y(n_2528)
);

BUFx3_ASAP7_75t_L g2529 ( 
.A(n_2035),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2071),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2072),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2082),
.Y(n_2532)
);

BUFx10_ASAP7_75t_L g2533 ( 
.A(n_2227),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2103),
.Y(n_2534)
);

CKINVDCx6p67_ASAP7_75t_R g2535 ( 
.A(n_2228),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2198),
.B(n_1262),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2105),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2101),
.B(n_1239),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_L g2539 ( 
.A(n_2185),
.B(n_1263),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2108),
.Y(n_2540)
);

INVx2_ASAP7_75t_SL g2541 ( 
.A(n_2311),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_2260),
.Y(n_2542)
);

INVx2_ASAP7_75t_SL g2543 ( 
.A(n_2314),
.Y(n_2543)
);

INVx2_ASAP7_75t_SL g2544 ( 
.A(n_2317),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2219),
.Y(n_2545)
);

INVx5_ASAP7_75t_L g2546 ( 
.A(n_2231),
.Y(n_2546)
);

BUFx8_ASAP7_75t_SL g2547 ( 
.A(n_2285),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2305),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2308),
.Y(n_2549)
);

OAI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2259),
.A2(n_2135),
.B1(n_2261),
.B2(n_2256),
.Y(n_2550)
);

BUFx2_ASAP7_75t_L g2551 ( 
.A(n_2254),
.Y(n_2551)
);

BUFx3_ASAP7_75t_L g2552 ( 
.A(n_2231),
.Y(n_2552)
);

BUFx2_ASAP7_75t_L g2553 ( 
.A(n_2254),
.Y(n_2553)
);

BUFx3_ASAP7_75t_L g2554 ( 
.A(n_2246),
.Y(n_2554)
);

AO21x2_ASAP7_75t_L g2555 ( 
.A1(n_2092),
.A2(n_1462),
.B(n_1460),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2111),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2058),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2063),
.Y(n_2558)
);

NOR3xp33_ASAP7_75t_L g2559 ( 
.A(n_2263),
.B(n_1383),
.C(n_1273),
.Y(n_2559)
);

INVx3_ASAP7_75t_L g2560 ( 
.A(n_2117),
.Y(n_2560)
);

OR2x2_ASAP7_75t_L g2561 ( 
.A(n_2273),
.B(n_1414),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2091),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2141),
.B(n_1265),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2101),
.B(n_1266),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2198),
.B(n_1275),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2095),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2070),
.Y(n_2567)
);

AND2x4_ASAP7_75t_L g2568 ( 
.A(n_2126),
.B(n_2183),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2198),
.B(n_1276),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2096),
.Y(n_2570)
);

INVx4_ASAP7_75t_L g2571 ( 
.A(n_2246),
.Y(n_2571)
);

XOR2xp5_ASAP7_75t_L g2572 ( 
.A(n_2275),
.B(n_2304),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2171),
.B(n_2189),
.Y(n_2573)
);

CKINVDCx6p67_ASAP7_75t_R g2574 ( 
.A(n_2269),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2129),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2085),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2086),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2265),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2088),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2120),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2151),
.A2(n_1284),
.B1(n_1290),
.B2(n_1281),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2127),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2187),
.B(n_2189),
.Y(n_2583)
);

BUFx6f_ASAP7_75t_L g2584 ( 
.A(n_2281),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2194),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2191),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2100),
.Y(n_2587)
);

INVxp33_ASAP7_75t_SL g2588 ( 
.A(n_2275),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2171),
.B(n_1295),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_SL g2590 ( 
.A(n_2126),
.B(n_1299),
.Y(n_2590)
);

NOR2x1p5_ASAP7_75t_L g2591 ( 
.A(n_2212),
.B(n_1305),
.Y(n_2591)
);

BUFx2_ASAP7_75t_L g2592 ( 
.A(n_2218),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2154),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2104),
.Y(n_2594)
);

AO21x2_ASAP7_75t_L g2595 ( 
.A1(n_2110),
.A2(n_1469),
.B(n_1465),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2207),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2233),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_SL g2598 ( 
.A(n_2221),
.B(n_1307),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2208),
.Y(n_2599)
);

INVx2_ASAP7_75t_SL g2600 ( 
.A(n_2151),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2213),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2106),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2112),
.Y(n_2603)
);

CKINVDCx5p33_ASAP7_75t_R g2604 ( 
.A(n_2248),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2215),
.Y(n_2605)
);

INVxp67_ASAP7_75t_SL g2606 ( 
.A(n_2099),
.Y(n_2606)
);

INVx3_ASAP7_75t_L g2607 ( 
.A(n_2115),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2118),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2250),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2121),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2217),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2282),
.Y(n_2612)
);

INVxp33_ASAP7_75t_L g2613 ( 
.A(n_2128),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2306),
.Y(n_2614)
);

INVx5_ASAP7_75t_L g2615 ( 
.A(n_2146),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2041),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2153),
.B(n_1308),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2276),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2319),
.Y(n_2619)
);

AND2x6_ASAP7_75t_L g2620 ( 
.A(n_2192),
.B(n_1449),
.Y(n_2620)
);

CKINVDCx16_ASAP7_75t_R g2621 ( 
.A(n_2193),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2320),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2199),
.Y(n_2623)
);

INVx2_ASAP7_75t_SL g2624 ( 
.A(n_2204),
.Y(n_2624)
);

BUFx6f_ASAP7_75t_L g2625 ( 
.A(n_2281),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2197),
.Y(n_2626)
);

NAND2xp33_ASAP7_75t_SL g2627 ( 
.A(n_2249),
.B(n_1346),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2247),
.B(n_1310),
.Y(n_2628)
);

INVxp67_ASAP7_75t_L g2629 ( 
.A(n_2258),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2257),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2264),
.Y(n_2631)
);

AO22x2_ASAP7_75t_L g2632 ( 
.A1(n_2262),
.A2(n_1550),
.B1(n_1622),
.B2(n_1468),
.Y(n_2632)
);

INVx3_ASAP7_75t_L g2633 ( 
.A(n_2235),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2200),
.Y(n_2634)
);

BUFx6f_ASAP7_75t_L g2635 ( 
.A(n_2293),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2235),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2235),
.Y(n_2637)
);

INVx3_ASAP7_75t_L g2638 ( 
.A(n_2280),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2280),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2280),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_2293),
.B(n_1313),
.Y(n_2641)
);

INVx1_ASAP7_75t_SL g2642 ( 
.A(n_2301),
.Y(n_2642)
);

OR2x6_ASAP7_75t_L g2643 ( 
.A(n_2301),
.B(n_1316),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2295),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2303),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2253),
.Y(n_2646)
);

BUFx3_ASAP7_75t_L g2647 ( 
.A(n_2253),
.Y(n_2647)
);

BUFx3_ASAP7_75t_L g2648 ( 
.A(n_2266),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2267),
.Y(n_2649)
);

BUFx3_ASAP7_75t_L g2650 ( 
.A(n_2270),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2272),
.B(n_1321),
.Y(n_2651)
);

INVx3_ASAP7_75t_L g2652 ( 
.A(n_2268),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2278),
.B(n_1322),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2279),
.B(n_1049),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2284),
.Y(n_2655)
);

OR2x2_ASAP7_75t_L g2656 ( 
.A(n_2286),
.B(n_1326),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2289),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_SL g2658 ( 
.A(n_2291),
.B(n_1327),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_2292),
.B(n_1329),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2294),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_SL g2661 ( 
.A(n_2299),
.B(n_1333),
.Y(n_2661)
);

INVx3_ASAP7_75t_L g2662 ( 
.A(n_2274),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2300),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2302),
.B(n_1334),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2309),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2277),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2283),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2287),
.Y(n_2668)
);

BUFx6f_ASAP7_75t_L g2669 ( 
.A(n_2288),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2290),
.B(n_1336),
.Y(n_2670)
);

INVx3_ASAP7_75t_L g2671 ( 
.A(n_2296),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2297),
.B(n_1338),
.Y(n_2672)
);

NAND3xp33_ASAP7_75t_L g2673 ( 
.A(n_2298),
.B(n_1342),
.C(n_1341),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2307),
.B(n_1344),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2031),
.Y(n_2675)
);

NAND2xp33_ASAP7_75t_R g2676 ( 
.A(n_2038),
.B(n_1348),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2174),
.Y(n_2677)
);

NAND2xp33_ASAP7_75t_L g2678 ( 
.A(n_2313),
.B(n_1356),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2174),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2031),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2031),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2031),
.Y(n_2682)
);

INVx3_ASAP7_75t_L g2683 ( 
.A(n_2313),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2031),
.Y(n_2684)
);

NOR2xp33_ASAP7_75t_L g2685 ( 
.A(n_2210),
.B(n_1357),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2031),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2174),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2174),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2031),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2031),
.Y(n_2690)
);

CKINVDCx6p67_ASAP7_75t_R g2691 ( 
.A(n_2216),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2031),
.Y(n_2692)
);

INVx4_ASAP7_75t_L g2693 ( 
.A(n_2313),
.Y(n_2693)
);

AND2x2_ASAP7_75t_SL g2694 ( 
.A(n_2022),
.B(n_1440),
.Y(n_2694)
);

INVxp67_ASAP7_75t_L g2695 ( 
.A(n_2067),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2031),
.Y(n_2696)
);

INVx1_ASAP7_75t_SL g2697 ( 
.A(n_2067),
.Y(n_2697)
);

INVx3_ASAP7_75t_L g2698 ( 
.A(n_2313),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2031),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2174),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2031),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2174),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_L g2703 ( 
.A(n_2210),
.B(n_1367),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_SL g2704 ( 
.A(n_2053),
.B(n_1376),
.Y(n_2704)
);

NAND2xp33_ASAP7_75t_L g2705 ( 
.A(n_2313),
.B(n_1377),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2031),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2195),
.B(n_1378),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2174),
.Y(n_2708)
);

BUFx2_ASAP7_75t_L g2709 ( 
.A(n_2053),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2195),
.B(n_1653),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2174),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2031),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2031),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2031),
.Y(n_2714)
);

INVxp33_ASAP7_75t_L g2715 ( 
.A(n_2067),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2031),
.Y(n_2716)
);

INVx2_ASAP7_75t_SL g2717 ( 
.A(n_2053),
.Y(n_2717)
);

INVx2_ASAP7_75t_SL g2718 ( 
.A(n_2053),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2031),
.Y(n_2719)
);

INVxp33_ASAP7_75t_L g2720 ( 
.A(n_2359),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2456),
.Y(n_2721)
);

AND2x4_ASAP7_75t_L g2722 ( 
.A(n_2385),
.B(n_1277),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2697),
.B(n_1101),
.Y(n_2723)
);

BUFx6f_ASAP7_75t_L g2724 ( 
.A(n_2523),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2346),
.B(n_1101),
.Y(n_2725)
);

INVx4_ASAP7_75t_L g2726 ( 
.A(n_2546),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2480),
.B(n_1101),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_SL g2728 ( 
.A(n_2695),
.B(n_1379),
.Y(n_2728)
);

NAND3x1_ASAP7_75t_L g2729 ( 
.A(n_2559),
.B(n_1596),
.C(n_1641),
.Y(n_2729)
);

OAI22xp33_ASAP7_75t_L g2730 ( 
.A1(n_2362),
.A2(n_1385),
.B1(n_1387),
.B2(n_1382),
.Y(n_2730)
);

BUFx3_ASAP7_75t_L g2731 ( 
.A(n_2330),
.Y(n_2731)
);

BUFx6f_ASAP7_75t_L g2732 ( 
.A(n_2523),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2465),
.Y(n_2733)
);

AO21x2_ASAP7_75t_L g2734 ( 
.A1(n_2502),
.A2(n_1480),
.B(n_1473),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2467),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2332),
.B(n_1388),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_SL g2737 ( 
.A(n_2368),
.B(n_1389),
.Y(n_2737)
);

BUFx3_ASAP7_75t_L g2738 ( 
.A(n_2334),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2687),
.Y(n_2739)
);

AND2x4_ASAP7_75t_L g2740 ( 
.A(n_2385),
.B(n_1282),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2687),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_SL g2742 ( 
.A(n_2358),
.B(n_2715),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2688),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2707),
.B(n_1138),
.Y(n_2744)
);

NAND2x1p5_ASAP7_75t_L g2745 ( 
.A(n_2329),
.B(n_1123),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2688),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2709),
.B(n_1390),
.Y(n_2747)
);

BUFx4f_ASAP7_75t_L g2748 ( 
.A(n_2691),
.Y(n_2748)
);

AO21x2_ASAP7_75t_L g2749 ( 
.A1(n_2502),
.A2(n_1484),
.B(n_1481),
.Y(n_2749)
);

BUFx8_ASAP7_75t_SL g2750 ( 
.A(n_2422),
.Y(n_2750)
);

AND2x4_ASAP7_75t_L g2751 ( 
.A(n_2385),
.B(n_1289),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_L g2752 ( 
.A(n_2460),
.B(n_1392),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2331),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2333),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2461),
.B(n_1302),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2677),
.Y(n_2756)
);

BUFx10_ASAP7_75t_L g2757 ( 
.A(n_2481),
.Y(n_2757)
);

INVx4_ASAP7_75t_SL g2758 ( 
.A(n_2365),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2679),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2700),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2702),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2708),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2711),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2343),
.Y(n_2764)
);

AND2x6_ASAP7_75t_L g2765 ( 
.A(n_2361),
.B(n_1055),
.Y(n_2765)
);

BUFx6f_ASAP7_75t_L g2766 ( 
.A(n_2523),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2710),
.B(n_1396),
.Y(n_2767)
);

CKINVDCx11_ASAP7_75t_R g2768 ( 
.A(n_2468),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2426),
.B(n_1397),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2361),
.Y(n_2770)
);

AOI22xp33_ASAP7_75t_SL g2771 ( 
.A1(n_2632),
.A2(n_1138),
.B1(n_1404),
.B2(n_1403),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2421),
.B(n_1406),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_2498),
.B(n_1408),
.Y(n_2773)
);

BUFx3_ASAP7_75t_L g2774 ( 
.A(n_2370),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2345),
.Y(n_2775)
);

NAND3x1_ASAP7_75t_L g2776 ( 
.A(n_2448),
.B(n_1655),
.C(n_1317),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2472),
.B(n_1415),
.Y(n_2777)
);

AND2x4_ASAP7_75t_L g2778 ( 
.A(n_2485),
.B(n_1314),
.Y(n_2778)
);

OAI22xp5_ASAP7_75t_L g2779 ( 
.A1(n_2562),
.A2(n_1418),
.B1(n_1422),
.B2(n_1416),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2364),
.Y(n_2780)
);

AND2x4_ASAP7_75t_L g2781 ( 
.A(n_2486),
.B(n_1339),
.Y(n_2781)
);

OAI22xp5_ASAP7_75t_SL g2782 ( 
.A1(n_2483),
.A2(n_1429),
.B1(n_1430),
.B2(n_1426),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2489),
.B(n_1433),
.Y(n_2783)
);

AND2x4_ASAP7_75t_L g2784 ( 
.A(n_2509),
.B(n_2510),
.Y(n_2784)
);

BUFx3_ASAP7_75t_L g2785 ( 
.A(n_2375),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2349),
.Y(n_2786)
);

NAND2x1p5_ASAP7_75t_L g2787 ( 
.A(n_2329),
.B(n_1298),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_2419),
.B(n_1435),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2352),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2481),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2685),
.B(n_2703),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2350),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2354),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2374),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2378),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2675),
.Y(n_2796)
);

BUFx6f_ASAP7_75t_L g2797 ( 
.A(n_2542),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2632),
.B(n_1138),
.Y(n_2798)
);

INVx8_ASAP7_75t_L g2799 ( 
.A(n_2546),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2542),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2524),
.B(n_1437),
.Y(n_2801)
);

AO22x2_ASAP7_75t_L g2802 ( 
.A1(n_2504),
.A2(n_1409),
.B1(n_1399),
.B2(n_1494),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2392),
.Y(n_2803)
);

AND2x4_ASAP7_75t_L g2804 ( 
.A(n_2717),
.B(n_1345),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2561),
.B(n_1441),
.Y(n_2805)
);

INVx3_ASAP7_75t_L g2806 ( 
.A(n_2542),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2643),
.Y(n_2807)
);

BUFx6f_ASAP7_75t_L g2808 ( 
.A(n_2584),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2680),
.Y(n_2809)
);

INVxp67_ASAP7_75t_SL g2810 ( 
.A(n_2584),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2364),
.B(n_1446),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_SL g2812 ( 
.A(n_2718),
.B(n_1451),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2584),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2681),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2463),
.B(n_1452),
.Y(n_2815)
);

AO22x2_ASAP7_75t_L g2816 ( 
.A1(n_2504),
.A2(n_1496),
.B1(n_1501),
.B2(n_1495),
.Y(n_2816)
);

NOR2x1p5_ASAP7_75t_L g2817 ( 
.A(n_2436),
.B(n_1453),
.Y(n_2817)
);

BUFx3_ASAP7_75t_L g2818 ( 
.A(n_2546),
.Y(n_2818)
);

NOR2xp33_ASAP7_75t_L g2819 ( 
.A(n_2551),
.B(n_1456),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2393),
.B(n_1457),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2682),
.Y(n_2821)
);

OAI221xp5_ASAP7_75t_L g2822 ( 
.A1(n_2367),
.A2(n_1463),
.B1(n_1464),
.B2(n_1459),
.C(n_1458),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2643),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2396),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2400),
.Y(n_2825)
);

AND2x4_ASAP7_75t_L g2826 ( 
.A(n_2591),
.B(n_1347),
.Y(n_2826)
);

INVx4_ASAP7_75t_SL g2827 ( 
.A(n_2529),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2625),
.Y(n_2828)
);

BUFx6f_ASAP7_75t_L g2829 ( 
.A(n_2625),
.Y(n_2829)
);

INVx3_ASAP7_75t_L g2830 ( 
.A(n_2625),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2694),
.B(n_1472),
.Y(n_2831)
);

NAND2x1p5_ASAP7_75t_L g2832 ( 
.A(n_2693),
.B(n_2425),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_L g2833 ( 
.A(n_2553),
.B(n_1475),
.Y(n_2833)
);

AND2x4_ASAP7_75t_L g2834 ( 
.A(n_2413),
.B(n_1354),
.Y(n_2834)
);

INVx1_ASAP7_75t_SL g2835 ( 
.A(n_2342),
.Y(n_2835)
);

AOI22xp5_ASAP7_75t_L g2836 ( 
.A1(n_2676),
.A2(n_1490),
.B1(n_1493),
.B2(n_1489),
.Y(n_2836)
);

AND2x4_ASAP7_75t_L g2837 ( 
.A(n_2427),
.B(n_1359),
.Y(n_2837)
);

BUFx6f_ASAP7_75t_L g2838 ( 
.A(n_2635),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2513),
.B(n_1498),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2429),
.Y(n_2840)
);

INVx2_ASAP7_75t_SL g2841 ( 
.A(n_2468),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2684),
.Y(n_2842)
);

BUFx3_ASAP7_75t_L g2843 ( 
.A(n_2535),
.Y(n_2843)
);

BUFx6f_ASAP7_75t_L g2844 ( 
.A(n_2635),
.Y(n_2844)
);

BUFx2_ASAP7_75t_L g2845 ( 
.A(n_2450),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2336),
.B(n_1499),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2338),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2686),
.Y(n_2848)
);

AOI22xp33_ASAP7_75t_L g2849 ( 
.A1(n_2627),
.A2(n_1504),
.B1(n_1505),
.B2(n_1502),
.Y(n_2849)
);

AOI22xp5_ASAP7_75t_L g2850 ( 
.A1(n_2455),
.A2(n_1532),
.B1(n_1533),
.B2(n_1528),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2689),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2690),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2339),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2341),
.B(n_1361),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2692),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2696),
.Y(n_2856)
);

NAND2x1p5_ASAP7_75t_L g2857 ( 
.A(n_2693),
.B(n_1055),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2430),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2407),
.Y(n_2859)
);

BUFx3_ASAP7_75t_L g2860 ( 
.A(n_2377),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2433),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_L g2862 ( 
.A(n_2573),
.B(n_1534),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2699),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2701),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2443),
.Y(n_2865)
);

INVx1_ASAP7_75t_SL g2866 ( 
.A(n_2451),
.Y(n_2866)
);

BUFx6f_ASAP7_75t_L g2867 ( 
.A(n_2635),
.Y(n_2867)
);

BUFx6f_ASAP7_75t_L g2868 ( 
.A(n_2363),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2444),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2414),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2373),
.B(n_1536),
.Y(n_2871)
);

BUFx3_ASAP7_75t_L g2872 ( 
.A(n_2425),
.Y(n_2872)
);

CKINVDCx5p33_ASAP7_75t_R g2873 ( 
.A(n_2507),
.Y(n_2873)
);

CKINVDCx11_ASAP7_75t_R g2874 ( 
.A(n_2533),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2417),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2431),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2432),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2706),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2466),
.B(n_1538),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_2383),
.B(n_1541),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_SL g2881 ( 
.A1(n_2328),
.A2(n_1546),
.B1(n_1547),
.B2(n_1545),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2600),
.B(n_1549),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2380),
.B(n_1554),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2452),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2386),
.B(n_1557),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2453),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2712),
.Y(n_2887)
);

AO21x2_ASAP7_75t_L g2888 ( 
.A1(n_2428),
.A2(n_1507),
.B(n_1503),
.Y(n_2888)
);

INVx3_ASAP7_75t_L g2889 ( 
.A(n_2337),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2328),
.B(n_1560),
.Y(n_2890)
);

CKINVDCx5p33_ASAP7_75t_R g2891 ( 
.A(n_2574),
.Y(n_2891)
);

NOR2x1p5_ASAP7_75t_L g2892 ( 
.A(n_2473),
.B(n_2337),
.Y(n_2892)
);

AND2x4_ASAP7_75t_L g2893 ( 
.A(n_2548),
.B(n_1365),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2415),
.Y(n_2894)
);

OR2x2_ASAP7_75t_L g2895 ( 
.A(n_2621),
.B(n_1561),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2562),
.A2(n_1564),
.B1(n_1565),
.B2(n_1563),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2713),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2415),
.Y(n_2898)
);

AO22x2_ASAP7_75t_L g2899 ( 
.A1(n_2526),
.A2(n_1524),
.B1(n_1530),
.B2(n_1519),
.Y(n_2899)
);

OR2x2_ASAP7_75t_L g2900 ( 
.A(n_2335),
.B(n_1566),
.Y(n_2900)
);

INVx2_ASAP7_75t_SL g2901 ( 
.A(n_2552),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_SL g2902 ( 
.A(n_2568),
.B(n_1569),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2549),
.B(n_1368),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2714),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2434),
.B(n_1573),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2716),
.Y(n_2906)
);

INVx3_ASAP7_75t_L g2907 ( 
.A(n_2344),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2719),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2351),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2353),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2564),
.B(n_1574),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2355),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2402),
.B(n_1575),
.Y(n_2913)
);

INVx4_ASAP7_75t_L g2914 ( 
.A(n_2344),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2435),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2356),
.Y(n_2916)
);

AND2x4_ASAP7_75t_L g2917 ( 
.A(n_2568),
.B(n_1375),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2464),
.B(n_1577),
.Y(n_2918)
);

AND2x4_ASAP7_75t_L g2919 ( 
.A(n_2340),
.B(n_1411),
.Y(n_2919)
);

NAND2x1p5_ASAP7_75t_L g2920 ( 
.A(n_2683),
.B(n_1055),
.Y(n_2920)
);

INVx4_ASAP7_75t_L g2921 ( 
.A(n_2683),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2357),
.Y(n_2922)
);

BUFx3_ASAP7_75t_L g2923 ( 
.A(n_2554),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2360),
.Y(n_2924)
);

AND2x4_ASAP7_75t_L g2925 ( 
.A(n_2389),
.B(n_1420),
.Y(n_2925)
);

AND2x2_ASAP7_75t_SL g2926 ( 
.A(n_2501),
.B(n_2678),
.Y(n_2926)
);

OR2x2_ASAP7_75t_L g2927 ( 
.A(n_2348),
.B(n_1578),
.Y(n_2927)
);

AND2x4_ASAP7_75t_L g2928 ( 
.A(n_2593),
.B(n_2476),
.Y(n_2928)
);

BUFx6f_ASAP7_75t_L g2929 ( 
.A(n_2363),
.Y(n_2929)
);

INVx8_ASAP7_75t_L g2930 ( 
.A(n_2482),
.Y(n_2930)
);

INVx3_ASAP7_75t_L g2931 ( 
.A(n_2698),
.Y(n_2931)
);

INVx4_ASAP7_75t_L g2932 ( 
.A(n_2698),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2437),
.Y(n_2933)
);

INVx1_ASAP7_75t_SL g2934 ( 
.A(n_2514),
.Y(n_2934)
);

BUFx3_ASAP7_75t_L g2935 ( 
.A(n_2533),
.Y(n_2935)
);

BUFx6f_ASAP7_75t_L g2936 ( 
.A(n_2363),
.Y(n_2936)
);

INVx4_ASAP7_75t_L g2937 ( 
.A(n_2571),
.Y(n_2937)
);

BUFx6f_ASAP7_75t_L g2938 ( 
.A(n_2391),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2449),
.Y(n_2939)
);

BUFx6f_ASAP7_75t_L g2940 ( 
.A(n_2391),
.Y(n_2940)
);

AO22x2_ASAP7_75t_L g2941 ( 
.A1(n_2366),
.A2(n_2371),
.B1(n_2550),
.B2(n_2538),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_SL g2942 ( 
.A(n_2497),
.B(n_1581),
.Y(n_2942)
);

HB1xp67_ASAP7_75t_L g2943 ( 
.A(n_2514),
.Y(n_2943)
);

AO22x2_ASAP7_75t_L g2944 ( 
.A1(n_2366),
.A2(n_1548),
.B1(n_1551),
.B2(n_1537),
.Y(n_2944)
);

NAND3xp33_ASAP7_75t_L g2945 ( 
.A(n_2405),
.B(n_1585),
.C(n_1584),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2596),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2454),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2506),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2445),
.B(n_1588),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2590),
.B(n_1592),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2409),
.B(n_1595),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2516),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2599),
.Y(n_2953)
);

BUFx6f_ASAP7_75t_L g2954 ( 
.A(n_2391),
.Y(n_2954)
);

AND2x4_ASAP7_75t_L g2955 ( 
.A(n_2490),
.B(n_1432),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2475),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2478),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2517),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2518),
.Y(n_2959)
);

AND2x4_ASAP7_75t_L g2960 ( 
.A(n_2462),
.B(n_1434),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2492),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2601),
.Y(n_2962)
);

AO21x2_ASAP7_75t_L g2963 ( 
.A1(n_2428),
.A2(n_1568),
.B(n_1562),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2522),
.Y(n_2964)
);

AO22x2_ASAP7_75t_L g2965 ( 
.A1(n_2538),
.A2(n_1576),
.B1(n_1586),
.B2(n_1571),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_L g2966 ( 
.A(n_2446),
.B(n_1597),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2567),
.B(n_1436),
.Y(n_2967)
);

INVx2_ASAP7_75t_SL g2968 ( 
.A(n_2482),
.Y(n_2968)
);

OAI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2488),
.A2(n_1602),
.B1(n_1607),
.B2(n_1599),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2440),
.B(n_1613),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2605),
.Y(n_2971)
);

AND2x4_ASAP7_75t_L g2972 ( 
.A(n_2571),
.B(n_1439),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2611),
.Y(n_2973)
);

BUFx6f_ASAP7_75t_L g2974 ( 
.A(n_2403),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_L g2975 ( 
.A(n_2459),
.B(n_1618),
.Y(n_2975)
);

BUFx3_ASAP7_75t_L g2976 ( 
.A(n_2399),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2539),
.B(n_1624),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2528),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2418),
.B(n_1628),
.Y(n_2979)
);

INVx5_ASAP7_75t_L g2980 ( 
.A(n_2369),
.Y(n_2980)
);

AND2x2_ASAP7_75t_L g2981 ( 
.A(n_2420),
.B(n_1631),
.Y(n_2981)
);

AND2x2_ASAP7_75t_SL g2982 ( 
.A(n_2705),
.B(n_1471),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_SL g2983 ( 
.A(n_2495),
.B(n_1634),
.Y(n_2983)
);

AND2x4_ASAP7_75t_L g2984 ( 
.A(n_2458),
.B(n_1448),
.Y(n_2984)
);

INVx4_ASAP7_75t_L g2985 ( 
.A(n_2369),
.Y(n_2985)
);

BUFx6f_ASAP7_75t_L g2986 ( 
.A(n_2403),
.Y(n_2986)
);

INVx5_ASAP7_75t_L g2987 ( 
.A(n_2369),
.Y(n_2987)
);

BUFx3_ASAP7_75t_L g2988 ( 
.A(n_2457),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2442),
.B(n_1635),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2494),
.Y(n_2990)
);

INVx4_ASAP7_75t_L g2991 ( 
.A(n_2369),
.Y(n_2991)
);

HB1xp67_ASAP7_75t_L g2992 ( 
.A(n_2479),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2438),
.B(n_1642),
.Y(n_2993)
);

AO22x2_ASAP7_75t_L g2994 ( 
.A1(n_2471),
.A2(n_1589),
.B1(n_1591),
.B2(n_1587),
.Y(n_2994)
);

AND2x6_ASAP7_75t_L g2995 ( 
.A(n_2511),
.B(n_1055),
.Y(n_2995)
);

NAND2x1p5_ASAP7_75t_L g2996 ( 
.A(n_2493),
.B(n_1208),
.Y(n_2996)
);

INVxp67_ASAP7_75t_L g2997 ( 
.A(n_2469),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2508),
.B(n_1647),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2496),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2566),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2347),
.B(n_1650),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2566),
.Y(n_3002)
);

INVx3_ASAP7_75t_L g3003 ( 
.A(n_2372),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2570),
.Y(n_3004)
);

NOR2xp33_ASAP7_75t_L g3005 ( 
.A(n_2589),
.B(n_1024),
.Y(n_3005)
);

INVx3_ASAP7_75t_L g3006 ( 
.A(n_2372),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2404),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2575),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2404),
.Y(n_3009)
);

INVx3_ASAP7_75t_L g3010 ( 
.A(n_2372),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2558),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2515),
.B(n_1030),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2586),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2583),
.B(n_1034),
.Y(n_3014)
);

CKINVDCx6p67_ASAP7_75t_R g3015 ( 
.A(n_2615),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2382),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2379),
.Y(n_3017)
);

AND2x4_ASAP7_75t_L g3018 ( 
.A(n_2458),
.B(n_1477),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2581),
.B(n_1593),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2398),
.B(n_2592),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2381),
.Y(n_3021)
);

OR2x6_ASAP7_75t_L g3022 ( 
.A(n_2503),
.B(n_1316),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2384),
.Y(n_3023)
);

BUFx6f_ASAP7_75t_L g3024 ( 
.A(n_2403),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2387),
.Y(n_3025)
);

BUFx6f_ASAP7_75t_L g3026 ( 
.A(n_2477),
.Y(n_3026)
);

NAND2x1p5_ASAP7_75t_L g3027 ( 
.A(n_2642),
.B(n_1208),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2390),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2394),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2395),
.Y(n_3030)
);

NAND3xp33_ASAP7_75t_L g3031 ( 
.A(n_2447),
.B(n_1254),
.C(n_1208),
.Y(n_3031)
);

OR2x2_ASAP7_75t_L g3032 ( 
.A(n_2617),
.B(n_1037),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2397),
.Y(n_3033)
);

CKINVDCx14_ASAP7_75t_R g3034 ( 
.A(n_2572),
.Y(n_3034)
);

CKINVDCx5p33_ASAP7_75t_R g3035 ( 
.A(n_2547),
.Y(n_3035)
);

AND2x6_ASAP7_75t_L g3036 ( 
.A(n_2570),
.B(n_1208),
.Y(n_3036)
);

AND2x4_ASAP7_75t_L g3037 ( 
.A(n_2470),
.B(n_1486),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2411),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2412),
.Y(n_3039)
);

INVx4_ASAP7_75t_L g3040 ( 
.A(n_2372),
.Y(n_3040)
);

NOR2xp33_ASAP7_75t_L g3041 ( 
.A(n_2704),
.B(n_1042),
.Y(n_3041)
);

AND2x4_ASAP7_75t_L g3042 ( 
.A(n_2470),
.B(n_1492),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_SL g3043 ( 
.A(n_2441),
.B(n_2536),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2484),
.B(n_1601),
.Y(n_3044)
);

INVx6_ASAP7_75t_L g3045 ( 
.A(n_2615),
.Y(n_3045)
);

NAND2x1p5_ASAP7_75t_L g3046 ( 
.A(n_2615),
.B(n_1254),
.Y(n_3046)
);

AOI22xp33_ASAP7_75t_L g3047 ( 
.A1(n_2585),
.A2(n_1064),
.B1(n_1093),
.B2(n_1062),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2519),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_2613),
.B(n_1118),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2656),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2595),
.Y(n_3051)
);

AO22x2_ASAP7_75t_L g3052 ( 
.A1(n_2471),
.A2(n_1608),
.B1(n_1609),
.B2(n_1604),
.Y(n_3052)
);

INVx3_ASAP7_75t_L g3053 ( 
.A(n_2633),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2576),
.Y(n_3054)
);

OR2x2_ASAP7_75t_L g3055 ( 
.A(n_2505),
.B(n_1125),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2487),
.B(n_1610),
.Y(n_3056)
);

INVx4_ASAP7_75t_SL g3057 ( 
.A(n_2620),
.Y(n_3057)
);

AND2x4_ASAP7_75t_L g3058 ( 
.A(n_2624),
.B(n_1500),
.Y(n_3058)
);

BUFx3_ASAP7_75t_L g3059 ( 
.A(n_2610),
.Y(n_3059)
);

BUFx4f_ASAP7_75t_L g3060 ( 
.A(n_2620),
.Y(n_3060)
);

BUFx6f_ASAP7_75t_L g3061 ( 
.A(n_2477),
.Y(n_3061)
);

AND2x6_ASAP7_75t_L g3062 ( 
.A(n_2521),
.B(n_2545),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2577),
.Y(n_3063)
);

NOR2xp33_ASAP7_75t_L g3064 ( 
.A(n_2439),
.B(n_1127),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2579),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2491),
.B(n_1133),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2670),
.Y(n_3067)
);

BUFx2_ASAP7_75t_L g3068 ( 
.A(n_2620),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2672),
.Y(n_3069)
);

BUFx6f_ASAP7_75t_L g3070 ( 
.A(n_2477),
.Y(n_3070)
);

NAND2x1p5_ASAP7_75t_L g3071 ( 
.A(n_2633),
.B(n_1254),
.Y(n_3071)
);

NAND2x1p5_ASAP7_75t_L g3072 ( 
.A(n_2638),
.B(n_1254),
.Y(n_3072)
);

BUFx3_ASAP7_75t_L g3073 ( 
.A(n_2597),
.Y(n_3073)
);

INVx2_ASAP7_75t_SL g3074 ( 
.A(n_2604),
.Y(n_3074)
);

INVx1_ASAP7_75t_SL g3075 ( 
.A(n_2620),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2565),
.B(n_1139),
.Y(n_3076)
);

INVx2_ASAP7_75t_SL g3077 ( 
.A(n_2376),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2630),
.Y(n_3078)
);

AND2x2_ASAP7_75t_SL g3079 ( 
.A(n_2499),
.B(n_1520),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2569),
.B(n_1144),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2587),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_2654),
.B(n_1146),
.Y(n_3082)
);

OA22x2_ASAP7_75t_L g3083 ( 
.A1(n_2631),
.A2(n_1159),
.B1(n_1161),
.B2(n_1151),
.Y(n_3083)
);

INVx3_ASAP7_75t_L g3084 ( 
.A(n_2638),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2424),
.B(n_1164),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_SL g3086 ( 
.A(n_2580),
.B(n_1170),
.Y(n_3086)
);

AO21x2_ASAP7_75t_L g3087 ( 
.A1(n_2555),
.A2(n_1629),
.B(n_1627),
.Y(n_3087)
);

AND2x6_ASAP7_75t_L g3088 ( 
.A(n_2582),
.B(n_1256),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2653),
.Y(n_3089)
);

AO22x2_ASAP7_75t_L g3090 ( 
.A1(n_2512),
.A2(n_2500),
.B1(n_2388),
.B2(n_2623),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_SL g3091 ( 
.A(n_2616),
.B(n_1632),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2664),
.Y(n_3092)
);

NOR2xp33_ASAP7_75t_L g3093 ( 
.A(n_2629),
.B(n_1175),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2557),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2520),
.B(n_2628),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2594),
.Y(n_3096)
);

INVx1_ASAP7_75t_SL g3097 ( 
.A(n_2609),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2606),
.B(n_2578),
.Y(n_3098)
);

INVx1_ASAP7_75t_SL g3099 ( 
.A(n_2609),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2602),
.Y(n_3100)
);

AND2x4_ASAP7_75t_L g3101 ( 
.A(n_2578),
.B(n_1518),
.Y(n_3101)
);

INVx3_ASAP7_75t_L g3102 ( 
.A(n_2648),
.Y(n_3102)
);

AND2x4_ASAP7_75t_L g3103 ( 
.A(n_2673),
.B(n_1525),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_SL g3104 ( 
.A(n_2619),
.B(n_2622),
.Y(n_3104)
);

AO22x2_ASAP7_75t_L g3105 ( 
.A1(n_2512),
.A2(n_1640),
.B1(n_1643),
.B2(n_1633),
.Y(n_3105)
);

INVx3_ASAP7_75t_L g3106 ( 
.A(n_2650),
.Y(n_3106)
);

CKINVDCx16_ASAP7_75t_R g3107 ( 
.A(n_2525),
.Y(n_3107)
);

HB1xp67_ASAP7_75t_L g3108 ( 
.A(n_2541),
.Y(n_3108)
);

AND2x2_ASAP7_75t_L g3109 ( 
.A(n_2543),
.B(n_1176),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2603),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2608),
.Y(n_3111)
);

OR2x2_ASAP7_75t_L g3112 ( 
.A(n_2544),
.B(n_1194),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2651),
.Y(n_3113)
);

AND2x4_ASAP7_75t_L g3114 ( 
.A(n_2563),
.B(n_2658),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2659),
.Y(n_3115)
);

BUFx6f_ASAP7_75t_L g3116 ( 
.A(n_2669),
.Y(n_3116)
);

AND2x4_ASAP7_75t_L g3117 ( 
.A(n_2661),
.B(n_1526),
.Y(n_3117)
);

INVx4_ASAP7_75t_L g3118 ( 
.A(n_2406),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2674),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2598),
.B(n_1644),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_SL g3121 ( 
.A(n_2647),
.B(n_1197),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2641),
.B(n_1203),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2657),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2660),
.Y(n_3124)
);

HB1xp67_ASAP7_75t_L g3125 ( 
.A(n_2645),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2665),
.Y(n_3126)
);

BUFx6f_ASAP7_75t_L g3127 ( 
.A(n_2669),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2406),
.Y(n_3128)
);

BUFx2_ASAP7_75t_L g3129 ( 
.A(n_2636),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2408),
.B(n_1645),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2646),
.Y(n_3131)
);

AO22x2_ASAP7_75t_L g3132 ( 
.A1(n_2474),
.A2(n_1651),
.B1(n_1648),
.B2(n_1542),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2408),
.B(n_1205),
.Y(n_3133)
);

AND2x4_ASAP7_75t_L g3134 ( 
.A(n_2423),
.B(n_1529),
.Y(n_3134)
);

AO22x2_ASAP7_75t_L g3135 ( 
.A1(n_2637),
.A2(n_1603),
.B1(n_1606),
.B2(n_1600),
.Y(n_3135)
);

AND2x6_ASAP7_75t_L g3136 ( 
.A(n_2639),
.B(n_1256),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2612),
.Y(n_3137)
);

INVx4_ASAP7_75t_L g3138 ( 
.A(n_2410),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2614),
.Y(n_3139)
);

BUFx3_ASAP7_75t_L g3140 ( 
.A(n_2640),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2530),
.Y(n_3141)
);

INVx4_ASAP7_75t_L g3142 ( 
.A(n_2410),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2618),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2416),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2531),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2416),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_2588),
.A2(n_1209),
.B1(n_1214),
.B2(n_1207),
.Y(n_3147)
);

INVx2_ASAP7_75t_SL g3148 ( 
.A(n_2644),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2532),
.Y(n_3149)
);

INVx1_ASAP7_75t_SL g3150 ( 
.A(n_2667),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2607),
.B(n_1220),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2607),
.B(n_1222),
.Y(n_3152)
);

INVx2_ASAP7_75t_SL g3153 ( 
.A(n_2649),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2655),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_2634),
.B(n_1232),
.Y(n_3155)
);

CKINVDCx16_ASAP7_75t_R g3156 ( 
.A(n_2668),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2537),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2663),
.Y(n_3158)
);

INVx3_ASAP7_75t_L g3159 ( 
.A(n_2527),
.Y(n_3159)
);

INVx4_ASAP7_75t_L g3160 ( 
.A(n_2669),
.Y(n_3160)
);

BUFx6f_ASAP7_75t_L g3161 ( 
.A(n_2527),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_2540),
.Y(n_3162)
);

BUFx6f_ASAP7_75t_L g3163 ( 
.A(n_2534),
.Y(n_3163)
);

NAND2x1p5_ASAP7_75t_L g3164 ( 
.A(n_2534),
.B(n_1256),
.Y(n_3164)
);

NAND2x1p5_ASAP7_75t_L g3165 ( 
.A(n_2560),
.B(n_1256),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2556),
.Y(n_3166)
);

CKINVDCx5p33_ASAP7_75t_R g3167 ( 
.A(n_2560),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2626),
.B(n_1234),
.Y(n_3168)
);

OAI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_2666),
.A2(n_1544),
.B1(n_1555),
.B2(n_1520),
.Y(n_3169)
);

AND2x6_ASAP7_75t_L g3170 ( 
.A(n_2652),
.B(n_1649),
.Y(n_3170)
);

AOI22xp5_ASAP7_75t_L g3171 ( 
.A1(n_2401),
.A2(n_1243),
.B1(n_1259),
.B2(n_1255),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_2652),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2662),
.Y(n_3173)
);

INVxp67_ASAP7_75t_L g3174 ( 
.A(n_2662),
.Y(n_3174)
);

BUFx3_ASAP7_75t_L g3175 ( 
.A(n_2671),
.Y(n_3175)
);

INVx4_ASAP7_75t_L g3176 ( 
.A(n_2671),
.Y(n_3176)
);

BUFx6f_ASAP7_75t_L g3177 ( 
.A(n_2523),
.Y(n_3177)
);

BUFx6f_ASAP7_75t_L g3178 ( 
.A(n_2523),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2465),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2697),
.B(n_1278),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2467),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2467),
.Y(n_3182)
);

AND2x4_ASAP7_75t_L g3183 ( 
.A(n_2385),
.B(n_1612),
.Y(n_3183)
);

AND2x4_ASAP7_75t_L g3184 ( 
.A(n_2385),
.B(n_1619),
.Y(n_3184)
);

BUFx6f_ASAP7_75t_L g3185 ( 
.A(n_2523),
.Y(n_3185)
);

BUFx3_ASAP7_75t_L g3186 ( 
.A(n_2330),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_2697),
.B(n_1280),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2467),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2467),
.Y(n_3189)
);

AOI22xp5_ASAP7_75t_L g3190 ( 
.A1(n_2359),
.A2(n_1285),
.B1(n_1296),
.B2(n_1283),
.Y(n_3190)
);

INVxp67_ASAP7_75t_SL g3191 ( 
.A(n_2695),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2467),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2467),
.Y(n_3193)
);

INVx1_ASAP7_75t_SL g3194 ( 
.A(n_2697),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2467),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2467),
.Y(n_3196)
);

INVx4_ASAP7_75t_L g3197 ( 
.A(n_2546),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_2697),
.B(n_1297),
.Y(n_3198)
);

INVx3_ASAP7_75t_L g3199 ( 
.A(n_2523),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2467),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_SL g3201 ( 
.A(n_2697),
.B(n_1300),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2467),
.Y(n_3202)
);

OAI22xp33_ASAP7_75t_SL g3203 ( 
.A1(n_2362),
.A2(n_1309),
.B1(n_1315),
.B2(n_1304),
.Y(n_3203)
);

AND2x4_ASAP7_75t_L g3204 ( 
.A(n_2385),
.B(n_1621),
.Y(n_3204)
);

AND3x4_ASAP7_75t_L g3205 ( 
.A(n_2330),
.B(n_1352),
.C(n_1320),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2465),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_2523),
.Y(n_3207)
);

AOI22xp33_ASAP7_75t_L g3208 ( 
.A1(n_2559),
.A2(n_1331),
.B1(n_1351),
.B2(n_1325),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2465),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2467),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2358),
.B(n_1353),
.Y(n_3211)
);

INVxp67_ASAP7_75t_SL g3212 ( 
.A(n_2695),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2467),
.Y(n_3213)
);

NAND2xp33_ASAP7_75t_R g3214 ( 
.A(n_2456),
.B(n_0),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_2697),
.B(n_1355),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2332),
.B(n_1360),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_SL g3217 ( 
.A(n_2697),
.B(n_1363),
.Y(n_3217)
);

INVx5_ASAP7_75t_L g3218 ( 
.A(n_2523),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2465),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2465),
.Y(n_3220)
);

AND2x6_ASAP7_75t_L g3221 ( 
.A(n_2687),
.B(n_1649),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2465),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2467),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_2358),
.B(n_1366),
.Y(n_3224)
);

AND2x4_ASAP7_75t_L g3225 ( 
.A(n_2385),
.B(n_1623),
.Y(n_3225)
);

INVx3_ASAP7_75t_L g3226 ( 
.A(n_2523),
.Y(n_3226)
);

BUFx6f_ASAP7_75t_L g3227 ( 
.A(n_2523),
.Y(n_3227)
);

AND2x2_ASAP7_75t_L g3228 ( 
.A(n_2697),
.B(n_1371),
.Y(n_3228)
);

AO22x2_ASAP7_75t_L g3229 ( 
.A1(n_2362),
.A2(n_1626),
.B1(n_1352),
.B2(n_1559),
.Y(n_3229)
);

BUFx6f_ASAP7_75t_L g3230 ( 
.A(n_2523),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2467),
.Y(n_3231)
);

INVxp67_ASAP7_75t_L g3232 ( 
.A(n_2697),
.Y(n_3232)
);

AND2x4_ASAP7_75t_L g3233 ( 
.A(n_2385),
.B(n_1320),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2467),
.Y(n_3234)
);

INVxp67_ASAP7_75t_SL g3235 ( 
.A(n_2695),
.Y(n_3235)
);

NAND3x1_ASAP7_75t_L g3236 ( 
.A(n_2559),
.B(n_0),
.C(n_1),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_2330),
.Y(n_3237)
);

AND2x2_ASAP7_75t_L g3238 ( 
.A(n_2697),
.B(n_1391),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2465),
.Y(n_3239)
);

INVx4_ASAP7_75t_L g3240 ( 
.A(n_2546),
.Y(n_3240)
);

CKINVDCx20_ASAP7_75t_R g3241 ( 
.A(n_2456),
.Y(n_3241)
);

AND2x6_ASAP7_75t_L g3242 ( 
.A(n_2687),
.B(n_1649),
.Y(n_3242)
);

BUFx6f_ASAP7_75t_L g3243 ( 
.A(n_2523),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2467),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2332),
.B(n_1393),
.Y(n_3245)
);

AND2x4_ASAP7_75t_L g3246 ( 
.A(n_2385),
.B(n_1559),
.Y(n_3246)
);

AND2x4_ASAP7_75t_L g3247 ( 
.A(n_2385),
.B(n_1611),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2467),
.Y(n_3248)
);

INVx3_ASAP7_75t_L g3249 ( 
.A(n_2523),
.Y(n_3249)
);

AND2x4_ASAP7_75t_L g3250 ( 
.A(n_2385),
.B(n_1611),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2467),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_2697),
.B(n_1400),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2697),
.B(n_1401),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_SL g3254 ( 
.A(n_2697),
.B(n_1598),
.Y(n_3254)
);

AO22x2_ASAP7_75t_L g3255 ( 
.A1(n_2362),
.A2(n_1652),
.B1(n_1616),
.B2(n_1555),
.Y(n_3255)
);

AND2x6_ASAP7_75t_L g3256 ( 
.A(n_2687),
.B(n_1649),
.Y(n_3256)
);

BUFx2_ASAP7_75t_L g3257 ( 
.A(n_2697),
.Y(n_3257)
);

INVx5_ASAP7_75t_L g3258 ( 
.A(n_2523),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2467),
.Y(n_3259)
);

OR2x6_ASAP7_75t_L g3260 ( 
.A(n_2330),
.B(n_1616),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2465),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2467),
.Y(n_3262)
);

AOI22xp5_ASAP7_75t_L g3263 ( 
.A1(n_2359),
.A2(n_1417),
.B1(n_1442),
.B2(n_1407),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2467),
.Y(n_3264)
);

CKINVDCx5p33_ASAP7_75t_R g3265 ( 
.A(n_2456),
.Y(n_3265)
);

AOI22xp5_ASAP7_75t_L g3266 ( 
.A1(n_2359),
.A2(n_1450),
.B1(n_1467),
.B2(n_1445),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_2465),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_2697),
.B(n_1474),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2687),
.Y(n_3269)
);

AND2x4_ASAP7_75t_L g3270 ( 
.A(n_2385),
.B(n_1652),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_2359),
.A2(n_1479),
.B1(n_1487),
.B2(n_1478),
.Y(n_3271)
);

CKINVDCx20_ASAP7_75t_R g3272 ( 
.A(n_2456),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2465),
.Y(n_3273)
);

OR2x6_ASAP7_75t_L g3274 ( 
.A(n_2330),
.B(n_1625),
.Y(n_3274)
);

NAND2x1p5_ASAP7_75t_L g3275 ( 
.A(n_2330),
.B(n_1654),
.Y(n_3275)
);

AND2x4_ASAP7_75t_L g3276 ( 
.A(n_2385),
.B(n_1639),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_2523),
.Y(n_3277)
);

BUFx6f_ASAP7_75t_L g3278 ( 
.A(n_2523),
.Y(n_3278)
);

BUFx3_ASAP7_75t_L g3279 ( 
.A(n_2330),
.Y(n_3279)
);

NOR2xp33_ASAP7_75t_SL g3280 ( 
.A(n_2456),
.B(n_1491),
.Y(n_3280)
);

NOR2xp33_ASAP7_75t_L g3281 ( 
.A(n_2358),
.B(n_1497),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_2332),
.B(n_1506),
.Y(n_3282)
);

INVx4_ASAP7_75t_L g3283 ( 
.A(n_2546),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2687),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2332),
.B(n_1509),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_L g3286 ( 
.A(n_2358),
.B(n_1510),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_SL g3287 ( 
.A(n_2697),
.B(n_1617),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2332),
.B(n_1512),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2465),
.Y(n_3289)
);

INVx3_ASAP7_75t_L g3290 ( 
.A(n_2523),
.Y(n_3290)
);

AND2x4_ASAP7_75t_L g3291 ( 
.A(n_2385),
.B(n_1630),
.Y(n_3291)
);

BUFx3_ASAP7_75t_L g3292 ( 
.A(n_2330),
.Y(n_3292)
);

INVx4_ASAP7_75t_L g3293 ( 
.A(n_2546),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2687),
.Y(n_3294)
);

BUFx6f_ASAP7_75t_L g3295 ( 
.A(n_2523),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2687),
.Y(n_3296)
);

AND2x2_ASAP7_75t_L g3297 ( 
.A(n_2697),
.B(n_1522),
.Y(n_3297)
);

NOR2xp33_ASAP7_75t_L g3298 ( 
.A(n_2358),
.B(n_1531),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_2465),
.Y(n_3299)
);

AND2x6_ASAP7_75t_L g3300 ( 
.A(n_2687),
.B(n_1654),
.Y(n_3300)
);

INVx4_ASAP7_75t_L g3301 ( 
.A(n_2546),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_2332),
.B(n_1535),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_2523),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2687),
.Y(n_3304)
);

AOI22xp33_ASAP7_75t_L g3305 ( 
.A1(n_2559),
.A2(n_1540),
.B1(n_1553),
.B2(n_1539),
.Y(n_3305)
);

AOI22xp5_ASAP7_75t_SL g3306 ( 
.A1(n_2483),
.A2(n_1558),
.B1(n_1567),
.B2(n_1556),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2687),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_2465),
.Y(n_3308)
);

INVx4_ASAP7_75t_L g3309 ( 
.A(n_2546),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_2697),
.B(n_1570),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_2687),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_2687),
.Y(n_3312)
);

OR2x2_ASAP7_75t_L g3313 ( 
.A(n_2362),
.B(n_1572),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2687),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_2465),
.Y(n_3315)
);

OR2x6_ASAP7_75t_L g3316 ( 
.A(n_2330),
.B(n_1544),
.Y(n_3316)
);

BUFx6f_ASAP7_75t_L g3317 ( 
.A(n_2523),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_2697),
.B(n_1579),
.Y(n_3318)
);

INVxp67_ASAP7_75t_L g3319 ( 
.A(n_2697),
.Y(n_3319)
);

INVx4_ASAP7_75t_L g3320 ( 
.A(n_2546),
.Y(n_3320)
);

INVx2_ASAP7_75t_SL g3321 ( 
.A(n_2468),
.Y(n_3321)
);

BUFx6f_ASAP7_75t_L g3322 ( 
.A(n_2523),
.Y(n_3322)
);

INVx4_ASAP7_75t_L g3323 ( 
.A(n_2546),
.Y(n_3323)
);

INVx3_ASAP7_75t_L g3324 ( 
.A(n_2523),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2687),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2687),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_L g3327 ( 
.A(n_2358),
.B(n_1582),
.Y(n_3327)
);

INVxp33_ASAP7_75t_L g3328 ( 
.A(n_2359),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_2358),
.B(n_1625),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_2697),
.B(n_1630),
.Y(n_3330)
);

NOR2xp33_ASAP7_75t_L g3331 ( 
.A(n_2358),
.B(n_1639),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2687),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2332),
.B(n_1),
.Y(n_3333)
);

BUFx2_ASAP7_75t_L g3334 ( 
.A(n_2697),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_2697),
.B(n_1),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2467),
.Y(n_3336)
);

BUFx8_ASAP7_75t_SL g3337 ( 
.A(n_2456),
.Y(n_3337)
);

AND2x4_ASAP7_75t_L g3338 ( 
.A(n_2385),
.B(n_2),
.Y(n_3338)
);

INVx3_ASAP7_75t_L g3339 ( 
.A(n_2523),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2467),
.Y(n_3340)
);

BUFx6f_ASAP7_75t_L g3341 ( 
.A(n_2523),
.Y(n_3341)
);

INVx4_ASAP7_75t_L g3342 ( 
.A(n_2546),
.Y(n_3342)
);

OA22x2_ASAP7_75t_L g3343 ( 
.A1(n_2376),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_2697),
.B(n_2),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_2332),
.B(n_3),
.Y(n_3345)
);

INVx4_ASAP7_75t_L g3346 ( 
.A(n_2546),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2467),
.Y(n_3347)
);

BUFx6f_ASAP7_75t_L g3348 ( 
.A(n_2523),
.Y(n_3348)
);

BUFx2_ASAP7_75t_L g3349 ( 
.A(n_2697),
.Y(n_3349)
);

BUFx6f_ASAP7_75t_L g3350 ( 
.A(n_2523),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_2467),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_2467),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_2332),
.B(n_3),
.Y(n_3353)
);

BUFx3_ASAP7_75t_L g3354 ( 
.A(n_2330),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_2465),
.Y(n_3355)
);

INVx2_ASAP7_75t_SL g3356 ( 
.A(n_2468),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_SL g3357 ( 
.A(n_2697),
.B(n_1654),
.Y(n_3357)
);

AND2x4_ASAP7_75t_L g3358 ( 
.A(n_2385),
.B(n_5),
.Y(n_3358)
);

NOR3xp33_ASAP7_75t_L g3359 ( 
.A(n_2342),
.B(n_7),
.C(n_6),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_2697),
.B(n_5),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_2697),
.B(n_5),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_2332),
.B(n_6),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_2465),
.Y(n_3363)
);

AND2x6_ASAP7_75t_L g3364 ( 
.A(n_2687),
.B(n_1654),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_2358),
.B(n_7),
.Y(n_3365)
);

NOR2xp33_ASAP7_75t_L g3366 ( 
.A(n_2358),
.B(n_7),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_2465),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_2467),
.Y(n_3368)
);

INVx4_ASAP7_75t_SL g3369 ( 
.A(n_2330),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_2332),
.B(n_8),
.Y(n_3370)
);

INVx4_ASAP7_75t_L g3371 ( 
.A(n_2546),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_2465),
.Y(n_3372)
);

AND2x4_ASAP7_75t_L g3373 ( 
.A(n_2385),
.B(n_8),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_2465),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_2559),
.A2(n_1274),
.B1(n_1240),
.B2(n_10),
.Y(n_3375)
);

BUFx3_ASAP7_75t_L g3376 ( 
.A(n_2330),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_2332),
.B(n_8),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_SL g3378 ( 
.A(n_3156),
.B(n_3060),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_2735),
.Y(n_3379)
);

AOI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_3007),
.A2(n_1274),
.B(n_1240),
.Y(n_3380)
);

NOR3x1_ASAP7_75t_L g3381 ( 
.A(n_3077),
.B(n_18),
.C(n_9),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_2720),
.B(n_9),
.Y(n_3382)
);

BUFx3_ASAP7_75t_L g3383 ( 
.A(n_2799),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_3060),
.B(n_1240),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3000),
.B(n_9),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_L g3386 ( 
.A(n_3328),
.B(n_11),
.Y(n_3386)
);

CKINVDCx5p33_ASAP7_75t_R g3387 ( 
.A(n_2750),
.Y(n_3387)
);

BUFx12f_ASAP7_75t_SL g3388 ( 
.A(n_3274),
.Y(n_3388)
);

AOI21xp5_ASAP7_75t_L g3389 ( 
.A1(n_3009),
.A2(n_1274),
.B(n_1240),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3000),
.B(n_12),
.Y(n_3390)
);

INVx4_ASAP7_75t_L g3391 ( 
.A(n_2799),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_2791),
.A2(n_1274),
.B1(n_14),
.B2(n_12),
.Y(n_3392)
);

NAND2xp33_ASAP7_75t_L g3393 ( 
.A(n_3062),
.B(n_12),
.Y(n_3393)
);

INVx2_ASAP7_75t_SL g3394 ( 
.A(n_2748),
.Y(n_3394)
);

AOI22xp5_ASAP7_75t_L g3395 ( 
.A1(n_2788),
.A2(n_2782),
.B1(n_2730),
.B2(n_3194),
.Y(n_3395)
);

NAND2xp33_ASAP7_75t_L g3396 ( 
.A(n_3062),
.B(n_13),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_2789),
.Y(n_3397)
);

NOR2xp33_ASAP7_75t_L g3398 ( 
.A(n_2997),
.B(n_13),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3002),
.B(n_13),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2793),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3002),
.B(n_14),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3004),
.B(n_15),
.Y(n_3402)
);

AOI22xp5_ASAP7_75t_L g3403 ( 
.A1(n_2798),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_3004),
.Y(n_3404)
);

NAND2x1p5_ASAP7_75t_L g3405 ( 
.A(n_2748),
.B(n_16),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_2884),
.B(n_17),
.Y(n_3406)
);

O2A1O1Ixp33_ASAP7_75t_L g3407 ( 
.A1(n_3095),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_3407)
);

INVx4_ASAP7_75t_L g3408 ( 
.A(n_2768),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2884),
.B(n_18),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_2769),
.B(n_19),
.Y(n_3410)
);

INVx8_ASAP7_75t_L g3411 ( 
.A(n_2930),
.Y(n_3411)
);

NOR3xp33_ASAP7_75t_L g3412 ( 
.A(n_2771),
.B(n_2881),
.C(n_3043),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_SL g3413 ( 
.A(n_3257),
.B(n_834),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2886),
.B(n_20),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_SL g3415 ( 
.A(n_3334),
.B(n_834),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_2886),
.B(n_3094),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_2894),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3094),
.B(n_20),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_2894),
.Y(n_3419)
);

AND2x4_ASAP7_75t_L g3420 ( 
.A(n_3057),
.B(n_20),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_2898),
.B(n_21),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_2898),
.B(n_21),
.Y(n_3422)
);

BUFx3_ASAP7_75t_L g3423 ( 
.A(n_2731),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3349),
.B(n_835),
.Y(n_3424)
);

A2O1A1Ixp33_ASAP7_75t_L g3425 ( 
.A1(n_3089),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_3425)
);

NOR2xp33_ASAP7_75t_L g3426 ( 
.A(n_2831),
.B(n_22),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_2770),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_2770),
.Y(n_3428)
);

OR2x2_ASAP7_75t_L g3429 ( 
.A(n_3232),
.B(n_3319),
.Y(n_3429)
);

INVx2_ASAP7_75t_SL g3430 ( 
.A(n_2930),
.Y(n_3430)
);

OAI22xp5_ASAP7_75t_L g3431 ( 
.A1(n_3022),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_3431)
);

O2A1O1Ixp33_ASAP7_75t_L g3432 ( 
.A1(n_3203),
.A2(n_26),
.B(n_23),
.C(n_25),
.Y(n_3432)
);

AOI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_2772),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_3050),
.B(n_25),
.Y(n_3434)
);

INVx2_ASAP7_75t_SL g3435 ( 
.A(n_2818),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_2780),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2794),
.Y(n_3437)
);

INVx2_ASAP7_75t_SL g3438 ( 
.A(n_2892),
.Y(n_3438)
);

AND2x2_ASAP7_75t_L g3439 ( 
.A(n_2805),
.B(n_26),
.Y(n_3439)
);

NAND2xp33_ASAP7_75t_L g3440 ( 
.A(n_3062),
.B(n_27),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_2795),
.Y(n_3441)
);

INVx8_ASAP7_75t_L g3442 ( 
.A(n_3337),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_2780),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2784),
.B(n_28),
.Y(n_3444)
);

INVx4_ASAP7_75t_L g3445 ( 
.A(n_3369),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_2733),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3179),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_2803),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_2784),
.B(n_28),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_2757),
.B(n_2835),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_SL g3451 ( 
.A(n_2757),
.B(n_836),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_2847),
.B(n_29),
.Y(n_3452)
);

BUFx5_ASAP7_75t_L g3453 ( 
.A(n_3062),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3206),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3209),
.Y(n_3455)
);

BUFx6f_ASAP7_75t_L g3456 ( 
.A(n_2724),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_3218),
.B(n_836),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3219),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3220),
.Y(n_3459)
);

BUFx8_ASAP7_75t_L g3460 ( 
.A(n_2738),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3222),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2853),
.B(n_29),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_SL g3463 ( 
.A(n_3218),
.B(n_837),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_2756),
.B(n_29),
.Y(n_3464)
);

NOR2xp33_ASAP7_75t_L g3465 ( 
.A(n_2790),
.B(n_30),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3239),
.Y(n_3466)
);

AOI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3191),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_3218),
.B(n_3258),
.Y(n_3468)
);

INVx4_ASAP7_75t_L g3469 ( 
.A(n_3369),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_2756),
.B(n_30),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_2905),
.B(n_31),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_2724),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3261),
.Y(n_3473)
);

HB1xp67_ASAP7_75t_L g3474 ( 
.A(n_3274),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_3258),
.B(n_837),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_2761),
.B(n_2762),
.Y(n_3476)
);

AO22x1_ASAP7_75t_L g3477 ( 
.A1(n_3205),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_3477)
);

OAI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_2736),
.A2(n_32),
.B(n_33),
.Y(n_3478)
);

INVxp67_ASAP7_75t_L g3479 ( 
.A(n_3212),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_2761),
.B(n_33),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_2824),
.Y(n_3481)
);

INVx3_ASAP7_75t_L g3482 ( 
.A(n_3040),
.Y(n_3482)
);

NOR2xp33_ASAP7_75t_L g3483 ( 
.A(n_2895),
.B(n_34),
.Y(n_3483)
);

INVx2_ASAP7_75t_SL g3484 ( 
.A(n_2843),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_SL g3485 ( 
.A(n_3258),
.B(n_838),
.Y(n_3485)
);

CKINVDCx5p33_ASAP7_75t_R g3486 ( 
.A(n_2874),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_2762),
.B(n_35),
.Y(n_3487)
);

INVx3_ASAP7_75t_L g3488 ( 
.A(n_3040),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3267),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2763),
.B(n_35),
.Y(n_3490)
);

NOR2xp33_ASAP7_75t_L g3491 ( 
.A(n_3313),
.B(n_35),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_2763),
.B(n_36),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_2825),
.Y(n_3493)
);

AOI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3235),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_2840),
.B(n_37),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3273),
.Y(n_3496)
);

O2A1O1Ixp5_ASAP7_75t_L g3497 ( 
.A1(n_3357),
.A2(n_41),
.B(n_37),
.C(n_40),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3181),
.Y(n_3498)
);

OAI22xp5_ASAP7_75t_SL g3499 ( 
.A1(n_2926),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_SL g3500 ( 
.A(n_2934),
.B(n_838),
.Y(n_3500)
);

INVx2_ASAP7_75t_SL g3501 ( 
.A(n_2935),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_2902),
.B(n_40),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_L g3503 ( 
.A(n_2845),
.B(n_42),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_2801),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_3504)
);

BUFx8_ASAP7_75t_L g3505 ( 
.A(n_2774),
.Y(n_3505)
);

AOI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_2779),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_3506)
);

AO22x1_ASAP7_75t_L g3507 ( 
.A1(n_2890),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3182),
.Y(n_3508)
);

NOR2x1_ASAP7_75t_L g3509 ( 
.A(n_2985),
.B(n_839),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_2943),
.B(n_46),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3188),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3330),
.B(n_46),
.Y(n_3512)
);

BUFx6f_ASAP7_75t_L g3513 ( 
.A(n_2724),
.Y(n_3513)
);

A2O1A1Ixp33_ASAP7_75t_L g3514 ( 
.A1(n_3092),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_SL g3515 ( 
.A(n_3057),
.B(n_839),
.Y(n_3515)
);

BUFx3_ASAP7_75t_L g3516 ( 
.A(n_2785),
.Y(n_3516)
);

NOR3xp33_ASAP7_75t_L g3517 ( 
.A(n_3359),
.B(n_47),
.C(n_48),
.Y(n_3517)
);

AND2x4_ASAP7_75t_L g3518 ( 
.A(n_2726),
.B(n_47),
.Y(n_3518)
);

AOI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_2896),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3189),
.B(n_50),
.Y(n_3520)
);

INVx2_ASAP7_75t_SL g3521 ( 
.A(n_3186),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3192),
.Y(n_3522)
);

INVx4_ASAP7_75t_L g3523 ( 
.A(n_2758),
.Y(n_3523)
);

NOR2xp33_ASAP7_75t_L g3524 ( 
.A(n_2742),
.B(n_50),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3193),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3195),
.B(n_51),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3196),
.B(n_52),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_2968),
.B(n_52),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3200),
.B(n_52),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3202),
.B(n_53),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3210),
.B(n_53),
.Y(n_3531)
);

NAND2xp33_ASAP7_75t_L g3532 ( 
.A(n_3036),
.B(n_53),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3377),
.A2(n_54),
.B(n_55),
.Y(n_3533)
);

INVx2_ASAP7_75t_SL g3534 ( 
.A(n_3237),
.Y(n_3534)
);

INVx2_ASAP7_75t_SL g3535 ( 
.A(n_3292),
.Y(n_3535)
);

AOI22xp33_ASAP7_75t_L g3536 ( 
.A1(n_2941),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_2745),
.B(n_840),
.Y(n_3537)
);

NOR2xp33_ASAP7_75t_L g3538 ( 
.A(n_2949),
.B(n_54),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3213),
.B(n_56),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3223),
.B(n_3231),
.Y(n_3540)
);

AOI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3180),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3234),
.B(n_58),
.Y(n_3542)
);

AOI21xp5_ASAP7_75t_L g3543 ( 
.A1(n_3370),
.A2(n_58),
.B(n_59),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3244),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_L g3545 ( 
.A(n_3001),
.B(n_2728),
.Y(n_3545)
);

NAND2x1_ASAP7_75t_L g3546 ( 
.A(n_3221),
.B(n_59),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3248),
.B(n_60),
.Y(n_3547)
);

OR2x6_ASAP7_75t_L g3548 ( 
.A(n_3316),
.B(n_60),
.Y(n_3548)
);

AND2x6_ASAP7_75t_L g3549 ( 
.A(n_3075),
.B(n_60),
.Y(n_3549)
);

BUFx6f_ASAP7_75t_L g3550 ( 
.A(n_2732),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_SL g3551 ( 
.A(n_2787),
.B(n_840),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_2982),
.B(n_841),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3251),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_2737),
.B(n_61),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_2965),
.B(n_61),
.Y(n_3555)
);

AND2x6_ASAP7_75t_SL g3556 ( 
.A(n_3316),
.B(n_62),
.Y(n_3556)
);

AND2x6_ASAP7_75t_SL g3557 ( 
.A(n_3260),
.B(n_62),
.Y(n_3557)
);

NAND3xp33_ASAP7_75t_SL g3558 ( 
.A(n_3280),
.B(n_62),
.C(n_63),
.Y(n_3558)
);

OAI22xp5_ASAP7_75t_L g3559 ( 
.A1(n_3022),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3259),
.B(n_3262),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3289),
.Y(n_3561)
);

OAI22xp5_ASAP7_75t_L g3562 ( 
.A1(n_2994),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3264),
.B(n_3336),
.Y(n_3563)
);

INVx2_ASAP7_75t_SL g3564 ( 
.A(n_3279),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3340),
.B(n_66),
.Y(n_3565)
);

CKINVDCx5p33_ASAP7_75t_R g3566 ( 
.A(n_2891),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3347),
.B(n_66),
.Y(n_3567)
);

BUFx5_ASAP7_75t_L g3568 ( 
.A(n_3170),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3351),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_3333),
.A2(n_67),
.B(n_68),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3352),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_SL g3572 ( 
.A(n_2866),
.B(n_841),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3368),
.B(n_67),
.Y(n_3573)
);

AOI21xp5_ASAP7_75t_L g3574 ( 
.A1(n_3345),
.A2(n_67),
.B(n_68),
.Y(n_3574)
);

AOI22x1_ASAP7_75t_L g3575 ( 
.A1(n_2899),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_3575)
);

INVx5_ASAP7_75t_L g3576 ( 
.A(n_2765),
.Y(n_3576)
);

INVx3_ASAP7_75t_L g3577 ( 
.A(n_2726),
.Y(n_3577)
);

AND2x2_ASAP7_75t_L g3578 ( 
.A(n_2965),
.B(n_69),
.Y(n_3578)
);

O2A1O1Ixp33_ASAP7_75t_L g3579 ( 
.A1(n_3353),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_2979),
.B(n_70),
.Y(n_3580)
);

AOI22xp5_ASAP7_75t_L g3581 ( 
.A1(n_3187),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_3581)
);

INVx2_ASAP7_75t_L g3582 ( 
.A(n_3299),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_3362),
.A2(n_72),
.B(n_73),
.Y(n_3583)
);

INVx3_ASAP7_75t_L g3584 ( 
.A(n_3197),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3308),
.Y(n_3585)
);

AOI22xp5_ASAP7_75t_L g3586 ( 
.A1(n_3198),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_3586)
);

AOI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3215),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_2981),
.B(n_2946),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_2773),
.B(n_75),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_2953),
.B(n_2962),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_3104),
.A2(n_75),
.B(n_76),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_SL g3592 ( 
.A(n_3079),
.B(n_842),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_2971),
.B(n_76),
.Y(n_3593)
);

NOR2xp33_ASAP7_75t_L g3594 ( 
.A(n_3012),
.B(n_77),
.Y(n_3594)
);

NOR3xp33_ASAP7_75t_L g3595 ( 
.A(n_2977),
.B(n_77),
.C(n_78),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_2858),
.Y(n_3596)
);

AOI22xp5_ASAP7_75t_L g3597 ( 
.A1(n_3228),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_3597)
);

NAND2xp33_ASAP7_75t_L g3598 ( 
.A(n_3036),
.B(n_79),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3044),
.A2(n_80),
.B(n_81),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_2861),
.Y(n_3600)
);

NOR2xp33_ASAP7_75t_L g3601 ( 
.A(n_2969),
.B(n_80),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_2865),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_2973),
.B(n_80),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3315),
.Y(n_3604)
);

AND2x4_ASAP7_75t_L g3605 ( 
.A(n_3197),
.B(n_81),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3008),
.B(n_3013),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_2869),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3355),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_SL g3609 ( 
.A(n_3068),
.B(n_842),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_2870),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_2752),
.B(n_82),
.Y(n_3611)
);

OAI22xp33_ASAP7_75t_L g3612 ( 
.A1(n_3260),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_2755),
.B(n_83),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2875),
.Y(n_3614)
);

AND2x2_ASAP7_75t_L g3615 ( 
.A(n_2944),
.B(n_83),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_2755),
.B(n_84),
.Y(n_3616)
);

OAI22xp33_ASAP7_75t_L g3617 ( 
.A1(n_3214),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3363),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_2980),
.B(n_843),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_3367),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_SL g3621 ( 
.A(n_2980),
.B(n_843),
.Y(n_3621)
);

NOR2xp67_ASAP7_75t_L g3622 ( 
.A(n_3240),
.B(n_85),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3067),
.B(n_86),
.Y(n_3623)
);

O2A1O1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_2879),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3069),
.B(n_87),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_2815),
.B(n_2739),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_2739),
.B(n_88),
.Y(n_3627)
);

INVx3_ASAP7_75t_L g3628 ( 
.A(n_3240),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_2876),
.Y(n_3629)
);

CKINVDCx5p33_ASAP7_75t_R g3630 ( 
.A(n_3241),
.Y(n_3630)
);

AND2x6_ASAP7_75t_SL g3631 ( 
.A(n_3272),
.B(n_88),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_2741),
.B(n_89),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_2877),
.Y(n_3633)
);

OR2x6_ASAP7_75t_L g3634 ( 
.A(n_3275),
.B(n_90),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_2944),
.B(n_90),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_2741),
.B(n_90),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_2915),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3372),
.Y(n_3638)
);

OR2x2_ASAP7_75t_L g3639 ( 
.A(n_3107),
.B(n_91),
.Y(n_3639)
);

INVx3_ASAP7_75t_L g3640 ( 
.A(n_3283),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3335),
.B(n_3344),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_2743),
.B(n_91),
.Y(n_3642)
);

A2O1A1Ixp33_ASAP7_75t_L g3643 ( 
.A1(n_3056),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_3643)
);

AOI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_3238),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_SL g3645 ( 
.A(n_2980),
.B(n_2987),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3011),
.Y(n_3646)
);

OAI22xp5_ASAP7_75t_SL g3647 ( 
.A1(n_3034),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3647)
);

O2A1O1Ixp5_ASAP7_75t_L g3648 ( 
.A1(n_3233),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_2743),
.B(n_95),
.Y(n_3649)
);

NOR2xp33_ASAP7_75t_L g3650 ( 
.A(n_2966),
.B(n_96),
.Y(n_3650)
);

AND2x2_ASAP7_75t_SL g3651 ( 
.A(n_2985),
.B(n_96),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_2933),
.Y(n_3652)
);

NAND3xp33_ASAP7_75t_L g3653 ( 
.A(n_3375),
.B(n_97),
.C(n_98),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_2933),
.Y(n_3654)
);

AND2x4_ASAP7_75t_L g3655 ( 
.A(n_3283),
.B(n_97),
.Y(n_3655)
);

AOI22xp33_ASAP7_75t_L g3656 ( 
.A1(n_2941),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_3656)
);

INVx6_ASAP7_75t_L g3657 ( 
.A(n_2758),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_2746),
.B(n_98),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_2939),
.Y(n_3659)
);

AND2x6_ASAP7_75t_SL g3660 ( 
.A(n_3035),
.B(n_99),
.Y(n_3660)
);

O2A1O1Ixp5_ASAP7_75t_L g3661 ( 
.A1(n_3233),
.A2(n_103),
.B(n_100),
.C(n_101),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_2746),
.B(n_100),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3269),
.B(n_101),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_2939),
.Y(n_3664)
);

BUFx3_ASAP7_75t_L g3665 ( 
.A(n_3354),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_2987),
.B(n_844),
.Y(n_3666)
);

NOR3x1_ASAP7_75t_L g3667 ( 
.A(n_2859),
.B(n_101),
.C(n_103),
.Y(n_3667)
);

INVxp67_ASAP7_75t_SL g3668 ( 
.A(n_2732),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_SL g3669 ( 
.A(n_2987),
.B(n_844),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3374),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_SL g3671 ( 
.A(n_3338),
.B(n_847),
.Y(n_3671)
);

AOI22xp5_ASAP7_75t_L g3672 ( 
.A1(n_3252),
.A2(n_106),
.B1(n_103),
.B2(n_104),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3360),
.B(n_104),
.Y(n_3673)
);

AOI22xp33_ASAP7_75t_L g3674 ( 
.A1(n_2918),
.A2(n_107),
.B1(n_104),
.B2(n_106),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_SL g3675 ( 
.A(n_3338),
.B(n_847),
.Y(n_3675)
);

AND2x4_ASAP7_75t_L g3676 ( 
.A(n_3293),
.B(n_106),
.Y(n_3676)
);

AOI22xp33_ASAP7_75t_L g3677 ( 
.A1(n_3255),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_3677)
);

INVxp67_ASAP7_75t_L g3678 ( 
.A(n_3253),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3078),
.Y(n_3679)
);

INVx2_ASAP7_75t_SL g3680 ( 
.A(n_3376),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3269),
.B(n_107),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3284),
.B(n_109),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_SL g3683 ( 
.A(n_3358),
.B(n_3373),
.Y(n_3683)
);

BUFx3_ASAP7_75t_L g3684 ( 
.A(n_2860),
.Y(n_3684)
);

INVx3_ASAP7_75t_L g3685 ( 
.A(n_3293),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3284),
.B(n_110),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3123),
.Y(n_3687)
);

AOI22xp33_ASAP7_75t_L g3688 ( 
.A1(n_3255),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_3688)
);

NAND2x1p5_ASAP7_75t_L g3689 ( 
.A(n_3301),
.B(n_110),
.Y(n_3689)
);

BUFx6f_ASAP7_75t_L g3690 ( 
.A(n_2732),
.Y(n_3690)
);

AOI22xp5_ASAP7_75t_L g3691 ( 
.A1(n_3268),
.A2(n_114),
.B1(n_111),
.B2(n_113),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_L g3692 ( 
.A(n_2975),
.B(n_113),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_L g3693 ( 
.A1(n_2826),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3294),
.B(n_114),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_SL g3695 ( 
.A(n_3358),
.B(n_848),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3294),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3296),
.B(n_115),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3296),
.B(n_116),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3304),
.B(n_116),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3304),
.Y(n_3700)
);

INVxp67_ASAP7_75t_L g3701 ( 
.A(n_3297),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3307),
.Y(n_3702)
);

NAND2x1p5_ASAP7_75t_L g3703 ( 
.A(n_3301),
.B(n_117),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3124),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3307),
.B(n_3311),
.Y(n_3705)
);

OR2x2_ASAP7_75t_L g3706 ( 
.A(n_3310),
.B(n_117),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3311),
.B(n_117),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3312),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3312),
.B(n_118),
.Y(n_3709)
);

NOR2xp33_ASAP7_75t_L g3710 ( 
.A(n_2900),
.B(n_2927),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3314),
.B(n_3325),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3361),
.B(n_118),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3314),
.B(n_119),
.Y(n_3713)
);

AOI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_2826),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3325),
.B(n_119),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3126),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3229),
.B(n_120),
.Y(n_3717)
);

NOR2xp67_ASAP7_75t_L g3718 ( 
.A(n_3309),
.B(n_3320),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3229),
.B(n_3318),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_SL g3720 ( 
.A(n_3373),
.B(n_848),
.Y(n_3720)
);

NOR2x2_ASAP7_75t_L g3721 ( 
.A(n_3306),
.B(n_121),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_2804),
.B(n_849),
.Y(n_3722)
);

BUFx6f_ASAP7_75t_L g3723 ( 
.A(n_2766),
.Y(n_3723)
);

OAI22xp33_ASAP7_75t_L g3724 ( 
.A1(n_2996),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_3724)
);

INVx8_ASAP7_75t_L g3725 ( 
.A(n_2721),
.Y(n_3725)
);

CKINVDCx5p33_ASAP7_75t_R g3726 ( 
.A(n_3265),
.Y(n_3726)
);

NOR2x2_ASAP7_75t_L g3727 ( 
.A(n_2873),
.B(n_125),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_L g3728 ( 
.A1(n_3083),
.A2(n_3366),
.B1(n_3365),
.B2(n_2802),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_3201),
.B(n_124),
.Y(n_3729)
);

BUFx3_ASAP7_75t_L g3730 ( 
.A(n_2923),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3326),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3326),
.B(n_124),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_2816),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3332),
.B(n_124),
.Y(n_3734)
);

AND2x4_ASAP7_75t_SL g3735 ( 
.A(n_3309),
.B(n_125),
.Y(n_3735)
);

BUFx6f_ASAP7_75t_SL g3736 ( 
.A(n_3073),
.Y(n_3736)
);

NAND2xp33_ASAP7_75t_L g3737 ( 
.A(n_3036),
.B(n_125),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3332),
.B(n_126),
.Y(n_3738)
);

AOI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_2729),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_2816),
.Y(n_3740)
);

AOI22xp5_ASAP7_75t_L g3741 ( 
.A1(n_2836),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_3741)
);

NOR2xp33_ASAP7_75t_L g3742 ( 
.A(n_3217),
.B(n_128),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_2764),
.Y(n_3743)
);

OAI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_2767),
.A2(n_129),
.B(n_130),
.Y(n_3744)
);

AOI22xp5_ASAP7_75t_L g3745 ( 
.A1(n_2802),
.A2(n_2833),
.B1(n_2819),
.B2(n_2862),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_2775),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_2753),
.B(n_130),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_2754),
.B(n_130),
.Y(n_3748)
);

NAND2x1p5_ASAP7_75t_L g3749 ( 
.A(n_3320),
.B(n_131),
.Y(n_3749)
);

NOR2xp67_ASAP7_75t_L g3750 ( 
.A(n_3323),
.B(n_131),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_2759),
.B(n_131),
.Y(n_3751)
);

AND2x6_ASAP7_75t_SL g3752 ( 
.A(n_3211),
.B(n_132),
.Y(n_3752)
);

INVx4_ASAP7_75t_L g3753 ( 
.A(n_3323),
.Y(n_3753)
);

NOR2xp33_ASAP7_75t_L g3754 ( 
.A(n_3254),
.B(n_132),
.Y(n_3754)
);

CKINVDCx5p33_ASAP7_75t_R g3755 ( 
.A(n_3015),
.Y(n_3755)
);

NOR2xp33_ASAP7_75t_L g3756 ( 
.A(n_3287),
.B(n_133),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_2760),
.B(n_133),
.Y(n_3757)
);

INVx2_ASAP7_75t_SL g3758 ( 
.A(n_3342),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_2786),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_2948),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_SL g3761 ( 
.A(n_2804),
.B(n_850),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_2744),
.B(n_133),
.Y(n_3762)
);

AOI22xp33_ASAP7_75t_L g3763 ( 
.A1(n_2919),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_3763)
);

INVxp67_ASAP7_75t_L g3764 ( 
.A(n_2723),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_2854),
.B(n_134),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_2911),
.B(n_134),
.Y(n_3766)
);

OAI22x1_ASAP7_75t_L g3767 ( 
.A1(n_2817),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_3767)
);

NAND2xp33_ASAP7_75t_L g3768 ( 
.A(n_3036),
.B(n_135),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_2952),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_2958),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_2854),
.B(n_136),
.Y(n_3771)
);

AOI22xp33_ASAP7_75t_L g3772 ( 
.A1(n_2919),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_3772)
);

NOR2xp33_ASAP7_75t_L g3773 ( 
.A(n_2950),
.B(n_137),
.Y(n_3773)
);

INVx8_ASAP7_75t_L g3774 ( 
.A(n_2765),
.Y(n_3774)
);

AO22x1_ASAP7_75t_L g3775 ( 
.A1(n_3088),
.A2(n_2995),
.B1(n_2765),
.B2(n_3364),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_2849),
.B(n_850),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_2959),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3019),
.B(n_138),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_2778),
.B(n_140),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_2839),
.B(n_140),
.Y(n_3780)
);

OAI221xp5_ASAP7_75t_L g3781 ( 
.A1(n_3208),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.C(n_143),
.Y(n_3781)
);

OAI22xp5_ASAP7_75t_L g3782 ( 
.A1(n_2994),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_3782)
);

NOR2xp33_ASAP7_75t_L g3783 ( 
.A(n_3190),
.B(n_144),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_2778),
.B(n_145),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_2781),
.B(n_145),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_2781),
.B(n_146),
.Y(n_3786)
);

BUFx8_ASAP7_75t_L g3787 ( 
.A(n_3074),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_2834),
.B(n_146),
.Y(n_3788)
);

NOR3xp33_ASAP7_75t_L g3789 ( 
.A(n_2945),
.B(n_146),
.C(n_147),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_2834),
.B(n_147),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_2925),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_3791)
);

OR2x2_ASAP7_75t_L g3792 ( 
.A(n_2822),
.B(n_148),
.Y(n_3792)
);

BUFx2_ASAP7_75t_L g3793 ( 
.A(n_3342),
.Y(n_3793)
);

NOR2xp33_ASAP7_75t_L g3794 ( 
.A(n_3263),
.B(n_148),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3051),
.A2(n_150),
.B(n_151),
.Y(n_3795)
);

OAI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3052),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_3796)
);

NAND2x1_ASAP7_75t_L g3797 ( 
.A(n_3221),
.B(n_152),
.Y(n_3797)
);

NOR2x1p5_ASAP7_75t_L g3798 ( 
.A(n_3346),
.B(n_153),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_SL g3799 ( 
.A(n_3346),
.B(n_851),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_SL g3800 ( 
.A(n_3371),
.B(n_851),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_2837),
.B(n_153),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_2837),
.B(n_153),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_2964),
.Y(n_3803)
);

OAI22xp33_ASAP7_75t_L g3804 ( 
.A1(n_3343),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_3804)
);

NOR2xp33_ASAP7_75t_L g3805 ( 
.A(n_3266),
.B(n_154),
.Y(n_3805)
);

BUFx3_ASAP7_75t_L g3806 ( 
.A(n_3059),
.Y(n_3806)
);

NOR2xp33_ASAP7_75t_L g3807 ( 
.A(n_3271),
.B(n_155),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_2960),
.B(n_156),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_2960),
.B(n_156),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_SL g3810 ( 
.A(n_3371),
.B(n_852),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_2978),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_SL g3812 ( 
.A(n_2722),
.B(n_852),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_2792),
.Y(n_3813)
);

OR2x2_ASAP7_75t_L g3814 ( 
.A(n_2850),
.B(n_157),
.Y(n_3814)
);

AOI22xp5_ASAP7_75t_L g3815 ( 
.A1(n_3224),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_2796),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_SL g3817 ( 
.A(n_2722),
.B(n_853),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_2967),
.B(n_157),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_2967),
.B(n_158),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3082),
.B(n_158),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3125),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_L g3822 ( 
.A(n_2983),
.B(n_2998),
.Y(n_3822)
);

NOR2xp33_ASAP7_75t_L g3823 ( 
.A(n_2747),
.B(n_2871),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_2893),
.B(n_159),
.Y(n_3824)
);

NOR2xp33_ASAP7_75t_L g3825 ( 
.A(n_2970),
.B(n_160),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3130),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_2989),
.B(n_160),
.Y(n_3827)
);

INVx3_ASAP7_75t_L g3828 ( 
.A(n_2991),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_2893),
.B(n_2903),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_2809),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_2903),
.B(n_161),
.Y(n_3831)
);

INVx1_ASAP7_75t_SL g3832 ( 
.A(n_3020),
.Y(n_3832)
);

AND2x6_ASAP7_75t_SL g3833 ( 
.A(n_3281),
.B(n_161),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_SL g3834 ( 
.A(n_2991),
.B(n_161),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_2956),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_2993),
.B(n_162),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_2725),
.B(n_162),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_2956),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_2811),
.B(n_163),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_2883),
.B(n_163),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_2885),
.B(n_163),
.Y(n_3841)
);

INVx6_ASAP7_75t_L g3842 ( 
.A(n_2827),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_2814),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_2913),
.B(n_164),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_2957),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_2807),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_L g3847 ( 
.A1(n_2925),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_2951),
.B(n_3058),
.Y(n_3848)
);

BUFx6f_ASAP7_75t_L g3849 ( 
.A(n_2766),
.Y(n_3849)
);

AOI22xp5_ASAP7_75t_L g3850 ( 
.A1(n_3286),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_3850)
);

INVxp67_ASAP7_75t_L g3851 ( 
.A(n_2727),
.Y(n_3851)
);

INVx2_ASAP7_75t_SL g3852 ( 
.A(n_2872),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3058),
.B(n_165),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_2957),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3135),
.B(n_166),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_2961),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_2846),
.B(n_167),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_2777),
.B(n_167),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_2783),
.B(n_167),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_SL g3860 ( 
.A(n_2740),
.B(n_853),
.Y(n_3860)
);

BUFx6f_ASAP7_75t_L g3861 ( 
.A(n_2766),
.Y(n_3861)
);

HB1xp67_ASAP7_75t_L g3862 ( 
.A(n_2823),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_2820),
.B(n_168),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_2821),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_2961),
.Y(n_3865)
);

INVxp67_ASAP7_75t_L g3866 ( 
.A(n_3135),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3329),
.B(n_168),
.Y(n_3867)
);

NOR2xp33_ASAP7_75t_R g3868 ( 
.A(n_2841),
.B(n_168),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3331),
.B(n_169),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_2928),
.B(n_169),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_2928),
.B(n_170),
.Y(n_3871)
);

INVxp67_ASAP7_75t_L g3872 ( 
.A(n_2992),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3216),
.B(n_3245),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3282),
.B(n_3285),
.Y(n_3874)
);

AOI22xp33_ASAP7_75t_L g3875 ( 
.A1(n_2955),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_3875)
);

INVx2_ASAP7_75t_SL g3876 ( 
.A(n_3045),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_SL g3877 ( 
.A(n_2740),
.B(n_854),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_SL g3878 ( 
.A(n_2751),
.B(n_855),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3288),
.B(n_3302),
.Y(n_3879)
);

OAI21xp5_ASAP7_75t_L g3880 ( 
.A1(n_3120),
.A2(n_171),
.B(n_172),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_SL g3881 ( 
.A(n_2751),
.B(n_855),
.Y(n_3881)
);

AND2x6_ASAP7_75t_SL g3882 ( 
.A(n_3298),
.B(n_171),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3005),
.B(n_172),
.Y(n_3883)
);

AOI22xp33_ASAP7_75t_L g3884 ( 
.A1(n_2955),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_3183),
.B(n_856),
.Y(n_3885)
);

BUFx3_ASAP7_75t_L g3886 ( 
.A(n_2976),
.Y(n_3886)
);

BUFx6f_ASAP7_75t_L g3887 ( 
.A(n_2797),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_L g3888 ( 
.A(n_3086),
.B(n_3327),
.Y(n_3888)
);

NOR2x1p5_ASAP7_75t_L g3889 ( 
.A(n_2937),
.B(n_173),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_2880),
.B(n_174),
.Y(n_3890)
);

O2A1O1Ixp5_ASAP7_75t_L g3891 ( 
.A1(n_3246),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_3183),
.B(n_856),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3150),
.B(n_176),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_3137),
.B(n_176),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3139),
.B(n_177),
.Y(n_3895)
);

NOR2xp33_ASAP7_75t_SL g3896 ( 
.A(n_2765),
.B(n_3221),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3017),
.B(n_177),
.Y(n_3897)
);

A2O1A1Ixp33_ASAP7_75t_L g3898 ( 
.A1(n_3085),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_3898)
);

NOR2xp67_ASAP7_75t_L g3899 ( 
.A(n_2937),
.B(n_178),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3021),
.B(n_2917),
.Y(n_3900)
);

AND2x6_ASAP7_75t_SL g3901 ( 
.A(n_2776),
.B(n_3049),
.Y(n_3901)
);

AOI22xp33_ASAP7_75t_L g3902 ( 
.A1(n_3103),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_3902)
);

INVx2_ASAP7_75t_SL g3903 ( 
.A(n_3045),
.Y(n_3903)
);

BUFx3_ASAP7_75t_L g3904 ( 
.A(n_2988),
.Y(n_3904)
);

NAND2xp33_ASAP7_75t_L g3905 ( 
.A(n_3088),
.B(n_180),
.Y(n_3905)
);

INVx2_ASAP7_75t_SL g3906 ( 
.A(n_3321),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_2917),
.B(n_180),
.Y(n_3907)
);

NOR3xp33_ASAP7_75t_L g3908 ( 
.A(n_2942),
.B(n_181),
.C(n_182),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3117),
.B(n_3129),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_2999),
.Y(n_3910)
);

NOR2xp33_ASAP7_75t_SL g3911 ( 
.A(n_3221),
.B(n_181),
.Y(n_3911)
);

AOI22xp5_ASAP7_75t_SL g3912 ( 
.A1(n_3184),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_3912)
);

NOR2xp33_ASAP7_75t_L g3913 ( 
.A(n_3091),
.B(n_182),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_2999),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3023),
.Y(n_3915)
);

NOR2xp33_ASAP7_75t_L g3916 ( 
.A(n_3041),
.B(n_183),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3117),
.B(n_183),
.Y(n_3917)
);

AND2x4_ASAP7_75t_SL g3918 ( 
.A(n_3356),
.B(n_184),
.Y(n_3918)
);

NOR2x2_ASAP7_75t_L g3919 ( 
.A(n_2827),
.B(n_185),
.Y(n_3919)
);

AND2x2_ASAP7_75t_L g3920 ( 
.A(n_3052),
.B(n_184),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_2842),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_SL g3922 ( 
.A(n_3184),
.B(n_3204),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_L g3923 ( 
.A(n_3014),
.B(n_184),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_2848),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3112),
.B(n_3055),
.Y(n_3925)
);

NOR2xp33_ASAP7_75t_L g3926 ( 
.A(n_3147),
.B(n_185),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3028),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3305),
.B(n_3105),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3030),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3105),
.B(n_185),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3098),
.B(n_186),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_2851),
.Y(n_3932)
);

INVx3_ASAP7_75t_L g3933 ( 
.A(n_2797),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3114),
.B(n_186),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3114),
.B(n_186),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_2882),
.B(n_187),
.Y(n_3936)
);

NOR2xp33_ASAP7_75t_L g3937 ( 
.A(n_3032),
.B(n_187),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3113),
.B(n_188),
.Y(n_3938)
);

INVx3_ASAP7_75t_L g3939 ( 
.A(n_2797),
.Y(n_3939)
);

A2O1A1Ixp33_ASAP7_75t_L g3940 ( 
.A1(n_3031),
.A2(n_3152),
.B(n_3103),
.C(n_3115),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_2899),
.B(n_188),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3133),
.B(n_189),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3033),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3047),
.B(n_190),
.Y(n_3944)
);

AOI221xp5_ASAP7_75t_L g3945 ( 
.A1(n_3101),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.C(n_193),
.Y(n_3945)
);

AOI22xp5_ASAP7_75t_L g3946 ( 
.A1(n_3093),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_2972),
.B(n_192),
.Y(n_3947)
);

NOR2xp33_ASAP7_75t_L g3948 ( 
.A(n_3064),
.B(n_193),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_2852),
.Y(n_3949)
);

INVx2_ASAP7_75t_SL g3950 ( 
.A(n_2832),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3404),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_SL g3952 ( 
.A(n_3651),
.B(n_3204),
.Y(n_3952)
);

AND2x4_ASAP7_75t_L g3953 ( 
.A(n_3718),
.B(n_3003),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3379),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3710),
.B(n_3066),
.Y(n_3955)
);

AOI22xp5_ASAP7_75t_L g3956 ( 
.A1(n_3548),
.A2(n_3236),
.B1(n_3291),
.B2(n_3276),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3696),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3417),
.Y(n_3958)
);

AND2x4_ASAP7_75t_L g3959 ( 
.A(n_3753),
.B(n_3003),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3412),
.A2(n_3247),
.B1(n_3250),
.B2(n_3246),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3588),
.B(n_2972),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3397),
.Y(n_3962)
);

BUFx3_ASAP7_75t_L g3963 ( 
.A(n_3460),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3400),
.Y(n_3964)
);

INVx1_ASAP7_75t_SL g3965 ( 
.A(n_3383),
.Y(n_3965)
);

INVx4_ASAP7_75t_L g3966 ( 
.A(n_3391),
.Y(n_3966)
);

BUFx12f_ASAP7_75t_L g3967 ( 
.A(n_3387),
.Y(n_3967)
);

NOR2x1p5_ASAP7_75t_L g3968 ( 
.A(n_3408),
.B(n_3391),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3419),
.Y(n_3969)
);

AND2x4_ASAP7_75t_L g3970 ( 
.A(n_3753),
.B(n_3006),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3626),
.B(n_3733),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3700),
.Y(n_3972)
);

CKINVDCx5p33_ASAP7_75t_R g3973 ( 
.A(n_3630),
.Y(n_3973)
);

CKINVDCx6p67_ASAP7_75t_R g3974 ( 
.A(n_3442),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3740),
.B(n_3038),
.Y(n_3975)
);

OAI221xp5_ASAP7_75t_L g3976 ( 
.A1(n_3745),
.A2(n_3122),
.B1(n_3119),
.B2(n_2812),
.C(n_3155),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3555),
.B(n_3225),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3702),
.Y(n_3978)
);

AND2x4_ASAP7_75t_L g3979 ( 
.A(n_3577),
.B(n_3006),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3517),
.A2(n_3250),
.B1(n_3270),
.B2(n_3247),
.Y(n_3980)
);

BUFx2_ASAP7_75t_L g3981 ( 
.A(n_3388),
.Y(n_3981)
);

INVx2_ASAP7_75t_SL g3982 ( 
.A(n_3411),
.Y(n_3982)
);

BUFx3_ASAP7_75t_L g3983 ( 
.A(n_3460),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3416),
.B(n_3039),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3437),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3641),
.B(n_3225),
.Y(n_3986)
);

INVx2_ASAP7_75t_L g3987 ( 
.A(n_3708),
.Y(n_3987)
);

INVxp33_ASAP7_75t_SL g3988 ( 
.A(n_3868),
.Y(n_3988)
);

AND2x4_ASAP7_75t_L g3989 ( 
.A(n_3577),
.B(n_3010),
.Y(n_3989)
);

BUFx3_ASAP7_75t_L g3990 ( 
.A(n_3505),
.Y(n_3990)
);

INVx2_ASAP7_75t_L g3991 ( 
.A(n_3731),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3441),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3678),
.B(n_3154),
.Y(n_3993)
);

BUFx2_ASAP7_75t_L g3994 ( 
.A(n_3684),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3701),
.B(n_3158),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3448),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3427),
.Y(n_3997)
);

INVx5_ASAP7_75t_L g3998 ( 
.A(n_3548),
.Y(n_3998)
);

INVxp67_ASAP7_75t_L g3999 ( 
.A(n_3429),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3481),
.B(n_3097),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3493),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3498),
.B(n_3099),
.Y(n_4002)
);

OR2x2_ASAP7_75t_L g4003 ( 
.A(n_3909),
.B(n_3276),
.Y(n_4003)
);

INVx5_ASAP7_75t_L g4004 ( 
.A(n_3774),
.Y(n_4004)
);

OAI22xp5_ASAP7_75t_L g4005 ( 
.A1(n_3866),
.A2(n_3132),
.B1(n_3291),
.B2(n_3270),
.Y(n_4005)
);

OAI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3650),
.A2(n_3169),
.B(n_3134),
.Y(n_4006)
);

AND2x4_ASAP7_75t_L g4007 ( 
.A(n_3584),
.B(n_3010),
.Y(n_4007)
);

INVx1_ASAP7_75t_SL g4008 ( 
.A(n_3423),
.Y(n_4008)
);

INVxp67_ASAP7_75t_L g4009 ( 
.A(n_3503),
.Y(n_4009)
);

OAI21xp33_ASAP7_75t_L g4010 ( 
.A1(n_3728),
.A2(n_3132),
.B(n_3134),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3508),
.B(n_3101),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3511),
.Y(n_4012)
);

BUFx4f_ASAP7_75t_SL g4013 ( 
.A(n_3505),
.Y(n_4013)
);

INVx2_ASAP7_75t_SL g4014 ( 
.A(n_3411),
.Y(n_4014)
);

BUFx3_ASAP7_75t_L g4015 ( 
.A(n_3516),
.Y(n_4015)
);

AOI22xp33_ASAP7_75t_SL g4016 ( 
.A1(n_3499),
.A2(n_3393),
.B1(n_3440),
.B2(n_3396),
.Y(n_4016)
);

CKINVDCx5p33_ASAP7_75t_R g4017 ( 
.A(n_3486),
.Y(n_4017)
);

BUFx6f_ASAP7_75t_L g4018 ( 
.A(n_3456),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3522),
.B(n_2901),
.Y(n_4019)
);

NOR2xp33_ASAP7_75t_SL g4020 ( 
.A(n_3408),
.B(n_3242),
.Y(n_4020)
);

INVx3_ASAP7_75t_L g4021 ( 
.A(n_3774),
.Y(n_4021)
);

INVx5_ASAP7_75t_L g4022 ( 
.A(n_3634),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3525),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3544),
.B(n_3153),
.Y(n_4024)
);

BUFx6f_ASAP7_75t_L g4025 ( 
.A(n_3456),
.Y(n_4025)
);

BUFx3_ASAP7_75t_L g4026 ( 
.A(n_3665),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_L g4027 ( 
.A(n_3553),
.B(n_3140),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3569),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3571),
.B(n_2984),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3428),
.Y(n_4030)
);

NOR2xp33_ASAP7_75t_L g4031 ( 
.A(n_3395),
.B(n_3048),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3596),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3600),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3602),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3607),
.Y(n_4035)
);

NAND3xp33_ASAP7_75t_L g4036 ( 
.A(n_3575),
.B(n_3018),
.C(n_2984),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3436),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3443),
.Y(n_4038)
);

BUFx2_ASAP7_75t_L g4039 ( 
.A(n_3793),
.Y(n_4039)
);

INVx2_ASAP7_75t_SL g4040 ( 
.A(n_3755),
.Y(n_4040)
);

BUFx2_ASAP7_75t_L g4041 ( 
.A(n_3886),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3679),
.Y(n_4042)
);

AND2x4_ASAP7_75t_L g4043 ( 
.A(n_3584),
.B(n_3053),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3687),
.Y(n_4044)
);

OAI22xp33_ASAP7_75t_L g4045 ( 
.A1(n_3634),
.A2(n_3046),
.B1(n_2857),
.B2(n_3071),
.Y(n_4045)
);

INVx3_ASAP7_75t_L g4046 ( 
.A(n_3576),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3719),
.A2(n_3018),
.B1(n_3042),
.B2(n_3037),
.Y(n_4047)
);

BUFx2_ASAP7_75t_L g4048 ( 
.A(n_3904),
.Y(n_4048)
);

INVxp67_ASAP7_75t_L g4049 ( 
.A(n_3474),
.Y(n_4049)
);

AOI22xp5_ASAP7_75t_L g4050 ( 
.A1(n_3426),
.A2(n_3109),
.B1(n_2995),
.B2(n_3088),
.Y(n_4050)
);

CKINVDCx5p33_ASAP7_75t_R g4051 ( 
.A(n_3442),
.Y(n_4051)
);

CKINVDCx6p67_ASAP7_75t_R g4052 ( 
.A(n_3725),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3704),
.Y(n_4053)
);

INVx2_ASAP7_75t_L g4054 ( 
.A(n_3646),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3716),
.Y(n_4055)
);

INVx2_ASAP7_75t_L g4056 ( 
.A(n_3446),
.Y(n_4056)
);

INVx2_ASAP7_75t_SL g4057 ( 
.A(n_3657),
.Y(n_4057)
);

AOI22xp5_ASAP7_75t_L g4058 ( 
.A1(n_3410),
.A2(n_2995),
.B1(n_3088),
.B2(n_3080),
.Y(n_4058)
);

NAND2x1_ASAP7_75t_L g4059 ( 
.A(n_3456),
.B(n_3242),
.Y(n_4059)
);

BUFx6f_ASAP7_75t_L g4060 ( 
.A(n_3472),
.Y(n_4060)
);

INVx2_ASAP7_75t_SL g4061 ( 
.A(n_3657),
.Y(n_4061)
);

INVx3_ASAP7_75t_L g4062 ( 
.A(n_3576),
.Y(n_4062)
);

AND2x4_ASAP7_75t_L g4063 ( 
.A(n_3628),
.B(n_3053),
.Y(n_4063)
);

OR2x6_ASAP7_75t_L g4064 ( 
.A(n_3725),
.B(n_2914),
.Y(n_4064)
);

HB1xp67_ASAP7_75t_L g4065 ( 
.A(n_3479),
.Y(n_4065)
);

BUFx12f_ASAP7_75t_L g4066 ( 
.A(n_3726),
.Y(n_4066)
);

HB1xp67_ASAP7_75t_L g4067 ( 
.A(n_3832),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3447),
.Y(n_4068)
);

AND2x4_ASAP7_75t_L g4069 ( 
.A(n_3628),
.B(n_3084),
.Y(n_4069)
);

AOI21x1_ASAP7_75t_L g4070 ( 
.A1(n_3775),
.A2(n_3090),
.B(n_3151),
.Y(n_4070)
);

AND2x4_ASAP7_75t_L g4071 ( 
.A(n_3640),
.B(n_3084),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3826),
.B(n_3037),
.Y(n_4072)
);

CKINVDCx5p33_ASAP7_75t_R g4073 ( 
.A(n_3566),
.Y(n_4073)
);

NAND2x1p5_ASAP7_75t_L g4074 ( 
.A(n_3445),
.B(n_3102),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3454),
.Y(n_4075)
);

BUFx3_ASAP7_75t_L g4076 ( 
.A(n_3787),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3821),
.Y(n_4077)
);

AND2x6_ASAP7_75t_SL g4078 ( 
.A(n_3721),
.B(n_3042),
.Y(n_4078)
);

AND3x1_ASAP7_75t_SL g4079 ( 
.A(n_3889),
.B(n_193),
.C(n_194),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3540),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_L g4081 ( 
.A(n_3491),
.B(n_3108),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3560),
.B(n_3143),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3455),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3563),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_3590),
.Y(n_4085)
);

AOI22xp5_ASAP7_75t_L g4086 ( 
.A1(n_3692),
.A2(n_2995),
.B1(n_3076),
.B2(n_3171),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3606),
.B(n_3054),
.Y(n_4087)
);

HB1xp67_ASAP7_75t_L g4088 ( 
.A(n_3829),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_3538),
.B(n_3063),
.Y(n_4089)
);

CKINVDCx5p33_ASAP7_75t_R g4090 ( 
.A(n_3787),
.Y(n_4090)
);

CKINVDCx5p33_ASAP7_75t_R g4091 ( 
.A(n_3556),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_3458),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3459),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3578),
.B(n_3167),
.Y(n_4094)
);

NOR2xp33_ASAP7_75t_L g4095 ( 
.A(n_3764),
.B(n_3121),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_SL g4096 ( 
.A(n_3834),
.B(n_2800),
.Y(n_4096)
);

OR2x6_ASAP7_75t_L g4097 ( 
.A(n_3445),
.B(n_2914),
.Y(n_4097)
);

CKINVDCx5p33_ASAP7_75t_R g4098 ( 
.A(n_3557),
.Y(n_4098)
);

BUFx3_ASAP7_75t_L g4099 ( 
.A(n_3730),
.Y(n_4099)
);

BUFx2_ASAP7_75t_L g4100 ( 
.A(n_3806),
.Y(n_4100)
);

BUFx3_ASAP7_75t_L g4101 ( 
.A(n_3501),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3610),
.Y(n_4102)
);

AOI22xp5_ASAP7_75t_L g4103 ( 
.A1(n_3594),
.A2(n_3090),
.B1(n_3256),
.B2(n_3242),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3825),
.B(n_3065),
.Y(n_4104)
);

INVx5_ASAP7_75t_L g4105 ( 
.A(n_3469),
.Y(n_4105)
);

AND2x4_ASAP7_75t_L g4106 ( 
.A(n_3640),
.B(n_2800),
.Y(n_4106)
);

CKINVDCx5p33_ASAP7_75t_R g4107 ( 
.A(n_3631),
.Y(n_4107)
);

BUFx6f_ASAP7_75t_L g4108 ( 
.A(n_3472),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3827),
.B(n_3081),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_3937),
.B(n_3096),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_3471),
.B(n_3100),
.Y(n_4111)
);

BUFx3_ASAP7_75t_L g4112 ( 
.A(n_3521),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3439),
.B(n_3110),
.Y(n_4113)
);

CKINVDCx5p33_ASAP7_75t_R g4114 ( 
.A(n_3736),
.Y(n_4114)
);

HB1xp67_ASAP7_75t_L g4115 ( 
.A(n_3942),
.Y(n_4115)
);

BUFx6f_ASAP7_75t_L g4116 ( 
.A(n_3472),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_3461),
.Y(n_4117)
);

AOI22xp5_ASAP7_75t_L g4118 ( 
.A1(n_3483),
.A2(n_3256),
.B1(n_3300),
.B2(n_3242),
.Y(n_4118)
);

INVx1_ASAP7_75t_SL g4119 ( 
.A(n_3852),
.Y(n_4119)
);

BUFx3_ASAP7_75t_L g4120 ( 
.A(n_3534),
.Y(n_4120)
);

INVx2_ASAP7_75t_L g4121 ( 
.A(n_3466),
.Y(n_4121)
);

NOR2xp33_ASAP7_75t_L g4122 ( 
.A(n_3851),
.B(n_3102),
.Y(n_4122)
);

BUFx3_ASAP7_75t_L g4123 ( 
.A(n_3535),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_3896),
.B(n_2800),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3614),
.Y(n_4125)
);

INVxp67_ASAP7_75t_SL g4126 ( 
.A(n_3683),
.Y(n_4126)
);

HB1xp67_ASAP7_75t_L g4127 ( 
.A(n_3900),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3476),
.B(n_3111),
.Y(n_4128)
);

CKINVDCx8_ASAP7_75t_R g4129 ( 
.A(n_3660),
.Y(n_4129)
);

A2O1A1Ixp33_ASAP7_75t_L g4130 ( 
.A1(n_3923),
.A2(n_3174),
.B(n_3106),
.C(n_3016),
.Y(n_4130)
);

OR2x4_ASAP7_75t_L g4131 ( 
.A(n_3639),
.B(n_3144),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3629),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3705),
.Y(n_4133)
);

BUFx6f_ASAP7_75t_L g4134 ( 
.A(n_3513),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_3633),
.Y(n_4135)
);

CKINVDCx5p33_ASAP7_75t_R g4136 ( 
.A(n_3736),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_3473),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3398),
.B(n_2990),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3637),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3489),
.Y(n_4140)
);

NAND2x1p5_ASAP7_75t_L g4141 ( 
.A(n_3469),
.B(n_3106),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_3496),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3561),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3915),
.Y(n_4144)
);

BUFx3_ASAP7_75t_L g4145 ( 
.A(n_3564),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3927),
.Y(n_4146)
);

AND2x2_ASAP7_75t_L g4147 ( 
.A(n_3855),
.B(n_3025),
.Y(n_4147)
);

AOI22xp33_ASAP7_75t_L g4148 ( 
.A1(n_3908),
.A2(n_3087),
.B1(n_3300),
.B2(n_3256),
.Y(n_4148)
);

BUFx2_ASAP7_75t_L g4149 ( 
.A(n_3685),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3929),
.Y(n_4150)
);

INVx2_ASAP7_75t_SL g4151 ( 
.A(n_3842),
.Y(n_4151)
);

BUFx2_ASAP7_75t_L g4152 ( 
.A(n_3685),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3582),
.Y(n_4153)
);

CKINVDCx5p33_ASAP7_75t_R g4154 ( 
.A(n_3752),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_3585),
.Y(n_4155)
);

NOR2xp33_ASAP7_75t_L g4156 ( 
.A(n_3925),
.B(n_3148),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_3873),
.B(n_3029),
.Y(n_4157)
);

AND2x6_ASAP7_75t_L g4158 ( 
.A(n_3453),
.B(n_2868),
.Y(n_4158)
);

INVx2_ASAP7_75t_SL g4159 ( 
.A(n_3842),
.Y(n_4159)
);

NOR2xp33_ASAP7_75t_L g4160 ( 
.A(n_3888),
.B(n_3146),
.Y(n_4160)
);

BUFx3_ASAP7_75t_L g4161 ( 
.A(n_3680),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_3604),
.Y(n_4162)
);

BUFx4f_ASAP7_75t_L g4163 ( 
.A(n_3405),
.Y(n_4163)
);

INVx5_ASAP7_75t_L g4164 ( 
.A(n_3523),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_3943),
.Y(n_4165)
);

BUFx3_ASAP7_75t_L g4166 ( 
.A(n_3430),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_3874),
.B(n_3166),
.Y(n_4167)
);

AND2x4_ASAP7_75t_L g4168 ( 
.A(n_3576),
.B(n_2808),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3652),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_3608),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3654),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_SL g4172 ( 
.A(n_3911),
.B(n_2808),
.Y(n_4172)
);

BUFx6f_ASAP7_75t_L g4173 ( 
.A(n_3513),
.Y(n_4173)
);

INVx2_ASAP7_75t_SL g4174 ( 
.A(n_3523),
.Y(n_4174)
);

CKINVDCx20_ASAP7_75t_R g4175 ( 
.A(n_3918),
.Y(n_4175)
);

INVxp67_ASAP7_75t_SL g4176 ( 
.A(n_3532),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_3618),
.Y(n_4177)
);

BUFx6f_ASAP7_75t_L g4178 ( 
.A(n_3513),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_3620),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3659),
.Y(n_4180)
);

AND2x4_ASAP7_75t_L g4181 ( 
.A(n_3798),
.B(n_3482),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_3879),
.B(n_3168),
.Y(n_4182)
);

BUFx3_ASAP7_75t_L g4183 ( 
.A(n_3435),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3664),
.B(n_3131),
.Y(n_4184)
);

BUFx2_ASAP7_75t_L g4185 ( 
.A(n_3950),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3760),
.Y(n_4186)
);

NOR2xp33_ASAP7_75t_L g4187 ( 
.A(n_3823),
.B(n_3118),
.Y(n_4187)
);

NOR2xp33_ASAP7_75t_L g4188 ( 
.A(n_3901),
.B(n_3118),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_L g4189 ( 
.A(n_3545),
.B(n_3128),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_3638),
.Y(n_4190)
);

AOI22xp33_ASAP7_75t_SL g4191 ( 
.A1(n_3615),
.A2(n_3300),
.B1(n_3364),
.B2(n_3256),
.Y(n_4191)
);

AOI22xp33_ASAP7_75t_SL g4192 ( 
.A1(n_3635),
.A2(n_3364),
.B1(n_3300),
.B2(n_3136),
.Y(n_4192)
);

CKINVDCx8_ASAP7_75t_R g4193 ( 
.A(n_3833),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3769),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_3670),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_3743),
.Y(n_4196)
);

BUFx6f_ASAP7_75t_L g4197 ( 
.A(n_3550),
.Y(n_4197)
);

INVx5_ASAP7_75t_L g4198 ( 
.A(n_3549),
.Y(n_4198)
);

NOR2xp33_ASAP7_75t_R g4199 ( 
.A(n_3394),
.B(n_3364),
.Y(n_4199)
);

INVx1_ASAP7_75t_SL g4200 ( 
.A(n_3919),
.Y(n_4200)
);

INVx2_ASAP7_75t_SL g4201 ( 
.A(n_3758),
.Y(n_4201)
);

OR2x6_ASAP7_75t_L g4202 ( 
.A(n_3378),
.B(n_2921),
.Y(n_4202)
);

HB1xp67_ASAP7_75t_L g4203 ( 
.A(n_3512),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_3746),
.Y(n_4204)
);

INVx4_ASAP7_75t_L g4205 ( 
.A(n_3549),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3770),
.Y(n_4206)
);

BUFx3_ASAP7_75t_L g4207 ( 
.A(n_3484),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_3777),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_3759),
.Y(n_4209)
);

BUFx2_ASAP7_75t_L g4210 ( 
.A(n_3438),
.Y(n_4210)
);

BUFx3_ASAP7_75t_L g4211 ( 
.A(n_3906),
.Y(n_4211)
);

AOI22xp5_ASAP7_75t_L g4212 ( 
.A1(n_3766),
.A2(n_3136),
.B1(n_2749),
.B2(n_2734),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3803),
.Y(n_4213)
);

INVx5_ASAP7_75t_L g4214 ( 
.A(n_3549),
.Y(n_4214)
);

BUFx3_ASAP7_75t_L g4215 ( 
.A(n_3876),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_3811),
.Y(n_4216)
);

AND3x1_ASAP7_75t_L g4217 ( 
.A(n_3717),
.B(n_2907),
.C(n_2889),
.Y(n_4217)
);

NOR2x1p5_ASAP7_75t_L g4218 ( 
.A(n_3546),
.B(n_2921),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_3813),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_3947),
.B(n_194),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_SL g4221 ( 
.A(n_3453),
.B(n_3568),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_SL g4222 ( 
.A(n_3453),
.B(n_2808),
.Y(n_4222)
);

INVx2_ASAP7_75t_SL g4223 ( 
.A(n_3735),
.Y(n_4223)
);

BUFx2_ASAP7_75t_L g4224 ( 
.A(n_3689),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3816),
.Y(n_4225)
);

BUFx2_ASAP7_75t_L g4226 ( 
.A(n_3703),
.Y(n_4226)
);

INVx2_ASAP7_75t_SL g4227 ( 
.A(n_3518),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_3830),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_3843),
.Y(n_4229)
);

INVx1_ASAP7_75t_SL g4230 ( 
.A(n_3706),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3835),
.Y(n_4231)
);

OR2x6_ASAP7_75t_L g4232 ( 
.A(n_3477),
.B(n_2932),
.Y(n_4232)
);

INVx3_ASAP7_75t_L g4233 ( 
.A(n_3828),
.Y(n_4233)
);

BUFx6f_ASAP7_75t_L g4234 ( 
.A(n_3550),
.Y(n_4234)
);

AND2x6_ASAP7_75t_L g4235 ( 
.A(n_3453),
.B(n_2868),
.Y(n_4235)
);

OR2x6_ASAP7_75t_L g4236 ( 
.A(n_3749),
.B(n_2932),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_3864),
.Y(n_4237)
);

CKINVDCx5p33_ASAP7_75t_R g4238 ( 
.A(n_3882),
.Y(n_4238)
);

NAND3xp33_ASAP7_75t_SL g4239 ( 
.A(n_3739),
.B(n_3072),
.C(n_3027),
.Y(n_4239)
);

INVx1_ASAP7_75t_SL g4240 ( 
.A(n_3903),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_3921),
.Y(n_4241)
);

INVx1_ASAP7_75t_SL g4242 ( 
.A(n_3846),
.Y(n_4242)
);

AND2x4_ASAP7_75t_L g4243 ( 
.A(n_3482),
.B(n_2813),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_3838),
.Y(n_4244)
);

AOI22xp5_ASAP7_75t_L g4245 ( 
.A1(n_3773),
.A2(n_3136),
.B1(n_3170),
.B2(n_2907),
.Y(n_4245)
);

INVxp67_ASAP7_75t_SL g4246 ( 
.A(n_3598),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_3848),
.B(n_2855),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_3845),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_3854),
.Y(n_4249)
);

AOI211xp5_ASAP7_75t_L g4250 ( 
.A1(n_3617),
.A2(n_3175),
.B(n_2931),
.C(n_2889),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_3856),
.B(n_2856),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_3453),
.B(n_3568),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_3865),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_SL g4254 ( 
.A(n_3568),
.B(n_2813),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_SL g4255 ( 
.A(n_3568),
.B(n_2813),
.Y(n_4255)
);

OR2x2_ASAP7_75t_L g4256 ( 
.A(n_3808),
.B(n_2863),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_3910),
.Y(n_4257)
);

INVx2_ASAP7_75t_L g4258 ( 
.A(n_3924),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_3914),
.Y(n_4259)
);

AOI22xp33_ASAP7_75t_L g4260 ( 
.A1(n_3595),
.A2(n_3136),
.B1(n_3170),
.B2(n_2963),
.Y(n_4260)
);

NAND2xp5_ASAP7_75t_L g4261 ( 
.A(n_3783),
.B(n_3794),
.Y(n_4261)
);

INVx2_ASAP7_75t_L g4262 ( 
.A(n_3932),
.Y(n_4262)
);

NAND2x1p5_ASAP7_75t_L g4263 ( 
.A(n_3468),
.B(n_2829),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_SL g4264 ( 
.A(n_3568),
.B(n_2829),
.Y(n_4264)
);

AND2x4_ASAP7_75t_L g4265 ( 
.A(n_3488),
.B(n_2829),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_3805),
.B(n_2864),
.Y(n_4266)
);

HB1xp67_ASAP7_75t_L g4267 ( 
.A(n_3780),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3807),
.B(n_3926),
.Y(n_4268)
);

AND2x4_ASAP7_75t_L g4269 ( 
.A(n_3488),
.B(n_2838),
.Y(n_4269)
);

AND2x4_ASAP7_75t_SL g4270 ( 
.A(n_3518),
.B(n_3128),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_3949),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_3580),
.B(n_2878),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_3434),
.B(n_2887),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_SL g4274 ( 
.A(n_3509),
.B(n_2838),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_3747),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3748),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_3837),
.B(n_2897),
.Y(n_4277)
);

OAI22xp33_ASAP7_75t_L g4278 ( 
.A1(n_3403),
.A2(n_3142),
.B1(n_3138),
.B2(n_3176),
.Y(n_4278)
);

INVx3_ASAP7_75t_L g4279 ( 
.A(n_3828),
.Y(n_4279)
);

BUFx6f_ASAP7_75t_L g4280 ( 
.A(n_3550),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_3711),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_3751),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_L g4283 ( 
.A(n_3623),
.B(n_2904),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3757),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_3452),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_3462),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_3625),
.B(n_2906),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_3673),
.B(n_194),
.Y(n_4288)
);

INVx2_ASAP7_75t_L g4289 ( 
.A(n_3385),
.Y(n_4289)
);

BUFx3_ASAP7_75t_L g4290 ( 
.A(n_3605),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_SL g4291 ( 
.A(n_3509),
.B(n_2838),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_3928),
.B(n_2908),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_3814),
.B(n_2909),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_3495),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3520),
.Y(n_4295)
);

NOR2xp33_ASAP7_75t_L g4296 ( 
.A(n_3916),
.B(n_3138),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_3526),
.Y(n_4297)
);

AND2x4_ASAP7_75t_L g4298 ( 
.A(n_3922),
.B(n_2844),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_3390),
.Y(n_4299)
);

BUFx2_ASAP7_75t_L g4300 ( 
.A(n_3420),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_3527),
.Y(n_4301)
);

BUFx6f_ASAP7_75t_L g4302 ( 
.A(n_3690),
.Y(n_4302)
);

INVx2_ASAP7_75t_SL g4303 ( 
.A(n_3605),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_3529),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_3712),
.B(n_195),
.Y(n_4305)
);

HB1xp67_ASAP7_75t_L g4306 ( 
.A(n_3862),
.Y(n_4306)
);

AOI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_3948),
.A2(n_3170),
.B1(n_2931),
.B2(n_3142),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_3530),
.Y(n_4308)
);

OR2x2_ASAP7_75t_L g4309 ( 
.A(n_3809),
.B(n_2910),
.Y(n_4309)
);

INVx2_ASAP7_75t_SL g4310 ( 
.A(n_3655),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_3399),
.Y(n_4311)
);

OR2x4_ASAP7_75t_L g4312 ( 
.A(n_3558),
.B(n_3161),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_3401),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_3402),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_3421),
.Y(n_4315)
);

INVxp67_ASAP7_75t_L g4316 ( 
.A(n_3382),
.Y(n_4316)
);

AND2x4_ASAP7_75t_L g4317 ( 
.A(n_3420),
.B(n_2844),
.Y(n_4317)
);

BUFx3_ASAP7_75t_L g4318 ( 
.A(n_3655),
.Y(n_4318)
);

INVx1_ASAP7_75t_SL g4319 ( 
.A(n_3676),
.Y(n_4319)
);

AOI22xp5_ASAP7_75t_L g4320 ( 
.A1(n_3601),
.A2(n_3173),
.B1(n_3145),
.B2(n_3149),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3531),
.Y(n_4321)
);

INVx2_ASAP7_75t_SL g4322 ( 
.A(n_3676),
.Y(n_4322)
);

NOR3xp33_ASAP7_75t_L g4323 ( 
.A(n_3647),
.B(n_3176),
.C(n_3159),
.Y(n_4323)
);

INVx3_ASAP7_75t_L g4324 ( 
.A(n_3690),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_SL g4325 ( 
.A(n_3899),
.B(n_2844),
.Y(n_4325)
);

BUFx2_ASAP7_75t_SL g4326 ( 
.A(n_3549),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_3539),
.Y(n_4327)
);

NOR2xp33_ASAP7_75t_L g4328 ( 
.A(n_3537),
.B(n_3159),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_3386),
.B(n_2912),
.Y(n_4329)
);

BUFx3_ASAP7_75t_L g4330 ( 
.A(n_3690),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_3406),
.B(n_3141),
.Y(n_4331)
);

INVx3_ASAP7_75t_L g4332 ( 
.A(n_3723),
.Y(n_4332)
);

AND2x4_ASAP7_75t_L g4333 ( 
.A(n_3622),
.B(n_2867),
.Y(n_4333)
);

INVx2_ASAP7_75t_L g4334 ( 
.A(n_3422),
.Y(n_4334)
);

BUFx12f_ASAP7_75t_L g4335 ( 
.A(n_3920),
.Y(n_4335)
);

INVx1_ASAP7_75t_SL g4336 ( 
.A(n_3727),
.Y(n_4336)
);

HB1xp67_ASAP7_75t_L g4337 ( 
.A(n_3872),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_3409),
.B(n_3157),
.Y(n_4338)
);

BUFx6f_ASAP7_75t_L g4339 ( 
.A(n_3723),
.Y(n_4339)
);

BUFx6f_ASAP7_75t_L g4340 ( 
.A(n_3723),
.Y(n_4340)
);

BUFx3_ASAP7_75t_L g4341 ( 
.A(n_3849),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_3627),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_3632),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_3542),
.Y(n_4344)
);

AOI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_3502),
.A2(n_3589),
.B1(n_3554),
.B2(n_3729),
.Y(n_4345)
);

AOI22xp33_ASAP7_75t_L g4346 ( 
.A1(n_3653),
.A2(n_2888),
.B1(n_3162),
.B2(n_2922),
.Y(n_4346)
);

INVxp67_ASAP7_75t_L g4347 ( 
.A(n_3528),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_3750),
.B(n_2867),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_3414),
.B(n_2916),
.Y(n_4349)
);

AOI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_3789),
.A2(n_2924),
.B1(n_2947),
.B2(n_3161),
.Y(n_4350)
);

AOI22xp33_ASAP7_75t_L g4351 ( 
.A1(n_3552),
.A2(n_3592),
.B1(n_3792),
.B2(n_3913),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_3547),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_3418),
.B(n_195),
.Y(n_4353)
);

NOR2xp33_ASAP7_75t_L g4354 ( 
.A(n_3551),
.B(n_2920),
.Y(n_4354)
);

INVx2_ASAP7_75t_SL g4355 ( 
.A(n_3450),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_3636),
.Y(n_4356)
);

INVxp67_ASAP7_75t_SL g4357 ( 
.A(n_3737),
.Y(n_4357)
);

OAI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_3940),
.A2(n_3165),
.B(n_3164),
.Y(n_4358)
);

OAI22xp33_ASAP7_75t_L g4359 ( 
.A1(n_3541),
.A2(n_3586),
.B1(n_3587),
.B2(n_3581),
.Y(n_4359)
);

NOR2xp33_ASAP7_75t_L g4360 ( 
.A(n_3613),
.B(n_3161),
.Y(n_4360)
);

HB1xp67_ASAP7_75t_L g4361 ( 
.A(n_3444),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_3565),
.Y(n_4362)
);

BUFx6f_ASAP7_75t_L g4363 ( 
.A(n_3849),
.Y(n_4363)
);

BUFx6f_ASAP7_75t_L g4364 ( 
.A(n_3849),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_SL g4365 ( 
.A(n_3930),
.B(n_2867),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_3567),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_3611),
.B(n_196),
.Y(n_4367)
);

BUFx12f_ASAP7_75t_L g4368 ( 
.A(n_3861),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_3642),
.Y(n_4369)
);

INVx4_ASAP7_75t_L g4370 ( 
.A(n_3861),
.Y(n_4370)
);

BUFx3_ASAP7_75t_L g4371 ( 
.A(n_3861),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_3649),
.Y(n_4372)
);

OR2x2_ASAP7_75t_SL g4373 ( 
.A(n_3941),
.B(n_3177),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_3839),
.B(n_196),
.Y(n_4374)
);

OR2x2_ASAP7_75t_L g4375 ( 
.A(n_3818),
.B(n_2806),
.Y(n_4375)
);

BUFx3_ASAP7_75t_L g4376 ( 
.A(n_3887),
.Y(n_4376)
);

NOR2xp33_ASAP7_75t_L g4377 ( 
.A(n_3616),
.B(n_3163),
.Y(n_4377)
);

BUFx2_ASAP7_75t_L g4378 ( 
.A(n_3933),
.Y(n_4378)
);

INVx3_ASAP7_75t_L g4379 ( 
.A(n_3887),
.Y(n_4379)
);

INVx2_ASAP7_75t_L g4380 ( 
.A(n_3658),
.Y(n_4380)
);

INVx5_ASAP7_75t_L g4381 ( 
.A(n_3887),
.Y(n_4381)
);

BUFx2_ASAP7_75t_L g4382 ( 
.A(n_3933),
.Y(n_4382)
);

BUFx6f_ASAP7_75t_L g4383 ( 
.A(n_3939),
.Y(n_4383)
);

AOI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_3671),
.A2(n_3163),
.B1(n_3172),
.B2(n_3160),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_3573),
.Y(n_4385)
);

HB1xp67_ASAP7_75t_L g4386 ( 
.A(n_3449),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_3593),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_3603),
.Y(n_4388)
);

INVx3_ASAP7_75t_L g4389 ( 
.A(n_3797),
.Y(n_4389)
);

HB1xp67_ASAP7_75t_L g4390 ( 
.A(n_3870),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_3894),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_3895),
.Y(n_4392)
);

CKINVDCx5p33_ASAP7_75t_R g4393 ( 
.A(n_3767),
.Y(n_4393)
);

INVxp67_ASAP7_75t_SL g4394 ( 
.A(n_3768),
.Y(n_4394)
);

AND2x4_ASAP7_75t_L g4395 ( 
.A(n_3645),
.B(n_3177),
.Y(n_4395)
);

AND2x4_ASAP7_75t_SL g4396 ( 
.A(n_3939),
.B(n_3341),
.Y(n_4396)
);

INVx2_ASAP7_75t_SL g4397 ( 
.A(n_3912),
.Y(n_4397)
);

AND2x2_ASAP7_75t_L g4398 ( 
.A(n_3667),
.B(n_197),
.Y(n_4398)
);

AND2x2_ASAP7_75t_SL g4399 ( 
.A(n_3667),
.B(n_3177),
.Y(n_4399)
);

INVx2_ASAP7_75t_L g4400 ( 
.A(n_3662),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_3663),
.Y(n_4401)
);

INVx2_ASAP7_75t_SL g4402 ( 
.A(n_3917),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_3893),
.Y(n_4403)
);

HB1xp67_ASAP7_75t_L g4404 ( 
.A(n_3871),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_3897),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_3778),
.B(n_197),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_3464),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_3681),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_3682),
.Y(n_4409)
);

BUFx2_ASAP7_75t_L g4410 ( 
.A(n_3668),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_3470),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_3480),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_SL g4413 ( 
.A(n_3562),
.B(n_3178),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_3487),
.Y(n_4414)
);

AOI21xp33_ASAP7_75t_L g4415 ( 
.A1(n_3836),
.A2(n_2810),
.B(n_3163),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_3867),
.B(n_198),
.Y(n_4416)
);

NAND2x1p5_ASAP7_75t_L g4417 ( 
.A(n_3675),
.B(n_3178),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_3490),
.Y(n_4418)
);

CKINVDCx5p33_ASAP7_75t_R g4419 ( 
.A(n_3524),
.Y(n_4419)
);

INVxp67_ASAP7_75t_SL g4420 ( 
.A(n_3905),
.Y(n_4420)
);

NAND2x2_ASAP7_75t_L g4421 ( 
.A(n_3381),
.B(n_198),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_3686),
.Y(n_4422)
);

AOI22xp33_ASAP7_75t_L g4423 ( 
.A1(n_3695),
.A2(n_3172),
.B1(n_3160),
.B2(n_2828),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_3492),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_3694),
.Y(n_4425)
);

BUFx12f_ASAP7_75t_L g4426 ( 
.A(n_3612),
.Y(n_4426)
);

INVx3_ASAP7_75t_SL g4427 ( 
.A(n_3720),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_3869),
.B(n_198),
.Y(n_4428)
);

CKINVDCx20_ASAP7_75t_R g4429 ( 
.A(n_3431),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_3693),
.B(n_199),
.Y(n_4430)
);

BUFx4f_ASAP7_75t_L g4431 ( 
.A(n_3724),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_3824),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_3697),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_3831),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_3819),
.Y(n_4435)
);

AND2x4_ASAP7_75t_L g4436 ( 
.A(n_3698),
.B(n_3178),
.Y(n_4436)
);

OR2x2_ASAP7_75t_L g4437 ( 
.A(n_3765),
.B(n_3277),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_3699),
.Y(n_4438)
);

AND2x4_ASAP7_75t_L g4439 ( 
.A(n_3707),
.B(n_3185),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_3709),
.Y(n_4440)
);

INVxp67_ASAP7_75t_SL g4441 ( 
.A(n_3931),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_3713),
.Y(n_4442)
);

OR2x2_ASAP7_75t_L g4443 ( 
.A(n_3771),
.B(n_3277),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_3715),
.Y(n_4444)
);

INVxp67_ASAP7_75t_L g4445 ( 
.A(n_3510),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_3820),
.B(n_199),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_3857),
.B(n_199),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_3732),
.Y(n_4448)
);

INVx3_ASAP7_75t_L g4449 ( 
.A(n_3734),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_3738),
.Y(n_4450)
);

BUFx6f_ASAP7_75t_L g4451 ( 
.A(n_3384),
.Y(n_4451)
);

AOI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_3742),
.A2(n_3172),
.B1(n_2828),
.B2(n_2830),
.Y(n_4452)
);

INVx1_ASAP7_75t_SL g4453 ( 
.A(n_3934),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_3648),
.Y(n_4454)
);

OR2x2_ASAP7_75t_L g4455 ( 
.A(n_3779),
.B(n_3303),
.Y(n_4455)
);

AOI22xp5_ASAP7_75t_L g4456 ( 
.A1(n_3754),
.A2(n_2830),
.B1(n_3199),
.B2(n_2806),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_3858),
.B(n_200),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_3859),
.B(n_200),
.Y(n_4458)
);

AND2x6_ASAP7_75t_SL g4459 ( 
.A(n_3465),
.B(n_201),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_3784),
.Y(n_4460)
);

INVx1_ASAP7_75t_SL g4461 ( 
.A(n_3935),
.Y(n_4461)
);

NOR2xp33_ASAP7_75t_L g4462 ( 
.A(n_3822),
.B(n_201),
.Y(n_4462)
);

BUFx2_ASAP7_75t_L g4463 ( 
.A(n_3853),
.Y(n_4463)
);

INVx2_ASAP7_75t_L g4464 ( 
.A(n_3661),
.Y(n_4464)
);

INVx3_ASAP7_75t_L g4465 ( 
.A(n_3944),
.Y(n_4465)
);

INVx2_ASAP7_75t_SL g4466 ( 
.A(n_3785),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_3863),
.B(n_201),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_3786),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_3891),
.Y(n_4469)
);

INVx1_ASAP7_75t_SL g4470 ( 
.A(n_3907),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_SL g4471 ( 
.A(n_3782),
.B(n_3185),
.Y(n_4471)
);

AOI22xp33_ASAP7_75t_L g4472 ( 
.A1(n_3722),
.A2(n_3339),
.B1(n_3199),
.B2(n_3226),
.Y(n_4472)
);

AOI22xp33_ASAP7_75t_L g4473 ( 
.A1(n_3761),
.A2(n_3207),
.B1(n_3290),
.B2(n_3226),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_3788),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_3840),
.B(n_202),
.Y(n_4475)
);

AOI22xp33_ASAP7_75t_L g4476 ( 
.A1(n_3883),
.A2(n_3207),
.B1(n_3290),
.B2(n_3249),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_L g4477 ( 
.A(n_3841),
.B(n_202),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_3844),
.B(n_202),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_3762),
.B(n_203),
.Y(n_4479)
);

AOI22xp33_ASAP7_75t_L g4480 ( 
.A1(n_3776),
.A2(n_3324),
.B1(n_3339),
.B2(n_3249),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_3790),
.Y(n_4481)
);

INVxp67_ASAP7_75t_L g4482 ( 
.A(n_3756),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_3936),
.B(n_203),
.Y(n_4483)
);

BUFx3_ASAP7_75t_L g4484 ( 
.A(n_3801),
.Y(n_4484)
);

NOR2x1p5_ASAP7_75t_L g4485 ( 
.A(n_3802),
.B(n_3303),
.Y(n_4485)
);

CKINVDCx5p33_ASAP7_75t_R g4486 ( 
.A(n_3507),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_3938),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_3599),
.B(n_204),
.Y(n_4488)
);

INVx4_ASAP7_75t_L g4489 ( 
.A(n_3515),
.Y(n_4489)
);

INVx1_ASAP7_75t_SL g4490 ( 
.A(n_3812),
.Y(n_4490)
);

BUFx2_ASAP7_75t_L g4491 ( 
.A(n_3880),
.Y(n_4491)
);

CKINVDCx5p33_ASAP7_75t_R g4492 ( 
.A(n_3559),
.Y(n_4492)
);

AND2x4_ASAP7_75t_L g4493 ( 
.A(n_3817),
.B(n_3185),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_3467),
.Y(n_4494)
);

AND2x4_ASAP7_75t_L g4495 ( 
.A(n_3860),
.B(n_3227),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_3497),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_3494),
.Y(n_4497)
);

A2O1A1Ixp33_ASAP7_75t_L g4498 ( 
.A1(n_3407),
.A2(n_3324),
.B(n_3230),
.C(n_3243),
.Y(n_4498)
);

BUFx6f_ASAP7_75t_L g4499 ( 
.A(n_3457),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_3597),
.Y(n_4500)
);

OR2x6_ASAP7_75t_L g4501 ( 
.A(n_3877),
.B(n_3878),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_3890),
.B(n_204),
.Y(n_4502)
);

INVx2_ASAP7_75t_SL g4503 ( 
.A(n_3881),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_3463),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_3674),
.B(n_204),
.Y(n_4505)
);

INVx2_ASAP7_75t_SL g4506 ( 
.A(n_3885),
.Y(n_4506)
);

A2O1A1Ixp33_ASAP7_75t_L g4507 ( 
.A1(n_3478),
.A2(n_3744),
.B(n_3624),
.C(n_3432),
.Y(n_4507)
);

INVxp67_ASAP7_75t_SL g4508 ( 
.A(n_3796),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_3504),
.B(n_205),
.Y(n_4509)
);

AND2x4_ASAP7_75t_L g4510 ( 
.A(n_3892),
.B(n_3227),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_3644),
.Y(n_4511)
);

OR2x2_ASAP7_75t_L g4512 ( 
.A(n_3677),
.B(n_205),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_3714),
.B(n_206),
.Y(n_4513)
);

OR2x6_ASAP7_75t_L g4514 ( 
.A(n_3966),
.B(n_3451),
.Y(n_4514)
);

BUFx3_ASAP7_75t_L g4515 ( 
.A(n_4076),
.Y(n_4515)
);

O2A1O1Ixp33_ASAP7_75t_SL g4516 ( 
.A1(n_3952),
.A2(n_3804),
.B(n_3898),
.C(n_3514),
.Y(n_4516)
);

O2A1O1Ixp33_ASAP7_75t_SL g4517 ( 
.A1(n_4200),
.A2(n_4336),
.B(n_4045),
.C(n_4397),
.Y(n_4517)
);

AOI21xp5_ASAP7_75t_L g4518 ( 
.A1(n_4358),
.A2(n_4172),
.B(n_4176),
.Y(n_4518)
);

O2A1O1Ixp5_ASAP7_75t_L g4519 ( 
.A1(n_4431),
.A2(n_3621),
.B(n_3666),
.C(n_3619),
.Y(n_4519)
);

OAI22xp5_ASAP7_75t_L g4520 ( 
.A1(n_4016),
.A2(n_3688),
.B1(n_3656),
.B2(n_3536),
.Y(n_4520)
);

OAI22xp5_ASAP7_75t_SL g4521 ( 
.A1(n_3988),
.A2(n_3902),
.B1(n_3691),
.B2(n_3672),
.Y(n_4521)
);

HB1xp67_ASAP7_75t_L g4522 ( 
.A(n_4039),
.Y(n_4522)
);

NOR2xp33_ASAP7_75t_L g4523 ( 
.A(n_4193),
.B(n_3413),
.Y(n_4523)
);

AOI22xp33_ASAP7_75t_L g4524 ( 
.A1(n_4426),
.A2(n_3781),
.B1(n_3945),
.B2(n_3415),
.Y(n_4524)
);

NOR2xp33_ASAP7_75t_L g4525 ( 
.A(n_4078),
.B(n_3424),
.Y(n_4525)
);

NAND3xp33_ASAP7_75t_SL g4526 ( 
.A(n_4175),
.B(n_3433),
.C(n_3815),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_4246),
.A2(n_3024),
.B(n_2868),
.Y(n_4527)
);

AO21x1_ASAP7_75t_L g4528 ( 
.A1(n_4005),
.A2(n_3800),
.B(n_3799),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_4080),
.B(n_3850),
.Y(n_4529)
);

A2O1A1Ixp33_ASAP7_75t_L g4530 ( 
.A1(n_4431),
.A2(n_3579),
.B(n_3519),
.C(n_3506),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_SL g4531 ( 
.A(n_4022),
.B(n_3227),
.Y(n_4531)
);

AOI21xp5_ASAP7_75t_L g4532 ( 
.A1(n_4357),
.A2(n_3026),
.B(n_2929),
.Y(n_4532)
);

NOR2xp33_ASAP7_75t_L g4533 ( 
.A(n_4419),
.B(n_3500),
.Y(n_4533)
);

AND2x2_ASAP7_75t_SL g4534 ( 
.A(n_4163),
.B(n_3763),
.Y(n_4534)
);

OR2x6_ASAP7_75t_L g4535 ( 
.A(n_3966),
.B(n_3810),
.Y(n_4535)
);

AOI21xp5_ASAP7_75t_L g4536 ( 
.A1(n_4394),
.A2(n_3026),
.B(n_2929),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4084),
.B(n_3946),
.Y(n_4537)
);

NOR2xp33_ASAP7_75t_L g4538 ( 
.A(n_3955),
.B(n_3572),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4077),
.Y(n_4539)
);

AOI21xp5_ASAP7_75t_L g4540 ( 
.A1(n_4420),
.A2(n_3026),
.B(n_2929),
.Y(n_4540)
);

NOR2xp33_ASAP7_75t_L g4541 ( 
.A(n_4335),
.B(n_3741),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4085),
.B(n_3772),
.Y(n_4542)
);

NOR2xp33_ASAP7_75t_R g4543 ( 
.A(n_4090),
.B(n_3230),
.Y(n_4543)
);

O2A1O1Ixp5_ASAP7_75t_L g4544 ( 
.A1(n_4205),
.A2(n_3669),
.B(n_3485),
.C(n_3475),
.Y(n_4544)
);

A2O1A1Ixp33_ASAP7_75t_L g4545 ( 
.A1(n_4163),
.A2(n_3643),
.B(n_3425),
.C(n_3543),
.Y(n_4545)
);

INVx3_ASAP7_75t_SL g4546 ( 
.A(n_4052),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_3954),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4230),
.B(n_3791),
.Y(n_4548)
);

BUFx2_ASAP7_75t_L g4549 ( 
.A(n_4368),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_4056),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_3962),
.Y(n_4551)
);

BUFx2_ASAP7_75t_L g4552 ( 
.A(n_3994),
.Y(n_4552)
);

NOR3xp33_ASAP7_75t_SL g4553 ( 
.A(n_4051),
.B(n_4107),
.C(n_4154),
.Y(n_4553)
);

BUFx3_ASAP7_75t_L g4554 ( 
.A(n_4013),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4127),
.B(n_3847),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_L g4556 ( 
.A(n_4133),
.B(n_4281),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_4068),
.Y(n_4557)
);

OAI22xp5_ASAP7_75t_SL g4558 ( 
.A1(n_4091),
.A2(n_3875),
.B1(n_3884),
.B2(n_3392),
.Y(n_4558)
);

O2A1O1Ixp33_ASAP7_75t_L g4559 ( 
.A1(n_3976),
.A2(n_3609),
.B(n_3570),
.C(n_3574),
.Y(n_4559)
);

AOI22xp33_ASAP7_75t_L g4560 ( 
.A1(n_4010),
.A2(n_3583),
.B1(n_3533),
.B2(n_3591),
.Y(n_4560)
);

INVx2_ASAP7_75t_L g4561 ( 
.A(n_4075),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_4288),
.B(n_206),
.Y(n_4562)
);

BUFx3_ASAP7_75t_L g4563 ( 
.A(n_4015),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_SL g4564 ( 
.A(n_4022),
.B(n_3230),
.Y(n_4564)
);

INVxp67_ASAP7_75t_L g4565 ( 
.A(n_4065),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_3964),
.Y(n_4566)
);

INVx1_ASAP7_75t_SL g4567 ( 
.A(n_3965),
.Y(n_4567)
);

A2O1A1Ixp33_ASAP7_75t_L g4568 ( 
.A1(n_4250),
.A2(n_4036),
.B(n_4050),
.C(n_4103),
.Y(n_4568)
);

OAI22xp5_ASAP7_75t_L g4569 ( 
.A1(n_4022),
.A2(n_3795),
.B1(n_3278),
.B2(n_3295),
.Y(n_4569)
);

BUFx2_ASAP7_75t_L g4570 ( 
.A(n_4290),
.Y(n_4570)
);

NAND3xp33_ASAP7_75t_L g4571 ( 
.A(n_4462),
.B(n_3389),
.C(n_3380),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_L g4572 ( 
.A(n_4133),
.B(n_206),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_4096),
.A2(n_2938),
.B(n_2936),
.Y(n_4573)
);

CKINVDCx14_ASAP7_75t_R g4574 ( 
.A(n_3974),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_L g4575 ( 
.A(n_4147),
.B(n_207),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_SL g4576 ( 
.A(n_3998),
.B(n_3243),
.Y(n_4576)
);

OAI22xp5_ASAP7_75t_L g4577 ( 
.A1(n_4429),
.A2(n_3278),
.B1(n_3295),
.B2(n_3243),
.Y(n_4577)
);

INVx2_ASAP7_75t_L g4578 ( 
.A(n_4083),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_3985),
.Y(n_4579)
);

OAI321xp33_ASAP7_75t_L g4580 ( 
.A1(n_4359),
.A2(n_3295),
.A3(n_3317),
.B1(n_3341),
.B2(n_3322),
.C(n_3278),
.Y(n_4580)
);

AO21x1_ASAP7_75t_L g4581 ( 
.A1(n_4205),
.A2(n_208),
.B(n_209),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_SL g4582 ( 
.A(n_3998),
.B(n_3317),
.Y(n_4582)
);

BUFx2_ASAP7_75t_L g4583 ( 
.A(n_4318),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_SL g4584 ( 
.A(n_3998),
.B(n_3317),
.Y(n_4584)
);

AOI21xp5_ASAP7_75t_L g4585 ( 
.A1(n_4274),
.A2(n_2938),
.B(n_2936),
.Y(n_4585)
);

INVx4_ASAP7_75t_L g4586 ( 
.A(n_4004),
.Y(n_4586)
);

O2A1O1Ixp5_ASAP7_75t_SL g4587 ( 
.A1(n_4291),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_4587)
);

O2A1O1Ixp33_ASAP7_75t_L g4588 ( 
.A1(n_4482),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4305),
.B(n_211),
.Y(n_4589)
);

NOR2xp33_ASAP7_75t_L g4590 ( 
.A(n_4238),
.B(n_211),
.Y(n_4590)
);

NOR2xp33_ASAP7_75t_L g4591 ( 
.A(n_4098),
.B(n_4393),
.Y(n_4591)
);

BUFx2_ASAP7_75t_SL g4592 ( 
.A(n_3968),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_SL g4593 ( 
.A(n_4198),
.B(n_3322),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4220),
.B(n_212),
.Y(n_4594)
);

BUFx3_ASAP7_75t_L g4595 ( 
.A(n_4026),
.Y(n_4595)
);

CKINVDCx20_ASAP7_75t_R g4596 ( 
.A(n_4017),
.Y(n_4596)
);

AOI21xp5_ASAP7_75t_L g4597 ( 
.A1(n_4498),
.A2(n_2938),
.B(n_2936),
.Y(n_4597)
);

AOI21xp5_ASAP7_75t_L g4598 ( 
.A1(n_4059),
.A2(n_2954),
.B(n_2940),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_3992),
.Y(n_4599)
);

NOR2xp33_ASAP7_75t_L g4600 ( 
.A(n_4347),
.B(n_212),
.Y(n_4600)
);

NOR3xp33_ASAP7_75t_L g4601 ( 
.A(n_4031),
.B(n_220),
.C(n_212),
.Y(n_4601)
);

INVx5_ASAP7_75t_L g4602 ( 
.A(n_4064),
.Y(n_4602)
);

BUFx3_ASAP7_75t_L g4603 ( 
.A(n_4099),
.Y(n_4603)
);

O2A1O1Ixp33_ASAP7_75t_L g4604 ( 
.A1(n_4261),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4267),
.B(n_213),
.Y(n_4605)
);

CKINVDCx8_ASAP7_75t_R g4606 ( 
.A(n_4073),
.Y(n_4606)
);

A2O1A1Ixp33_ASAP7_75t_L g4607 ( 
.A1(n_4270),
.A2(n_3341),
.B(n_3348),
.C(n_3322),
.Y(n_4607)
);

BUFx3_ASAP7_75t_L g4608 ( 
.A(n_3963),
.Y(n_4608)
);

AOI21x1_ASAP7_75t_L g4609 ( 
.A1(n_4059),
.A2(n_2954),
.B(n_2940),
.Y(n_4609)
);

NOR2xp33_ASAP7_75t_L g4610 ( 
.A(n_4223),
.B(n_213),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4092),
.Y(n_4611)
);

HB1xp67_ASAP7_75t_L g4612 ( 
.A(n_4067),
.Y(n_4612)
);

O2A1O1Ixp33_ASAP7_75t_L g4613 ( 
.A1(n_4268),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_L g4614 ( 
.A(n_4088),
.B(n_214),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_4435),
.B(n_215),
.Y(n_4615)
);

OR2x6_ASAP7_75t_SL g4616 ( 
.A(n_4486),
.B(n_216),
.Y(n_4616)
);

OAI22xp5_ASAP7_75t_L g4617 ( 
.A1(n_3956),
.A2(n_3348),
.B1(n_3350),
.B2(n_2954),
.Y(n_4617)
);

AOI21xp5_ASAP7_75t_L g4618 ( 
.A1(n_4254),
.A2(n_2986),
.B(n_2974),
.Y(n_4618)
);

A2O1A1Ixp33_ASAP7_75t_L g4619 ( 
.A1(n_4507),
.A2(n_3350),
.B(n_3348),
.C(n_2974),
.Y(n_4619)
);

INVx2_ASAP7_75t_L g4620 ( 
.A(n_4093),
.Y(n_4620)
);

INVxp67_ASAP7_75t_L g4621 ( 
.A(n_4185),
.Y(n_4621)
);

NOR2xp33_ASAP7_75t_L g4622 ( 
.A(n_4008),
.B(n_216),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_L g4623 ( 
.A(n_4432),
.B(n_217),
.Y(n_4623)
);

O2A1O1Ixp33_ASAP7_75t_L g4624 ( 
.A1(n_4182),
.A2(n_219),
.B(n_217),
.C(n_218),
.Y(n_4624)
);

BUFx3_ASAP7_75t_L g4625 ( 
.A(n_3983),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_3996),
.Y(n_4626)
);

AOI22xp33_ASAP7_75t_L g4627 ( 
.A1(n_4494),
.A2(n_3350),
.B1(n_3127),
.B2(n_3116),
.Y(n_4627)
);

AND2x6_ASAP7_75t_SL g4628 ( 
.A(n_4064),
.B(n_217),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4434),
.B(n_219),
.Y(n_4629)
);

O2A1O1Ixp33_ASAP7_75t_SL g4630 ( 
.A1(n_4174),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_4630)
);

BUFx3_ASAP7_75t_L g4631 ( 
.A(n_3990),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4460),
.B(n_220),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4001),
.Y(n_4633)
);

AO22x1_ASAP7_75t_L g4634 ( 
.A1(n_4181),
.A2(n_2974),
.B1(n_2986),
.B2(n_2940),
.Y(n_4634)
);

OAI22xp5_ASAP7_75t_L g4635 ( 
.A1(n_4421),
.A2(n_3024),
.B1(n_3061),
.B2(n_2986),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4468),
.B(n_221),
.Y(n_4636)
);

NOR2xp33_ASAP7_75t_R g4637 ( 
.A(n_3973),
.B(n_222),
.Y(n_4637)
);

HB1xp67_ASAP7_75t_L g4638 ( 
.A(n_4306),
.Y(n_4638)
);

NOR3xp33_ASAP7_75t_L g4639 ( 
.A(n_4081),
.B(n_230),
.C(n_222),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_SL g4640 ( 
.A(n_4198),
.B(n_3070),
.Y(n_4640)
);

A2O1A1Ixp33_ASAP7_75t_L g4641 ( 
.A1(n_4058),
.A2(n_3061),
.B(n_3070),
.C(n_3024),
.Y(n_4641)
);

BUFx3_ASAP7_75t_L g4642 ( 
.A(n_3982),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4115),
.B(n_223),
.Y(n_4643)
);

NAND3xp33_ASAP7_75t_SL g4644 ( 
.A(n_4129),
.B(n_223),
.C(n_224),
.Y(n_4644)
);

INVx1_ASAP7_75t_SL g4645 ( 
.A(n_4100),
.Y(n_4645)
);

AOI21xp5_ASAP7_75t_L g4646 ( 
.A1(n_4255),
.A2(n_3070),
.B(n_3061),
.Y(n_4646)
);

A2O1A1Ixp33_ASAP7_75t_L g4647 ( 
.A1(n_4006),
.A2(n_3127),
.B(n_3116),
.C(n_225),
.Y(n_4647)
);

AOI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4264),
.A2(n_3127),
.B(n_3116),
.Y(n_4648)
);

AND2x2_ASAP7_75t_SL g4649 ( 
.A(n_4399),
.B(n_223),
.Y(n_4649)
);

OAI22xp5_ASAP7_75t_L g4650 ( 
.A1(n_4492),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4474),
.B(n_224),
.Y(n_4651)
);

NOR2xp33_ASAP7_75t_L g4652 ( 
.A(n_4445),
.B(n_226),
.Y(n_4652)
);

BUFx3_ASAP7_75t_L g4653 ( 
.A(n_4014),
.Y(n_4653)
);

OAI21x1_ASAP7_75t_L g4654 ( 
.A1(n_4221),
.A2(n_867),
.B(n_859),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4012),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_SL g4656 ( 
.A(n_4198),
.B(n_227),
.Y(n_4656)
);

OAI21xp33_ASAP7_75t_L g4657 ( 
.A1(n_4345),
.A2(n_227),
.B(n_228),
.Y(n_4657)
);

NAND2xp5_ASAP7_75t_L g4658 ( 
.A(n_4481),
.B(n_4023),
.Y(n_4658)
);

NOR2xp33_ASAP7_75t_L g4659 ( 
.A(n_4009),
.B(n_227),
.Y(n_4659)
);

BUFx6f_ASAP7_75t_L g4660 ( 
.A(n_4018),
.Y(n_4660)
);

INVx3_ASAP7_75t_L g4661 ( 
.A(n_4181),
.Y(n_4661)
);

O2A1O1Ixp33_ASAP7_75t_L g4662 ( 
.A1(n_4130),
.A2(n_231),
.B(n_228),
.C(n_229),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4028),
.B(n_229),
.Y(n_4663)
);

OAI21x1_ASAP7_75t_L g4664 ( 
.A1(n_4252),
.A2(n_870),
.B(n_861),
.Y(n_4664)
);

CKINVDCx5p33_ASAP7_75t_R g4665 ( 
.A(n_4066),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_4117),
.Y(n_4666)
);

OAI22xp5_ASAP7_75t_L g4667 ( 
.A1(n_4232),
.A2(n_232),
.B1(n_229),
.B2(n_231),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4032),
.B(n_231),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4121),
.Y(n_4669)
);

AO21x2_ASAP7_75t_L g4670 ( 
.A1(n_4070),
.A2(n_232),
.B(n_233),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4033),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_SL g4672 ( 
.A(n_4214),
.B(n_232),
.Y(n_4672)
);

NOR2xp33_ASAP7_75t_L g4673 ( 
.A(n_4131),
.B(n_233),
.Y(n_4673)
);

AND2x4_ASAP7_75t_L g4674 ( 
.A(n_4214),
.B(n_233),
.Y(n_4674)
);

INVx4_ASAP7_75t_L g4675 ( 
.A(n_4004),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_SL g4676 ( 
.A(n_4214),
.B(n_234),
.Y(n_4676)
);

AOI22xp5_ASAP7_75t_L g4677 ( 
.A1(n_4497),
.A2(n_4500),
.B1(n_4511),
.B2(n_4316),
.Y(n_4677)
);

INVx2_ASAP7_75t_L g4678 ( 
.A(n_4137),
.Y(n_4678)
);

OAI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4232),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_4679)
);

BUFx12f_ASAP7_75t_L g4680 ( 
.A(n_3967),
.Y(n_4680)
);

BUFx8_ASAP7_75t_L g4681 ( 
.A(n_3981),
.Y(n_4681)
);

INVx2_ASAP7_75t_L g4682 ( 
.A(n_4140),
.Y(n_4682)
);

A2O1A1Ixp33_ASAP7_75t_L g4683 ( 
.A1(n_4118),
.A2(n_237),
.B(n_234),
.C(n_235),
.Y(n_4683)
);

OAI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_3960),
.A2(n_238),
.B1(n_235),
.B2(n_237),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_4034),
.B(n_237),
.Y(n_4685)
);

INVx4_ASAP7_75t_L g4686 ( 
.A(n_4004),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4035),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4042),
.B(n_238),
.Y(n_4688)
);

O2A1O1Ixp33_ASAP7_75t_L g4689 ( 
.A1(n_4367),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4142),
.Y(n_4690)
);

AOI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4124),
.A2(n_4325),
.B(n_4222),
.Y(n_4691)
);

O2A1O1Ixp33_ASAP7_75t_L g4692 ( 
.A1(n_4483),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4044),
.B(n_241),
.Y(n_4693)
);

AO21x1_ASAP7_75t_L g4694 ( 
.A1(n_4489),
.A2(n_241),
.B(n_242),
.Y(n_4694)
);

AOI21xp5_ASAP7_75t_L g4695 ( 
.A1(n_4454),
.A2(n_243),
.B(n_244),
.Y(n_4695)
);

AOI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4464),
.A2(n_243),
.B(n_244),
.Y(n_4696)
);

AND2x4_ASAP7_75t_L g4697 ( 
.A(n_4217),
.B(n_244),
.Y(n_4697)
);

NOR2xp33_ASAP7_75t_L g4698 ( 
.A(n_4119),
.B(n_245),
.Y(n_4698)
);

INVxp67_ASAP7_75t_SL g4699 ( 
.A(n_4203),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_SL g4700 ( 
.A(n_4020),
.B(n_4489),
.Y(n_4700)
);

AOI22xp5_ASAP7_75t_L g4701 ( 
.A1(n_4508),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_4701)
);

HB1xp67_ASAP7_75t_L g4702 ( 
.A(n_4242),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4053),
.B(n_245),
.Y(n_4703)
);

INVx4_ASAP7_75t_L g4704 ( 
.A(n_4105),
.Y(n_4704)
);

OAI21xp33_ASAP7_75t_L g4705 ( 
.A1(n_4398),
.A2(n_246),
.B(n_247),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4055),
.B(n_247),
.Y(n_4706)
);

OAI22xp5_ASAP7_75t_L g4707 ( 
.A1(n_3980),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_4707)
);

NAND2x1p5_ASAP7_75t_L g4708 ( 
.A(n_4105),
.B(n_248),
.Y(n_4708)
);

O2A1O1Ixp5_ASAP7_75t_L g4709 ( 
.A1(n_4413),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_4709)
);

NOR2xp33_ASAP7_75t_L g4710 ( 
.A(n_4459),
.B(n_250),
.Y(n_4710)
);

AOI21xp5_ASAP7_75t_L g4711 ( 
.A1(n_4469),
.A2(n_251),
.B(n_252),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_4102),
.B(n_251),
.Y(n_4712)
);

BUFx12f_ASAP7_75t_L g4713 ( 
.A(n_4114),
.Y(n_4713)
);

NOR2xp33_ASAP7_75t_L g4714 ( 
.A(n_4156),
.B(n_252),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4125),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4143),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_SL g4717 ( 
.A(n_4199),
.B(n_252),
.Y(n_4717)
);

NAND3xp33_ASAP7_75t_SL g4718 ( 
.A(n_4224),
.B(n_4226),
.C(n_4319),
.Y(n_4718)
);

OAI22xp5_ASAP7_75t_L g4719 ( 
.A1(n_4047),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_4719)
);

INVx3_ASAP7_75t_SL g4720 ( 
.A(n_4136),
.Y(n_4720)
);

NOR2xp33_ASAP7_75t_L g4721 ( 
.A(n_4427),
.B(n_254),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4132),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_SL g4723 ( 
.A(n_4192),
.B(n_4191),
.Y(n_4723)
);

AOI21xp5_ASAP7_75t_L g4724 ( 
.A1(n_4365),
.A2(n_254),
.B(n_255),
.Y(n_4724)
);

NOR3xp33_ASAP7_75t_SL g4725 ( 
.A(n_4188),
.B(n_256),
.C(n_257),
.Y(n_4725)
);

A2O1A1Ixp33_ASAP7_75t_L g4726 ( 
.A1(n_4296),
.A2(n_259),
.B(n_257),
.C(n_258),
.Y(n_4726)
);

OAI22xp5_ASAP7_75t_SL g4727 ( 
.A1(n_4236),
.A2(n_260),
.B1(n_257),
.B2(n_259),
.Y(n_4727)
);

AOI22xp33_ASAP7_75t_L g4728 ( 
.A1(n_4491),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_SL g4729 ( 
.A(n_4149),
.B(n_260),
.Y(n_4729)
);

AOI22xp5_ASAP7_75t_L g4730 ( 
.A1(n_4351),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_4730)
);

OAI22xp5_ASAP7_75t_L g4731 ( 
.A1(n_4312),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_4731)
);

AOI21xp5_ASAP7_75t_L g4732 ( 
.A1(n_4128),
.A2(n_263),
.B(n_264),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_4135),
.B(n_265),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_SL g4734 ( 
.A(n_4152),
.B(n_266),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4139),
.B(n_267),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4144),
.B(n_267),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4146),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4150),
.B(n_268),
.Y(n_4738)
);

O2A1O1Ixp33_ASAP7_75t_L g4739 ( 
.A1(n_4502),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4165),
.B(n_270),
.Y(n_4740)
);

AOI22xp33_ASAP7_75t_SL g4741 ( 
.A1(n_4326),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_4741)
);

BUFx3_ASAP7_75t_L g4742 ( 
.A(n_4041),
.Y(n_4742)
);

NOR2xp33_ASAP7_75t_L g4743 ( 
.A(n_3999),
.B(n_271),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4285),
.B(n_271),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4286),
.B(n_272),
.Y(n_4745)
);

BUFx3_ASAP7_75t_L g4746 ( 
.A(n_4048),
.Y(n_4746)
);

NAND3xp33_ASAP7_75t_L g4747 ( 
.A(n_4475),
.B(n_4478),
.C(n_4477),
.Y(n_4747)
);

NOR2xp67_ASAP7_75t_L g4748 ( 
.A(n_4105),
.B(n_4164),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4186),
.Y(n_4749)
);

BUFx6f_ASAP7_75t_L g4750 ( 
.A(n_4018),
.Y(n_4750)
);

AOI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_4278),
.A2(n_272),
.B(n_273),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4294),
.B(n_273),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_SL g4753 ( 
.A(n_4164),
.B(n_4300),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_SL g4754 ( 
.A(n_4164),
.B(n_274),
.Y(n_4754)
);

NAND2x1p5_ASAP7_75t_L g4755 ( 
.A(n_4101),
.B(n_274),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_SL g4756 ( 
.A(n_4381),
.B(n_274),
.Y(n_4756)
);

NAND2xp33_ASAP7_75t_SL g4757 ( 
.A(n_4218),
.B(n_275),
.Y(n_4757)
);

AO21x1_ASAP7_75t_L g4758 ( 
.A1(n_4126),
.A2(n_276),
.B(n_277),
.Y(n_4758)
);

O2A1O1Ixp33_ASAP7_75t_L g4759 ( 
.A1(n_4104),
.A2(n_278),
.B(n_276),
.C(n_277),
.Y(n_4759)
);

AOI21xp5_ASAP7_75t_L g4760 ( 
.A1(n_4471),
.A2(n_276),
.B(n_278),
.Y(n_4760)
);

AOI21xp5_ASAP7_75t_L g4761 ( 
.A1(n_3984),
.A2(n_278),
.B(n_279),
.Y(n_4761)
);

BUFx3_ASAP7_75t_L g4762 ( 
.A(n_4183),
.Y(n_4762)
);

AOI21xp5_ASAP7_75t_L g4763 ( 
.A1(n_4239),
.A2(n_279),
.B(n_280),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_SL g4764 ( 
.A(n_4381),
.B(n_279),
.Y(n_4764)
);

BUFx2_ASAP7_75t_L g4765 ( 
.A(n_4097),
.Y(n_4765)
);

OAI22xp5_ASAP7_75t_L g4766 ( 
.A1(n_4236),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_4766)
);

AOI22xp33_ASAP7_75t_L g4767 ( 
.A1(n_4465),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_4767)
);

AOI21xp5_ASAP7_75t_L g4768 ( 
.A1(n_4245),
.A2(n_4346),
.B(n_4212),
.Y(n_4768)
);

INVx4_ASAP7_75t_L g4769 ( 
.A(n_4097),
.Y(n_4769)
);

OR2x6_ASAP7_75t_L g4770 ( 
.A(n_4326),
.B(n_283),
.Y(n_4770)
);

OAI21xp33_ASAP7_75t_L g4771 ( 
.A1(n_4160),
.A2(n_283),
.B(n_284),
.Y(n_4771)
);

BUFx6f_ASAP7_75t_L g4772 ( 
.A(n_4018),
.Y(n_4772)
);

AO22x1_ASAP7_75t_L g4773 ( 
.A1(n_4227),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_4773)
);

INVx2_ASAP7_75t_L g4774 ( 
.A(n_4153),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4194),
.Y(n_4775)
);

AND2x2_ASAP7_75t_L g4776 ( 
.A(n_3977),
.B(n_284),
.Y(n_4776)
);

NAND2xp5_ASAP7_75t_SL g4777 ( 
.A(n_4381),
.B(n_285),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4295),
.B(n_286),
.Y(n_4778)
);

AO21x1_ASAP7_75t_L g4779 ( 
.A1(n_3957),
.A2(n_286),
.B(n_287),
.Y(n_4779)
);

O2A1O1Ixp33_ASAP7_75t_L g4780 ( 
.A1(n_4109),
.A2(n_289),
.B(n_286),
.C(n_288),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4155),
.Y(n_4781)
);

BUFx2_ASAP7_75t_L g4782 ( 
.A(n_4112),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_4297),
.B(n_288),
.Y(n_4783)
);

NAND2xp33_ASAP7_75t_L g4784 ( 
.A(n_4323),
.B(n_289),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_SL g4785 ( 
.A(n_4389),
.B(n_290),
.Y(n_4785)
);

NOR2xp33_ASAP7_75t_L g4786 ( 
.A(n_4166),
.B(n_290),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_SL g4787 ( 
.A(n_4389),
.B(n_290),
.Y(n_4787)
);

O2A1O1Ixp33_ASAP7_75t_L g4788 ( 
.A1(n_4447),
.A2(n_293),
.B(n_291),
.C(n_292),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4301),
.B(n_4304),
.Y(n_4789)
);

INVx3_ASAP7_75t_L g4790 ( 
.A(n_4046),
.Y(n_4790)
);

NOR2xp33_ASAP7_75t_L g4791 ( 
.A(n_4094),
.B(n_3986),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4308),
.B(n_291),
.Y(n_4792)
);

INVx1_ASAP7_75t_SL g4793 ( 
.A(n_4120),
.Y(n_4793)
);

INVx2_ASAP7_75t_L g4794 ( 
.A(n_4162),
.Y(n_4794)
);

OA22x2_ASAP7_75t_L g4795 ( 
.A1(n_4303),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_4795)
);

INVx3_ASAP7_75t_L g4796 ( 
.A(n_4046),
.Y(n_4796)
);

AOI21xp5_ASAP7_75t_L g4797 ( 
.A1(n_4106),
.A2(n_293),
.B(n_294),
.Y(n_4797)
);

OAI22xp5_ASAP7_75t_L g4798 ( 
.A1(n_4501),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4321),
.B(n_295),
.Y(n_4799)
);

BUFx3_ASAP7_75t_L g4800 ( 
.A(n_4123),
.Y(n_4800)
);

BUFx6f_ASAP7_75t_L g4801 ( 
.A(n_4025),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4327),
.B(n_296),
.Y(n_4802)
);

AOI21xp5_ASAP7_75t_L g4803 ( 
.A1(n_4106),
.A2(n_296),
.B(n_297),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_SL g4804 ( 
.A(n_4333),
.B(n_297),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4344),
.B(n_297),
.Y(n_4805)
);

OR2x2_ASAP7_75t_L g4806 ( 
.A(n_3957),
.B(n_298),
.Y(n_4806)
);

AND2x4_ASAP7_75t_L g4807 ( 
.A(n_4317),
.B(n_298),
.Y(n_4807)
);

AOI221xp5_ASAP7_75t_L g4808 ( 
.A1(n_4403),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.C(n_302),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4206),
.Y(n_4809)
);

OAI21xp33_ASAP7_75t_L g4810 ( 
.A1(n_4457),
.A2(n_299),
.B(n_300),
.Y(n_4810)
);

BUFx2_ASAP7_75t_L g4811 ( 
.A(n_4145),
.Y(n_4811)
);

AOI21xp5_ASAP7_75t_L g4812 ( 
.A1(n_4243),
.A2(n_300),
.B(n_301),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_SL g4813 ( 
.A(n_4333),
.B(n_301),
.Y(n_4813)
);

OAI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4501),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_4814)
);

INVx1_ASAP7_75t_SL g4815 ( 
.A(n_4161),
.Y(n_4815)
);

AOI21xp5_ASAP7_75t_L g4816 ( 
.A1(n_4243),
.A2(n_302),
.B(n_303),
.Y(n_4816)
);

BUFx2_ASAP7_75t_L g4817 ( 
.A(n_4410),
.Y(n_4817)
);

INVx2_ASAP7_75t_L g4818 ( 
.A(n_4170),
.Y(n_4818)
);

INVx2_ASAP7_75t_L g4819 ( 
.A(n_4177),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4208),
.Y(n_4820)
);

NOR2xp33_ASAP7_75t_L g4821 ( 
.A(n_4484),
.B(n_304),
.Y(n_4821)
);

NAND2x1p5_ASAP7_75t_L g4822 ( 
.A(n_4021),
.B(n_305),
.Y(n_4822)
);

OAI21x1_ASAP7_75t_L g4823 ( 
.A1(n_4324),
.A2(n_874),
.B(n_864),
.Y(n_4823)
);

AOI21xp5_ASAP7_75t_L g4824 ( 
.A1(n_4265),
.A2(n_4269),
.B(n_4496),
.Y(n_4824)
);

NOR2xp33_ASAP7_75t_L g4825 ( 
.A(n_4211),
.B(n_305),
.Y(n_4825)
);

INVx1_ASAP7_75t_SL g4826 ( 
.A(n_4207),
.Y(n_4826)
);

INVx5_ASAP7_75t_L g4827 ( 
.A(n_4021),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_SL g4828 ( 
.A(n_4348),
.B(n_305),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_L g4829 ( 
.A(n_4352),
.B(n_306),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4201),
.B(n_307),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_SL g4831 ( 
.A(n_4348),
.B(n_307),
.Y(n_4831)
);

NOR2xp33_ASAP7_75t_L g4832 ( 
.A(n_4240),
.B(n_307),
.Y(n_4832)
);

O2A1O1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4458),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4362),
.B(n_308),
.Y(n_4834)
);

AOI21xp5_ASAP7_75t_L g4835 ( 
.A1(n_4265),
.A2(n_308),
.B(n_309),
.Y(n_4835)
);

BUFx6f_ASAP7_75t_L g4836 ( 
.A(n_4025),
.Y(n_4836)
);

O2A1O1Ixp33_ASAP7_75t_L g4837 ( 
.A1(n_4467),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4213),
.Y(n_4838)
);

A2O1A1Ixp33_ASAP7_75t_SL g4839 ( 
.A1(n_4189),
.A2(n_4187),
.B(n_4328),
.C(n_4062),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_SL g4840 ( 
.A(n_4499),
.B(n_310),
.Y(n_4840)
);

INVxp67_ASAP7_75t_L g4841 ( 
.A(n_4337),
.Y(n_4841)
);

INVx2_ASAP7_75t_L g4842 ( 
.A(n_4179),
.Y(n_4842)
);

AOI21xp5_ASAP7_75t_L g4843 ( 
.A1(n_4269),
.A2(n_311),
.B(n_312),
.Y(n_4843)
);

NAND2xp5_ASAP7_75t_L g4844 ( 
.A(n_4366),
.B(n_311),
.Y(n_4844)
);

A2O1A1Ixp33_ASAP7_75t_L g4845 ( 
.A1(n_4086),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_4845)
);

INVx4_ASAP7_75t_L g4846 ( 
.A(n_4062),
.Y(n_4846)
);

NOR2xp33_ASAP7_75t_L g4847 ( 
.A(n_3961),
.B(n_312),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4054),
.B(n_313),
.Y(n_4848)
);

OR2x6_ASAP7_75t_SL g4849 ( 
.A(n_4079),
.B(n_314),
.Y(n_4849)
);

AOI21xp5_ASAP7_75t_L g4850 ( 
.A1(n_4493),
.A2(n_315),
.B(n_316),
.Y(n_4850)
);

AND2x4_ASAP7_75t_L g4851 ( 
.A(n_4317),
.B(n_315),
.Y(n_4851)
);

NOR2xp33_ASAP7_75t_L g4852 ( 
.A(n_4095),
.B(n_315),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4385),
.B(n_317),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_SL g4854 ( 
.A(n_4499),
.B(n_317),
.Y(n_4854)
);

INVx2_ASAP7_75t_L g4855 ( 
.A(n_4190),
.Y(n_4855)
);

INVx3_ASAP7_75t_L g4856 ( 
.A(n_4168),
.Y(n_4856)
);

AOI22xp5_ASAP7_75t_L g4857 ( 
.A1(n_4441),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_4857)
);

AOI21xp5_ASAP7_75t_L g4858 ( 
.A1(n_4493),
.A2(n_318),
.B(n_319),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4495),
.A2(n_318),
.B(n_320),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_SL g4860 ( 
.A(n_4499),
.B(n_320),
.Y(n_4860)
);

A2O1A1Ixp33_ASAP7_75t_L g4861 ( 
.A1(n_4354),
.A2(n_323),
.B(n_321),
.C(n_322),
.Y(n_4861)
);

INVx2_ASAP7_75t_L g4862 ( 
.A(n_4195),
.Y(n_4862)
);

NOR2xp33_ASAP7_75t_L g4863 ( 
.A(n_4215),
.B(n_321),
.Y(n_4863)
);

NAND2xp5_ASAP7_75t_L g4864 ( 
.A(n_4387),
.B(n_4388),
.Y(n_4864)
);

AOI21xp5_ASAP7_75t_L g4865 ( 
.A1(n_4495),
.A2(n_321),
.B(n_322),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4169),
.B(n_322),
.Y(n_4866)
);

A2O1A1Ixp33_ASAP7_75t_L g4867 ( 
.A1(n_4310),
.A2(n_325),
.B(n_323),
.C(n_324),
.Y(n_4867)
);

OAI22xp5_ASAP7_75t_L g4868 ( 
.A1(n_4148),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_4868)
);

NOR2xp33_ASAP7_75t_L g4869 ( 
.A(n_4122),
.B(n_4470),
.Y(n_4869)
);

OAI21xp5_ASAP7_75t_L g4870 ( 
.A1(n_4488),
.A2(n_325),
.B(n_326),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_SL g4871 ( 
.A(n_4322),
.B(n_326),
.Y(n_4871)
);

NOR2xp33_ASAP7_75t_L g4872 ( 
.A(n_4040),
.B(n_327),
.Y(n_4872)
);

CKINVDCx5p33_ASAP7_75t_R g4873 ( 
.A(n_4210),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4171),
.B(n_327),
.Y(n_4874)
);

OAI21xp5_ASAP7_75t_L g4875 ( 
.A1(n_4350),
.A2(n_327),
.B(n_328),
.Y(n_4875)
);

A2O1A1Ixp33_ASAP7_75t_L g4876 ( 
.A1(n_4260),
.A2(n_331),
.B(n_328),
.C(n_329),
.Y(n_4876)
);

INVxp67_ASAP7_75t_L g4877 ( 
.A(n_4019),
.Y(n_4877)
);

O2A1O1Ixp33_ASAP7_75t_L g4878 ( 
.A1(n_4487),
.A2(n_332),
.B(n_329),
.C(n_331),
.Y(n_4878)
);

NOR2xp33_ASAP7_75t_L g4879 ( 
.A(n_4463),
.B(n_329),
.Y(n_4879)
);

NOR2xp33_ASAP7_75t_R g4880 ( 
.A(n_4057),
.B(n_331),
.Y(n_4880)
);

OR2x2_ASAP7_75t_L g4881 ( 
.A(n_4113),
.B(n_332),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4196),
.Y(n_4882)
);

INVx4_ASAP7_75t_L g4883 ( 
.A(n_4202),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4204),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4180),
.B(n_4231),
.Y(n_4885)
);

CKINVDCx5p33_ASAP7_75t_R g4886 ( 
.A(n_4061),
.Y(n_4886)
);

AOI21xp5_ASAP7_75t_L g4887 ( 
.A1(n_4510),
.A2(n_332),
.B(n_333),
.Y(n_4887)
);

OAI22xp5_ASAP7_75t_L g4888 ( 
.A1(n_4512),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4209),
.Y(n_4889)
);

BUFx6f_ASAP7_75t_SL g4890 ( 
.A(n_4151),
.Y(n_4890)
);

AOI21xp5_ASAP7_75t_L g4891 ( 
.A1(n_4510),
.A2(n_334),
.B(n_335),
.Y(n_4891)
);

BUFx3_ASAP7_75t_L g4892 ( 
.A(n_4159),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4087),
.A2(n_334),
.B(n_335),
.Y(n_4893)
);

NOR2xp33_ASAP7_75t_L g4894 ( 
.A(n_4049),
.B(n_336),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4361),
.B(n_336),
.Y(n_4895)
);

A2O1A1Ixp33_ASAP7_75t_L g4896 ( 
.A1(n_4307),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4216),
.Y(n_4897)
);

NAND2xp5_ASAP7_75t_L g4898 ( 
.A(n_4244),
.B(n_338),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_SL g4899 ( 
.A(n_3953),
.B(n_338),
.Y(n_4899)
);

NAND2xp33_ASAP7_75t_SL g4900 ( 
.A(n_4485),
.B(n_339),
.Y(n_4900)
);

INVx3_ASAP7_75t_L g4901 ( 
.A(n_4168),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4386),
.B(n_339),
.Y(n_4902)
);

CKINVDCx16_ASAP7_75t_R g4903 ( 
.A(n_4003),
.Y(n_4903)
);

INVx11_ASAP7_75t_L g4904 ( 
.A(n_4158),
.Y(n_4904)
);

AOI22xp33_ASAP7_75t_L g4905 ( 
.A1(n_4465),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_SL g4906 ( 
.A(n_3953),
.B(n_340),
.Y(n_4906)
);

AOI21xp5_ASAP7_75t_L g4907 ( 
.A1(n_3951),
.A2(n_340),
.B(n_341),
.Y(n_4907)
);

O2A1O1Ixp33_ASAP7_75t_L g4908 ( 
.A1(n_4110),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_4908)
);

OAI21x1_ASAP7_75t_L g4909 ( 
.A1(n_4324),
.A2(n_869),
.B(n_860),
.Y(n_4909)
);

AOI21x1_ASAP7_75t_L g4910 ( 
.A1(n_4292),
.A2(n_342),
.B(n_343),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_SL g4911 ( 
.A(n_3959),
.B(n_343),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4248),
.B(n_344),
.Y(n_4912)
);

BUFx2_ASAP7_75t_L g4913 ( 
.A(n_4330),
.Y(n_4913)
);

NOR2xp33_ASAP7_75t_L g4914 ( 
.A(n_4453),
.B(n_344),
.Y(n_4914)
);

O2A1O1Ixp5_ASAP7_75t_L g4915 ( 
.A1(n_4370),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_SL g4916 ( 
.A(n_3959),
.B(n_345),
.Y(n_4916)
);

O2A1O1Ixp33_ASAP7_75t_L g4917 ( 
.A1(n_4374),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_4917)
);

NAND3xp33_ASAP7_75t_L g4918 ( 
.A(n_4416),
.B(n_347),
.C(n_348),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_SL g4919 ( 
.A(n_3970),
.B(n_348),
.Y(n_4919)
);

AOI21xp5_ASAP7_75t_L g4920 ( 
.A1(n_3958),
.A2(n_350),
.B(n_351),
.Y(n_4920)
);

OAI22xp5_ASAP7_75t_L g4921 ( 
.A1(n_4490),
.A2(n_4089),
.B1(n_4111),
.B2(n_4449),
.Y(n_4921)
);

OAI22xp5_ASAP7_75t_L g4922 ( 
.A1(n_4449),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_4922)
);

NOR2xp33_ASAP7_75t_L g4923 ( 
.A(n_4461),
.B(n_352),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4249),
.Y(n_4924)
);

AND2x2_ASAP7_75t_L g4925 ( 
.A(n_4390),
.B(n_352),
.Y(n_4925)
);

AOI21xp5_ASAP7_75t_L g4926 ( 
.A1(n_3969),
.A2(n_353),
.B(n_354),
.Y(n_4926)
);

INVx2_ASAP7_75t_L g4927 ( 
.A(n_4219),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_SL g4928 ( 
.A(n_3970),
.B(n_353),
.Y(n_4928)
);

AOI21xp5_ASAP7_75t_L g4929 ( 
.A1(n_3972),
.A2(n_354),
.B(n_355),
.Y(n_4929)
);

OR2x6_ASAP7_75t_L g4930 ( 
.A(n_4074),
.B(n_354),
.Y(n_4930)
);

BUFx2_ASAP7_75t_L g4931 ( 
.A(n_4341),
.Y(n_4931)
);

OAI22xp5_ASAP7_75t_L g4932 ( 
.A1(n_4072),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_4932)
);

AOI21xp5_ASAP7_75t_L g4933 ( 
.A1(n_3978),
.A2(n_3991),
.B(n_3987),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4253),
.B(n_355),
.Y(n_4934)
);

INVxp67_ASAP7_75t_SL g4935 ( 
.A(n_4025),
.Y(n_4935)
);

NOR2xp33_ASAP7_75t_L g4936 ( 
.A(n_3993),
.B(n_3995),
.Y(n_4936)
);

HB1xp67_ASAP7_75t_L g4937 ( 
.A(n_3997),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4030),
.A2(n_357),
.B(n_358),
.Y(n_4938)
);

AND2x4_ASAP7_75t_L g4939 ( 
.A(n_4298),
.B(n_357),
.Y(n_4939)
);

CKINVDCx5p33_ASAP7_75t_R g4940 ( 
.A(n_4355),
.Y(n_4940)
);

AOI21xp5_ASAP7_75t_L g4941 ( 
.A1(n_4037),
.A2(n_358),
.B(n_359),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_L g4942 ( 
.A(n_4257),
.B(n_359),
.Y(n_4942)
);

INVx5_ASAP7_75t_L g4943 ( 
.A(n_4060),
.Y(n_4943)
);

NAND3xp33_ASAP7_75t_SL g4944 ( 
.A(n_4141),
.B(n_359),
.C(n_360),
.Y(n_4944)
);

INVx5_ASAP7_75t_L g4945 ( 
.A(n_4060),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_SL g4946 ( 
.A(n_4370),
.B(n_360),
.Y(n_4946)
);

AOI21xp5_ASAP7_75t_L g4947 ( 
.A1(n_4038),
.A2(n_4439),
.B(n_4436),
.Y(n_4947)
);

AOI21xp5_ASAP7_75t_L g4948 ( 
.A1(n_4436),
.A2(n_360),
.B(n_361),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4259),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4000),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_3971),
.B(n_361),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4407),
.B(n_361),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4411),
.B(n_362),
.Y(n_4953)
);

NOR2xp33_ASAP7_75t_L g4954 ( 
.A(n_4027),
.B(n_4404),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4412),
.B(n_362),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_SL g4956 ( 
.A(n_4233),
.B(n_362),
.Y(n_4956)
);

INVx2_ASAP7_75t_SL g4957 ( 
.A(n_4043),
.Y(n_4957)
);

OAI22xp5_ASAP7_75t_L g4958 ( 
.A1(n_4503),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_4958)
);

A2O1A1Ixp33_ASAP7_75t_SL g4959 ( 
.A1(n_4504),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4002),
.Y(n_4960)
);

AND2x2_ASAP7_75t_L g4961 ( 
.A(n_4277),
.B(n_363),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4024),
.Y(n_4962)
);

NOR2xp33_ASAP7_75t_R g4963 ( 
.A(n_4233),
.B(n_365),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4466),
.B(n_366),
.Y(n_4964)
);

AND2x2_ASAP7_75t_L g4965 ( 
.A(n_4402),
.B(n_4167),
.Y(n_4965)
);

INVx4_ASAP7_75t_L g4966 ( 
.A(n_4202),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4414),
.B(n_4418),
.Y(n_4967)
);

INVx2_ASAP7_75t_L g4968 ( 
.A(n_4225),
.Y(n_4968)
);

NAND2xp33_ASAP7_75t_R g4969 ( 
.A(n_4279),
.B(n_366),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4228),
.B(n_366),
.Y(n_4970)
);

HB1xp67_ASAP7_75t_L g4971 ( 
.A(n_4229),
.Y(n_4971)
);

A2O1A1Ixp33_ASAP7_75t_L g4972 ( 
.A1(n_4506),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_4972)
);

BUFx2_ASAP7_75t_L g4973 ( 
.A(n_4371),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4237),
.Y(n_4974)
);

AOI21xp5_ASAP7_75t_L g4975 ( 
.A1(n_4439),
.A2(n_367),
.B(n_368),
.Y(n_4975)
);

INVx4_ASAP7_75t_L g4976 ( 
.A(n_4279),
.Y(n_4976)
);

INVxp67_ASAP7_75t_L g4977 ( 
.A(n_4157),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4424),
.B(n_367),
.Y(n_4978)
);

AND2x4_ASAP7_75t_L g4979 ( 
.A(n_4298),
.B(n_369),
.Y(n_4979)
);

BUFx12f_ASAP7_75t_L g4980 ( 
.A(n_4373),
.Y(n_4980)
);

OAI22xp5_ASAP7_75t_L g4981 ( 
.A1(n_4649),
.A2(n_4417),
.B1(n_4384),
.B2(n_4423),
.Y(n_4981)
);

AND2x2_ASAP7_75t_L g4982 ( 
.A(n_4965),
.B(n_4241),
.Y(n_4982)
);

AND2x4_ASAP7_75t_L g4983 ( 
.A(n_4742),
.B(n_4043),
.Y(n_4983)
);

AOI22xp5_ASAP7_75t_L g4984 ( 
.A1(n_4521),
.A2(n_4430),
.B1(n_4513),
.B2(n_4266),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4977),
.B(n_3975),
.Y(n_4985)
);

NAND2xp5_ASAP7_75t_L g4986 ( 
.A(n_4950),
.B(n_4440),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4903),
.B(n_4258),
.Y(n_4987)
);

HAxp5_ASAP7_75t_L g4988 ( 
.A(n_4616),
.B(n_370),
.CON(n_4988),
.SN(n_4988)
);

AOI22xp33_ASAP7_75t_L g4989 ( 
.A1(n_4526),
.A2(n_4450),
.B1(n_4442),
.B2(n_4299),
.Y(n_4989)
);

BUFx4f_ASAP7_75t_L g4990 ( 
.A(n_4546),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4547),
.Y(n_4991)
);

AOI22xp33_ASAP7_75t_L g4992 ( 
.A1(n_4601),
.A2(n_4311),
.B1(n_4313),
.B2(n_4289),
.Y(n_4992)
);

OAI21xp33_ASAP7_75t_L g4993 ( 
.A1(n_4710),
.A2(n_4880),
.B(n_4637),
.Y(n_4993)
);

BUFx2_ASAP7_75t_L g4994 ( 
.A(n_4817),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4960),
.B(n_4314),
.Y(n_4995)
);

OR2x2_ASAP7_75t_L g4996 ( 
.A(n_4699),
.B(n_4011),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4551),
.Y(n_4997)
);

AOI22xp33_ASAP7_75t_L g4998 ( 
.A1(n_4520),
.A2(n_4334),
.B1(n_4342),
.B2(n_4315),
.Y(n_4998)
);

AND2x4_ASAP7_75t_L g4999 ( 
.A(n_4746),
.B(n_4063),
.Y(n_4999)
);

BUFx3_ASAP7_75t_L g5000 ( 
.A(n_4563),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4566),
.Y(n_5001)
);

BUFx6f_ASAP7_75t_L g5002 ( 
.A(n_4595),
.Y(n_5002)
);

INVx2_ASAP7_75t_L g5003 ( 
.A(n_4971),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4937),
.B(n_4262),
.Y(n_5004)
);

OAI22xp5_ASAP7_75t_L g5005 ( 
.A1(n_4849),
.A2(n_4293),
.B1(n_4473),
.B2(n_4472),
.Y(n_5005)
);

INVx2_ASAP7_75t_SL g5006 ( 
.A(n_4603),
.Y(n_5006)
);

INVx6_ASAP7_75t_L g5007 ( 
.A(n_4681),
.Y(n_5007)
);

AOI22xp33_ASAP7_75t_SL g5008 ( 
.A1(n_4963),
.A2(n_4069),
.B1(n_4071),
.B2(n_4063),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4677),
.B(n_4343),
.Y(n_5009)
);

AOI22xp33_ASAP7_75t_L g5010 ( 
.A1(n_4558),
.A2(n_4369),
.B1(n_4372),
.B2(n_4356),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4962),
.B(n_4380),
.Y(n_5011)
);

BUFx3_ASAP7_75t_L g5012 ( 
.A(n_4515),
.Y(n_5012)
);

NOR2xp33_ASAP7_75t_L g5013 ( 
.A(n_4567),
.B(n_4029),
.Y(n_5013)
);

O2A1O1Ixp33_ASAP7_75t_L g5014 ( 
.A1(n_4639),
.A2(n_4428),
.B(n_4446),
.C(n_4479),
.Y(n_5014)
);

INVxp67_ASAP7_75t_L g5015 ( 
.A(n_4552),
.Y(n_5015)
);

BUFx6f_ASAP7_75t_L g5016 ( 
.A(n_4762),
.Y(n_5016)
);

AOI22xp5_ASAP7_75t_L g5017 ( 
.A1(n_4727),
.A2(n_4405),
.B1(n_4276),
.B2(n_4282),
.Y(n_5017)
);

AND2x2_ASAP7_75t_L g5018 ( 
.A(n_4522),
.B(n_4954),
.Y(n_5018)
);

INVx2_ASAP7_75t_L g5019 ( 
.A(n_4550),
.Y(n_5019)
);

INVx3_ASAP7_75t_L g5020 ( 
.A(n_4554),
.Y(n_5020)
);

INVx4_ASAP7_75t_L g5021 ( 
.A(n_4602),
.Y(n_5021)
);

OAI21xp33_ASAP7_75t_SL g5022 ( 
.A1(n_4700),
.A2(n_4082),
.B(n_4415),
.Y(n_5022)
);

BUFx6f_ASAP7_75t_L g5023 ( 
.A(n_4800),
.Y(n_5023)
);

AND2x4_ASAP7_75t_L g5024 ( 
.A(n_4602),
.B(n_4069),
.Y(n_5024)
);

OR2x6_ASAP7_75t_SL g5025 ( 
.A(n_4873),
.B(n_4400),
.Y(n_5025)
);

OAI22xp5_ASAP7_75t_L g5026 ( 
.A1(n_4770),
.A2(n_4320),
.B1(n_4476),
.B2(n_4408),
.Y(n_5026)
);

A2O1A1Ixp33_ASAP7_75t_L g5027 ( 
.A1(n_4757),
.A2(n_4071),
.B(n_4509),
.C(n_4505),
.Y(n_5027)
);

BUFx12f_ASAP7_75t_L g5028 ( 
.A(n_4680),
.Y(n_5028)
);

BUFx6f_ASAP7_75t_L g5029 ( 
.A(n_4642),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4579),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_4580),
.A2(n_4619),
.B(n_4607),
.Y(n_5031)
);

AOI22xp33_ASAP7_75t_SL g5032 ( 
.A1(n_4592),
.A2(n_4378),
.B1(n_4382),
.B2(n_4401),
.Y(n_5032)
);

CKINVDCx20_ASAP7_75t_R g5033 ( 
.A(n_4574),
.Y(n_5033)
);

AND2x4_ASAP7_75t_L g5034 ( 
.A(n_4602),
.B(n_4376),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_L g5035 ( 
.A(n_4653),
.B(n_4138),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_L g5036 ( 
.A(n_4936),
.B(n_4409),
.Y(n_5036)
);

BUFx12f_ASAP7_75t_L g5037 ( 
.A(n_4681),
.Y(n_5037)
);

CKINVDCx5p33_ASAP7_75t_R g5038 ( 
.A(n_4553),
.Y(n_5038)
);

BUFx2_ASAP7_75t_L g5039 ( 
.A(n_4765),
.Y(n_5039)
);

INVx3_ASAP7_75t_L g5040 ( 
.A(n_4608),
.Y(n_5040)
);

INVx4_ASAP7_75t_L g5041 ( 
.A(n_4549),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4599),
.Y(n_5042)
);

BUFx2_ASAP7_75t_L g5043 ( 
.A(n_4846),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4626),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4562),
.B(n_4589),
.Y(n_5045)
);

BUFx3_ASAP7_75t_L g5046 ( 
.A(n_4625),
.Y(n_5046)
);

BUFx6f_ASAP7_75t_L g5047 ( 
.A(n_4631),
.Y(n_5047)
);

NAND2x1p5_ASAP7_75t_L g5048 ( 
.A(n_4586),
.B(n_3979),
.Y(n_5048)
);

CKINVDCx5p33_ASAP7_75t_R g5049 ( 
.A(n_4713),
.Y(n_5049)
);

AOI22xp5_ASAP7_75t_L g5050 ( 
.A1(n_4784),
.A2(n_4284),
.B1(n_4275),
.B2(n_4391),
.Y(n_5050)
);

OR2x6_ASAP7_75t_L g5051 ( 
.A(n_4770),
.B(n_4263),
.Y(n_5051)
);

BUFx2_ASAP7_75t_L g5052 ( 
.A(n_4846),
.Y(n_5052)
);

A2O1A1Ixp33_ASAP7_75t_L g5053 ( 
.A1(n_4900),
.A2(n_3989),
.B(n_4007),
.C(n_3979),
.Y(n_5053)
);

OR2x6_ASAP7_75t_L g5054 ( 
.A(n_4769),
.B(n_4748),
.Y(n_5054)
);

INVx2_ASAP7_75t_L g5055 ( 
.A(n_4557),
.Y(n_5055)
);

NAND3xp33_ASAP7_75t_L g5056 ( 
.A(n_4673),
.B(n_4406),
.C(n_4353),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4633),
.Y(n_5057)
);

AOI22xp5_ASAP7_75t_L g5058 ( 
.A1(n_4969),
.A2(n_4534),
.B1(n_4679),
.B2(n_4667),
.Y(n_5058)
);

CKINVDCx8_ASAP7_75t_R g5059 ( 
.A(n_4628),
.Y(n_5059)
);

INVx4_ASAP7_75t_L g5060 ( 
.A(n_4586),
.Y(n_5060)
);

INVxp67_ASAP7_75t_SL g5061 ( 
.A(n_4638),
.Y(n_5061)
);

INVx2_ASAP7_75t_SL g5062 ( 
.A(n_4543),
.Y(n_5062)
);

BUFx3_ASAP7_75t_L g5063 ( 
.A(n_4782),
.Y(n_5063)
);

BUFx12f_ASAP7_75t_L g5064 ( 
.A(n_4665),
.Y(n_5064)
);

AND2x4_ASAP7_75t_L g5065 ( 
.A(n_4769),
.B(n_3989),
.Y(n_5065)
);

OAI22xp33_ASAP7_75t_L g5066 ( 
.A1(n_4930),
.A2(n_4247),
.B1(n_4425),
.B2(n_4422),
.Y(n_5066)
);

BUFx6f_ASAP7_75t_L g5067 ( 
.A(n_4811),
.Y(n_5067)
);

O2A1O1Ixp33_ASAP7_75t_L g5068 ( 
.A1(n_4644),
.A2(n_4329),
.B(n_4392),
.C(n_4433),
.Y(n_5068)
);

BUFx4f_ASAP7_75t_L g5069 ( 
.A(n_4930),
.Y(n_5069)
);

NAND3xp33_ASAP7_75t_L g5070 ( 
.A(n_4725),
.B(n_4444),
.C(n_4438),
.Y(n_5070)
);

AND2x2_ASAP7_75t_L g5071 ( 
.A(n_4594),
.B(n_4271),
.Y(n_5071)
);

INVx1_ASAP7_75t_L g5072 ( 
.A(n_4655),
.Y(n_5072)
);

INVx3_ASAP7_75t_L g5073 ( 
.A(n_4675),
.Y(n_5073)
);

BUFx2_ASAP7_75t_L g5074 ( 
.A(n_4913),
.Y(n_5074)
);

OAI22xp5_ASAP7_75t_L g5075 ( 
.A1(n_4524),
.A2(n_4448),
.B1(n_4452),
.B2(n_4456),
.Y(n_5075)
);

AND2x4_ASAP7_75t_L g5076 ( 
.A(n_4645),
.B(n_4883),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_4671),
.Y(n_5077)
);

INVxp67_ASAP7_75t_L g5078 ( 
.A(n_4702),
.Y(n_5078)
);

INVx3_ASAP7_75t_L g5079 ( 
.A(n_4675),
.Y(n_5079)
);

BUFx2_ASAP7_75t_L g5080 ( 
.A(n_4931),
.Y(n_5080)
);

OR2x2_ASAP7_75t_L g5081 ( 
.A(n_4612),
.B(n_4256),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4687),
.Y(n_5082)
);

OR2x4_ASAP7_75t_L g5083 ( 
.A(n_4591),
.B(n_4360),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4715),
.Y(n_5084)
);

OAI22xp5_ASAP7_75t_L g5085 ( 
.A1(n_4741),
.A2(n_4287),
.B1(n_4283),
.B2(n_4331),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4722),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4737),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4924),
.Y(n_5088)
);

OR2x6_ASAP7_75t_L g5089 ( 
.A(n_4883),
.B(n_4007),
.Y(n_5089)
);

BUFx2_ASAP7_75t_L g5090 ( 
.A(n_4973),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_4791),
.B(n_4377),
.Y(n_5091)
);

OR2x6_ASAP7_75t_L g5092 ( 
.A(n_4966),
.B(n_4395),
.Y(n_5092)
);

AOI21xp5_ASAP7_75t_L g5093 ( 
.A1(n_4518),
.A2(n_4395),
.B(n_4379),
.Y(n_5093)
);

NAND2x1p5_ASAP7_75t_L g5094 ( 
.A(n_4686),
.B(n_4704),
.Y(n_5094)
);

INVx2_ASAP7_75t_L g5095 ( 
.A(n_4561),
.Y(n_5095)
);

INVx3_ASAP7_75t_L g5096 ( 
.A(n_4686),
.Y(n_5096)
);

BUFx2_ASAP7_75t_L g5097 ( 
.A(n_4570),
.Y(n_5097)
);

AND2x4_ASAP7_75t_L g5098 ( 
.A(n_4966),
.B(n_4379),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4949),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4539),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_4749),
.Y(n_5101)
);

BUFx3_ASAP7_75t_L g5102 ( 
.A(n_4892),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_4775),
.Y(n_5103)
);

HB1xp67_ASAP7_75t_L g5104 ( 
.A(n_4565),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_4809),
.Y(n_5105)
);

OAI22xp5_ASAP7_75t_L g5106 ( 
.A1(n_4530),
.A2(n_4349),
.B1(n_4338),
.B2(n_4309),
.Y(n_5106)
);

INVx4_ASAP7_75t_L g5107 ( 
.A(n_4890),
.Y(n_5107)
);

INVx2_ASAP7_75t_SL g5108 ( 
.A(n_4793),
.Y(n_5108)
);

INVx1_ASAP7_75t_SL g5109 ( 
.A(n_4815),
.Y(n_5109)
);

AOI22xp33_ASAP7_75t_L g5110 ( 
.A1(n_4705),
.A2(n_4697),
.B1(n_4944),
.B2(n_4939),
.Y(n_5110)
);

HB1xp67_ASAP7_75t_L g5111 ( 
.A(n_4841),
.Y(n_5111)
);

AOI22xp5_ASAP7_75t_L g5112 ( 
.A1(n_4541),
.A2(n_4272),
.B1(n_4273),
.B2(n_4375),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_4578),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4820),
.Y(n_5114)
);

INVx3_ASAP7_75t_L g5115 ( 
.A(n_4704),
.Y(n_5115)
);

OR2x6_ASAP7_75t_L g5116 ( 
.A(n_4535),
.B(n_4184),
.Y(n_5116)
);

INVx4_ASAP7_75t_L g5117 ( 
.A(n_4886),
.Y(n_5117)
);

BUFx2_ASAP7_75t_L g5118 ( 
.A(n_4583),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4838),
.Y(n_5119)
);

BUFx3_ASAP7_75t_L g5120 ( 
.A(n_4606),
.Y(n_5120)
);

AOI21xp5_ASAP7_75t_L g5121 ( 
.A1(n_4641),
.A2(n_4332),
.B(n_4396),
.Y(n_5121)
);

INVx5_ASAP7_75t_L g5122 ( 
.A(n_4514),
.Y(n_5122)
);

OAI22xp33_ASAP7_75t_L g5123 ( 
.A1(n_4535),
.A2(n_4455),
.B1(n_4437),
.B2(n_4443),
.Y(n_5123)
);

CKINVDCx5p33_ASAP7_75t_R g5124 ( 
.A(n_4596),
.Y(n_5124)
);

INVx3_ASAP7_75t_L g5125 ( 
.A(n_4827),
.Y(n_5125)
);

AOI22xp33_ASAP7_75t_L g5126 ( 
.A1(n_4697),
.A2(n_4480),
.B1(n_4451),
.B2(n_4383),
.Y(n_5126)
);

OR2x2_ASAP7_75t_L g5127 ( 
.A(n_4556),
.B(n_4251),
.Y(n_5127)
);

AND2x4_ASAP7_75t_L g5128 ( 
.A(n_4661),
.B(n_4332),
.Y(n_5128)
);

NOR2xp33_ASAP7_75t_L g5129 ( 
.A(n_4826),
.B(n_370),
.Y(n_5129)
);

AOI22xp33_ASAP7_75t_L g5130 ( 
.A1(n_4939),
.A2(n_4451),
.B1(n_4383),
.B2(n_4235),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_4897),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_4885),
.Y(n_5132)
);

BUFx6f_ASAP7_75t_L g5133 ( 
.A(n_4660),
.Y(n_5133)
);

CKINVDCx5p33_ASAP7_75t_R g5134 ( 
.A(n_4720),
.Y(n_5134)
);

BUFx12f_ASAP7_75t_L g5135 ( 
.A(n_4940),
.Y(n_5135)
);

OR2x6_ASAP7_75t_L g5136 ( 
.A(n_4980),
.B(n_4383),
.Y(n_5136)
);

OR2x6_ASAP7_75t_L g5137 ( 
.A(n_4514),
.B(n_4451),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4658),
.Y(n_5138)
);

BUFx2_ASAP7_75t_L g5139 ( 
.A(n_4976),
.Y(n_5139)
);

INVx5_ASAP7_75t_L g5140 ( 
.A(n_4827),
.Y(n_5140)
);

INVx2_ASAP7_75t_L g5141 ( 
.A(n_4611),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_4967),
.Y(n_5142)
);

INVx1_ASAP7_75t_SL g5143 ( 
.A(n_4830),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_4789),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4864),
.Y(n_5145)
);

INVx2_ASAP7_75t_SL g5146 ( 
.A(n_4827),
.Y(n_5146)
);

BUFx6f_ASAP7_75t_L g5147 ( 
.A(n_4660),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_4620),
.Y(n_5148)
);

INVx2_ASAP7_75t_L g5149 ( 
.A(n_4666),
.Y(n_5149)
);

NOR2xp33_ASAP7_75t_L g5150 ( 
.A(n_4877),
.B(n_370),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_4669),
.Y(n_5151)
);

INVx4_ASAP7_75t_L g5152 ( 
.A(n_4904),
.Y(n_5152)
);

NOR2xp33_ASAP7_75t_R g5153 ( 
.A(n_4718),
.B(n_371),
.Y(n_5153)
);

INVx2_ASAP7_75t_L g5154 ( 
.A(n_4678),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_4682),
.Y(n_5155)
);

CKINVDCx5p33_ASAP7_75t_R g5156 ( 
.A(n_4590),
.Y(n_5156)
);

CKINVDCx5p33_ASAP7_75t_R g5157 ( 
.A(n_4872),
.Y(n_5157)
);

CKINVDCx11_ASAP7_75t_R g5158 ( 
.A(n_4674),
.Y(n_5158)
);

OAI22xp5_ASAP7_75t_L g5159 ( 
.A1(n_4568),
.A2(n_4108),
.B1(n_4116),
.B2(n_4060),
.Y(n_5159)
);

BUFx8_ASAP7_75t_L g5160 ( 
.A(n_4674),
.Y(n_5160)
);

AND2x4_ASAP7_75t_L g5161 ( 
.A(n_4661),
.B(n_4976),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_SL g5162 ( 
.A(n_4528),
.B(n_4108),
.Y(n_5162)
);

BUFx6f_ASAP7_75t_L g5163 ( 
.A(n_4660),
.Y(n_5163)
);

INVx4_ASAP7_75t_L g5164 ( 
.A(n_4708),
.Y(n_5164)
);

BUFx6f_ASAP7_75t_L g5165 ( 
.A(n_4750),
.Y(n_5165)
);

INVx1_ASAP7_75t_L g5166 ( 
.A(n_4690),
.Y(n_5166)
);

AOI21x1_ASAP7_75t_L g5167 ( 
.A1(n_4634),
.A2(n_4609),
.B(n_4753),
.Y(n_5167)
);

AND2x4_ASAP7_75t_L g5168 ( 
.A(n_4957),
.B(n_4807),
.Y(n_5168)
);

BUFx5_ASAP7_75t_L g5169 ( 
.A(n_4807),
.Y(n_5169)
);

BUFx6f_ASAP7_75t_L g5170 ( 
.A(n_4750),
.Y(n_5170)
);

NAND2x1p5_ASAP7_75t_L g5171 ( 
.A(n_4531),
.B(n_4108),
.Y(n_5171)
);

NOR2xp33_ASAP7_75t_L g5172 ( 
.A(n_4523),
.B(n_371),
.Y(n_5172)
);

BUFx3_ASAP7_75t_L g5173 ( 
.A(n_4856),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_4716),
.Y(n_5174)
);

BUFx4f_ASAP7_75t_SL g5175 ( 
.A(n_4851),
.Y(n_5175)
);

BUFx2_ASAP7_75t_L g5176 ( 
.A(n_4621),
.Y(n_5176)
);

INVx3_ASAP7_75t_L g5177 ( 
.A(n_4755),
.Y(n_5177)
);

BUFx2_ASAP7_75t_L g5178 ( 
.A(n_4935),
.Y(n_5178)
);

INVxp67_ASAP7_75t_L g5179 ( 
.A(n_4879),
.Y(n_5179)
);

AND2x4_ASAP7_75t_L g5180 ( 
.A(n_4851),
.B(n_4116),
.Y(n_5180)
);

AOI22xp5_ASAP7_75t_L g5181 ( 
.A1(n_4538),
.A2(n_4235),
.B1(n_4158),
.B2(n_4134),
.Y(n_5181)
);

INVx2_ASAP7_75t_L g5182 ( 
.A(n_4774),
.Y(n_5182)
);

AND2x2_ASAP7_75t_L g5183 ( 
.A(n_4776),
.B(n_4116),
.Y(n_5183)
);

AOI22xp33_ASAP7_75t_L g5184 ( 
.A1(n_4979),
.A2(n_4723),
.B1(n_4771),
.B2(n_4731),
.Y(n_5184)
);

INVx2_ASAP7_75t_L g5185 ( 
.A(n_4781),
.Y(n_5185)
);

OAI22xp5_ASAP7_75t_L g5186 ( 
.A1(n_4647),
.A2(n_4173),
.B1(n_4178),
.B2(n_4134),
.Y(n_5186)
);

INVx4_ASAP7_75t_L g5187 ( 
.A(n_4943),
.Y(n_5187)
);

AOI22xp33_ASAP7_75t_L g5188 ( 
.A1(n_4979),
.A2(n_4158),
.B1(n_4235),
.B2(n_4173),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_SL g5189 ( 
.A(n_4577),
.B(n_4134),
.Y(n_5189)
);

NOR2xp33_ASAP7_75t_L g5190 ( 
.A(n_4533),
.B(n_371),
.Y(n_5190)
);

AND2x2_ASAP7_75t_L g5191 ( 
.A(n_4869),
.B(n_4794),
.Y(n_5191)
);

INVx1_ASAP7_75t_SL g5192 ( 
.A(n_4605),
.Y(n_5192)
);

HB1xp67_ASAP7_75t_L g5193 ( 
.A(n_4921),
.Y(n_5193)
);

INVx4_ASAP7_75t_L g5194 ( 
.A(n_4943),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_4818),
.Y(n_5195)
);

OAI22xp33_ASAP7_75t_L g5196 ( 
.A1(n_4795),
.A2(n_4339),
.B1(n_4340),
.B2(n_4302),
.Y(n_5196)
);

AND2x4_ASAP7_75t_L g5197 ( 
.A(n_4856),
.B(n_4173),
.Y(n_5197)
);

AND2x2_ASAP7_75t_L g5198 ( 
.A(n_4819),
.B(n_4178),
.Y(n_5198)
);

AND2x2_ASAP7_75t_L g5199 ( 
.A(n_4842),
.B(n_4178),
.Y(n_5199)
);

AND2x2_ASAP7_75t_L g5200 ( 
.A(n_4855),
.B(n_4197),
.Y(n_5200)
);

INVx2_ASAP7_75t_L g5201 ( 
.A(n_4862),
.Y(n_5201)
);

CKINVDCx8_ASAP7_75t_R g5202 ( 
.A(n_4786),
.Y(n_5202)
);

AND2x2_ASAP7_75t_L g5203 ( 
.A(n_4882),
.B(n_4197),
.Y(n_5203)
);

AND2x4_ASAP7_75t_L g5204 ( 
.A(n_4901),
.B(n_4790),
.Y(n_5204)
);

NOR2xp33_ASAP7_75t_L g5205 ( 
.A(n_4517),
.B(n_372),
.Y(n_5205)
);

AND2x2_ASAP7_75t_SL g5206 ( 
.A(n_4721),
.B(n_4340),
.Y(n_5206)
);

AOI22xp5_ASAP7_75t_L g5207 ( 
.A1(n_4525),
.A2(n_4235),
.B1(n_4158),
.B2(n_4234),
.Y(n_5207)
);

NOR2xp67_ASAP7_75t_L g5208 ( 
.A(n_4821),
.B(n_372),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_4884),
.B(n_4197),
.Y(n_5209)
);

INVx5_ASAP7_75t_L g5210 ( 
.A(n_4943),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_4889),
.Y(n_5211)
);

NAND2xp5_ASAP7_75t_L g5212 ( 
.A(n_4927),
.B(n_372),
.Y(n_5212)
);

INVx1_ASAP7_75t_SL g5213 ( 
.A(n_4643),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_4968),
.Y(n_5214)
);

BUFx2_ASAP7_75t_L g5215 ( 
.A(n_4790),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_4974),
.Y(n_5216)
);

BUFx10_ASAP7_75t_L g5217 ( 
.A(n_4863),
.Y(n_5217)
);

AOI22xp33_ASAP7_75t_L g5218 ( 
.A1(n_4657),
.A2(n_4280),
.B1(n_4302),
.B2(n_4234),
.Y(n_5218)
);

INVx2_ASAP7_75t_L g5219 ( 
.A(n_4970),
.Y(n_5219)
);

INVx2_ASAP7_75t_L g5220 ( 
.A(n_4848),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_4961),
.B(n_373),
.Y(n_5221)
);

NOR2x1_ASAP7_75t_SL g5222 ( 
.A(n_4635),
.B(n_4234),
.Y(n_5222)
);

BUFx6f_ASAP7_75t_L g5223 ( 
.A(n_4750),
.Y(n_5223)
);

OAI211xp5_ASAP7_75t_SL g5224 ( 
.A1(n_4600),
.A2(n_375),
.B(n_373),
.C(n_374),
.Y(n_5224)
);

INVx3_ASAP7_75t_L g5225 ( 
.A(n_4822),
.Y(n_5225)
);

AND2x2_ASAP7_75t_L g5226 ( 
.A(n_4895),
.B(n_4902),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_4806),
.Y(n_5227)
);

BUFx4f_ASAP7_75t_L g5228 ( 
.A(n_4964),
.Y(n_5228)
);

BUFx3_ASAP7_75t_L g5229 ( 
.A(n_4901),
.Y(n_5229)
);

AND2x4_ASAP7_75t_L g5230 ( 
.A(n_4796),
.B(n_4280),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_4933),
.Y(n_5231)
);

INVx2_ASAP7_75t_SL g5232 ( 
.A(n_4945),
.Y(n_5232)
);

NAND2x1p5_ASAP7_75t_L g5233 ( 
.A(n_4564),
.B(n_4280),
.Y(n_5233)
);

BUFx2_ASAP7_75t_L g5234 ( 
.A(n_4796),
.Y(n_5234)
);

AOI22xp5_ASAP7_75t_L g5235 ( 
.A1(n_4852),
.A2(n_4339),
.B1(n_4340),
.B2(n_4302),
.Y(n_5235)
);

AOI22xp33_ASAP7_75t_L g5236 ( 
.A1(n_4747),
.A2(n_4363),
.B1(n_4364),
.B2(n_4339),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_4925),
.Y(n_5237)
);

AOI221xp5_ASAP7_75t_L g5238 ( 
.A1(n_4650),
.A2(n_4364),
.B1(n_4363),
.B2(n_375),
.C(n_373),
.Y(n_5238)
);

BUFx8_ASAP7_75t_SL g5239 ( 
.A(n_4575),
.Y(n_5239)
);

AND2x4_ASAP7_75t_L g5240 ( 
.A(n_4945),
.B(n_4363),
.Y(n_5240)
);

INVx1_ASAP7_75t_L g5241 ( 
.A(n_4663),
.Y(n_5241)
);

BUFx12f_ASAP7_75t_L g5242 ( 
.A(n_4945),
.Y(n_5242)
);

BUFx6f_ASAP7_75t_L g5243 ( 
.A(n_4772),
.Y(n_5243)
);

INVxp67_ASAP7_75t_L g5244 ( 
.A(n_4825),
.Y(n_5244)
);

BUFx6f_ASAP7_75t_L g5245 ( 
.A(n_4772),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_4951),
.B(n_374),
.Y(n_5246)
);

INVx4_ASAP7_75t_L g5247 ( 
.A(n_4772),
.Y(n_5247)
);

BUFx6f_ASAP7_75t_L g5248 ( 
.A(n_4801),
.Y(n_5248)
);

OAI22xp5_ASAP7_75t_L g5249 ( 
.A1(n_4726),
.A2(n_4364),
.B1(n_377),
.B2(n_374),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_4668),
.Y(n_5250)
);

BUFx10_ASAP7_75t_L g5251 ( 
.A(n_4610),
.Y(n_5251)
);

AOI22xp5_ASAP7_75t_L g5252 ( 
.A1(n_4798),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_4881),
.B(n_376),
.Y(n_5253)
);

AOI22xp33_ASAP7_75t_L g5254 ( 
.A1(n_4814),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_5254)
);

INVx2_ASAP7_75t_SL g5255 ( 
.A(n_4576),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_4555),
.B(n_378),
.Y(n_5256)
);

INVx2_ASAP7_75t_L g5257 ( 
.A(n_4801),
.Y(n_5257)
);

AOI22xp33_ASAP7_75t_L g5258 ( 
.A1(n_4868),
.A2(n_382),
.B1(n_379),
.B2(n_381),
.Y(n_5258)
);

AOI22xp5_ASAP7_75t_L g5259 ( 
.A1(n_4684),
.A2(n_382),
.B1(n_379),
.B2(n_381),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_4542),
.B(n_381),
.Y(n_5260)
);

INVx2_ASAP7_75t_SL g5261 ( 
.A(n_4582),
.Y(n_5261)
);

NOR2xp33_ASAP7_75t_L g5262 ( 
.A(n_4622),
.B(n_382),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_4685),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_4572),
.B(n_383),
.Y(n_5264)
);

BUFx10_ASAP7_75t_L g5265 ( 
.A(n_4698),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_4688),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_4693),
.Y(n_5267)
);

CKINVDCx5p33_ASAP7_75t_R g5268 ( 
.A(n_4832),
.Y(n_5268)
);

NOR2xp33_ASAP7_75t_L g5269 ( 
.A(n_4714),
.B(n_383),
.Y(n_5269)
);

OAI22xp5_ASAP7_75t_L g5270 ( 
.A1(n_4701),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_4703),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_4537),
.B(n_384),
.Y(n_5272)
);

INVx1_ASAP7_75t_L g5273 ( 
.A(n_4706),
.Y(n_5273)
);

INVx2_ASAP7_75t_SL g5274 ( 
.A(n_4584),
.Y(n_5274)
);

CKINVDCx20_ASAP7_75t_R g5275 ( 
.A(n_4652),
.Y(n_5275)
);

A2O1A1Ixp33_ASAP7_75t_L g5276 ( 
.A1(n_4604),
.A2(n_387),
.B(n_385),
.C(n_386),
.Y(n_5276)
);

INVx2_ASAP7_75t_L g5277 ( 
.A(n_4801),
.Y(n_5277)
);

CKINVDCx8_ASAP7_75t_R g5278 ( 
.A(n_4743),
.Y(n_5278)
);

NAND2xp5_ASAP7_75t_L g5279 ( 
.A(n_4529),
.B(n_4847),
.Y(n_5279)
);

BUFx6f_ASAP7_75t_L g5280 ( 
.A(n_4836),
.Y(n_5280)
);

A2O1A1Ixp33_ASAP7_75t_L g5281 ( 
.A1(n_4613),
.A2(n_387),
.B(n_385),
.C(n_386),
.Y(n_5281)
);

BUFx3_ASAP7_75t_L g5282 ( 
.A(n_4836),
.Y(n_5282)
);

CKINVDCx20_ASAP7_75t_R g5283 ( 
.A(n_5033),
.Y(n_5283)
);

AOI22xp33_ASAP7_75t_L g5284 ( 
.A1(n_5010),
.A2(n_4694),
.B1(n_4581),
.B2(n_4758),
.Y(n_5284)
);

A2O1A1Ixp33_ASAP7_75t_L g5285 ( 
.A1(n_5069),
.A2(n_4624),
.B(n_4908),
.C(n_4780),
.Y(n_5285)
);

INVx2_ASAP7_75t_SL g5286 ( 
.A(n_5047),
.Y(n_5286)
);

CKINVDCx5p33_ASAP7_75t_R g5287 ( 
.A(n_5037),
.Y(n_5287)
);

A2O1A1Ixp33_ASAP7_75t_L g5288 ( 
.A1(n_4993),
.A2(n_5008),
.B(n_5022),
.C(n_5058),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_4991),
.Y(n_5289)
);

AND2x2_ASAP7_75t_L g5290 ( 
.A(n_5191),
.B(n_4947),
.Y(n_5290)
);

A2O1A1Ixp33_ASAP7_75t_L g5291 ( 
.A1(n_5205),
.A2(n_4759),
.B(n_4692),
.C(n_4739),
.Y(n_5291)
);

INVx2_ASAP7_75t_L g5292 ( 
.A(n_5003),
.Y(n_5292)
);

OAI221xp5_ASAP7_75t_L g5293 ( 
.A1(n_4989),
.A2(n_4839),
.B1(n_4870),
.B2(n_4659),
.C(n_4857),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_4997),
.Y(n_5294)
);

AOI21xp5_ASAP7_75t_L g5295 ( 
.A1(n_5031),
.A2(n_5162),
.B(n_5066),
.Y(n_5295)
);

INVx5_ASAP7_75t_SL g5296 ( 
.A(n_5047),
.Y(n_5296)
);

AOI21xp5_ASAP7_75t_L g5297 ( 
.A1(n_5189),
.A2(n_4597),
.B(n_4824),
.Y(n_5297)
);

AND2x4_ASAP7_75t_L g5298 ( 
.A(n_5043),
.B(n_4836),
.Y(n_5298)
);

O2A1O1Ixp33_ASAP7_75t_L g5299 ( 
.A1(n_4988),
.A2(n_4614),
.B(n_4745),
.C(n_4744),
.Y(n_5299)
);

INVx1_ASAP7_75t_L g5300 ( 
.A(n_5001),
.Y(n_5300)
);

BUFx3_ASAP7_75t_L g5301 ( 
.A(n_5012),
.Y(n_5301)
);

OR2x2_ASAP7_75t_L g5302 ( 
.A(n_4994),
.B(n_4712),
.Y(n_5302)
);

NAND2xp5_ASAP7_75t_L g5303 ( 
.A(n_5142),
.B(n_4914),
.Y(n_5303)
);

AOI21x1_ASAP7_75t_L g5304 ( 
.A1(n_5167),
.A2(n_4910),
.B(n_4773),
.Y(n_5304)
);

OAI22xp33_ASAP7_75t_L g5305 ( 
.A1(n_5025),
.A2(n_5175),
.B1(n_5116),
.B2(n_5050),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_5144),
.B(n_4923),
.Y(n_5306)
);

AOI21xp5_ASAP7_75t_L g5307 ( 
.A1(n_5052),
.A2(n_5186),
.B(n_5106),
.Y(n_5307)
);

OAI21x1_ASAP7_75t_L g5308 ( 
.A1(n_5094),
.A2(n_5093),
.B(n_5115),
.Y(n_5308)
);

O2A1O1Ixp33_ASAP7_75t_L g5309 ( 
.A1(n_5014),
.A2(n_4778),
.B(n_4783),
.C(n_4752),
.Y(n_5309)
);

A2O1A1Ixp33_ASAP7_75t_L g5310 ( 
.A1(n_5228),
.A2(n_4689),
.B(n_4833),
.C(n_4788),
.Y(n_5310)
);

O2A1O1Ixp33_ASAP7_75t_L g5311 ( 
.A1(n_5068),
.A2(n_4792),
.B(n_4802),
.C(n_4799),
.Y(n_5311)
);

O2A1O1Ixp33_ASAP7_75t_L g5312 ( 
.A1(n_5224),
.A2(n_5281),
.B(n_5276),
.C(n_5256),
.Y(n_5312)
);

NOR2xp33_ASAP7_75t_L g5313 ( 
.A(n_5059),
.B(n_4894),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_5030),
.Y(n_5314)
);

AOI221xp5_ASAP7_75t_L g5315 ( 
.A1(n_5056),
.A2(n_4766),
.B1(n_4588),
.B2(n_4917),
.C(n_4837),
.Y(n_5315)
);

BUFx2_ASAP7_75t_R g5316 ( 
.A(n_5038),
.Y(n_5316)
);

NOR2xp33_ASAP7_75t_L g5317 ( 
.A(n_5041),
.B(n_4805),
.Y(n_5317)
);

AOI21xp5_ASAP7_75t_L g5318 ( 
.A1(n_5121),
.A2(n_4598),
.B(n_4593),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_5042),
.Y(n_5319)
);

INVx2_ASAP7_75t_L g5320 ( 
.A(n_5178),
.Y(n_5320)
);

INVxp67_ASAP7_75t_L g5321 ( 
.A(n_5074),
.Y(n_5321)
);

BUFx12f_ASAP7_75t_L g5322 ( 
.A(n_5028),
.Y(n_5322)
);

AOI22xp5_ASAP7_75t_L g5323 ( 
.A1(n_5184),
.A2(n_4810),
.B1(n_4918),
.B2(n_4754),
.Y(n_5323)
);

AOI21xp5_ASAP7_75t_L g5324 ( 
.A1(n_5116),
.A2(n_4640),
.B(n_4768),
.Y(n_5324)
);

NAND2x1p5_ASAP7_75t_L g5325 ( 
.A(n_4990),
.B(n_4717),
.Y(n_5325)
);

O2A1O1Ixp33_ASAP7_75t_L g5326 ( 
.A1(n_5272),
.A2(n_4834),
.B(n_4844),
.C(n_4829),
.Y(n_5326)
);

AO31x2_ASAP7_75t_L g5327 ( 
.A1(n_5139),
.A2(n_4779),
.A3(n_4617),
.B(n_4691),
.Y(n_5327)
);

AO31x2_ASAP7_75t_L g5328 ( 
.A1(n_5222),
.A2(n_4569),
.A3(n_4763),
.B(n_4896),
.Y(n_5328)
);

NOR2xp67_ASAP7_75t_SL g5329 ( 
.A(n_5140),
.B(n_4656),
.Y(n_5329)
);

BUFx6f_ASAP7_75t_L g5330 ( 
.A(n_5242),
.Y(n_5330)
);

BUFx2_ASAP7_75t_L g5331 ( 
.A(n_5054),
.Y(n_5331)
);

O2A1O1Ixp33_ASAP7_75t_SL g5332 ( 
.A1(n_5062),
.A2(n_4911),
.B(n_4919),
.C(n_4916),
.Y(n_5332)
);

INVxp67_ASAP7_75t_L g5333 ( 
.A(n_5080),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_5044),
.Y(n_5334)
);

AO31x2_ASAP7_75t_L g5335 ( 
.A1(n_5159),
.A2(n_4922),
.A3(n_4683),
.B(n_4876),
.Y(n_5335)
);

BUFx6f_ASAP7_75t_L g5336 ( 
.A(n_5029),
.Y(n_5336)
);

AOI21xp5_ASAP7_75t_L g5337 ( 
.A1(n_5053),
.A2(n_4532),
.B(n_4527),
.Y(n_5337)
);

OR2x2_ASAP7_75t_L g5338 ( 
.A(n_5061),
.B(n_4733),
.Y(n_5338)
);

AOI21xp5_ASAP7_75t_L g5339 ( 
.A1(n_5196),
.A2(n_4540),
.B(n_4536),
.Y(n_5339)
);

A2O1A1Ixp33_ASAP7_75t_L g5340 ( 
.A1(n_5208),
.A2(n_5017),
.B(n_5225),
.C(n_5110),
.Y(n_5340)
);

AOI31xp67_ASAP7_75t_L g5341 ( 
.A1(n_5257),
.A2(n_4676),
.A3(n_4672),
.B(n_4840),
.Y(n_5341)
);

AO31x2_ASAP7_75t_L g5342 ( 
.A1(n_5215),
.A2(n_4874),
.A3(n_4898),
.B(n_4866),
.Y(n_5342)
);

AOI22xp5_ASAP7_75t_L g5343 ( 
.A1(n_4984),
.A2(n_4730),
.B1(n_4888),
.B2(n_4813),
.Y(n_5343)
);

O2A1O1Ixp33_ASAP7_75t_SL g5344 ( 
.A1(n_5006),
.A2(n_4928),
.B(n_4861),
.C(n_4906),
.Y(n_5344)
);

BUFx10_ASAP7_75t_L g5345 ( 
.A(n_5007),
.Y(n_5345)
);

AO31x2_ASAP7_75t_L g5346 ( 
.A1(n_5234),
.A2(n_4934),
.A3(n_4942),
.B(n_4912),
.Y(n_5346)
);

CKINVDCx11_ASAP7_75t_R g5347 ( 
.A(n_5064),
.Y(n_5347)
);

AND2x4_ASAP7_75t_L g5348 ( 
.A(n_5161),
.B(n_4946),
.Y(n_5348)
);

AOI22xp5_ASAP7_75t_L g5349 ( 
.A1(n_5085),
.A2(n_4828),
.B1(n_4831),
.B2(n_4804),
.Y(n_5349)
);

AND2x2_ASAP7_75t_L g5350 ( 
.A(n_5018),
.B(n_4627),
.Y(n_5350)
);

NOR2xp33_ASAP7_75t_L g5351 ( 
.A(n_5002),
.B(n_4853),
.Y(n_5351)
);

O2A1O1Ixp33_ASAP7_75t_SL g5352 ( 
.A1(n_5040),
.A2(n_4899),
.B(n_4734),
.C(n_4729),
.Y(n_5352)
);

OAI21x1_ASAP7_75t_L g5353 ( 
.A1(n_5073),
.A2(n_5096),
.B(n_5079),
.Y(n_5353)
);

INVx1_ASAP7_75t_SL g5354 ( 
.A(n_5046),
.Y(n_5354)
);

AND2x2_ASAP7_75t_L g5355 ( 
.A(n_4987),
.B(n_4735),
.Y(n_5355)
);

INVx2_ASAP7_75t_L g5356 ( 
.A(n_5004),
.Y(n_5356)
);

NAND2xp33_ASAP7_75t_L g5357 ( 
.A(n_5153),
.B(n_4845),
.Y(n_5357)
);

OR2x6_ASAP7_75t_L g5358 ( 
.A(n_5054),
.B(n_4751),
.Y(n_5358)
);

A2O1A1Ixp33_ASAP7_75t_L g5359 ( 
.A1(n_5177),
.A2(n_4878),
.B(n_4662),
.C(n_4761),
.Y(n_5359)
);

NOR2xp33_ASAP7_75t_L g5360 ( 
.A(n_5002),
.B(n_5067),
.Y(n_5360)
);

INVxp67_ASAP7_75t_SL g5361 ( 
.A(n_5097),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_5057),
.Y(n_5362)
);

A2O1A1Ixp33_ASAP7_75t_L g5363 ( 
.A1(n_5269),
.A2(n_4858),
.B(n_4859),
.C(n_4850),
.Y(n_5363)
);

HB1xp67_ASAP7_75t_L g5364 ( 
.A(n_5090),
.Y(n_5364)
);

NAND2xp5_ASAP7_75t_L g5365 ( 
.A(n_5145),
.B(n_4952),
.Y(n_5365)
);

AO32x2_ASAP7_75t_L g5366 ( 
.A1(n_5108),
.A2(n_4958),
.A3(n_4932),
.B1(n_4719),
.B2(n_4707),
.Y(n_5366)
);

OR2x6_ASAP7_75t_L g5367 ( 
.A(n_5092),
.B(n_4760),
.Y(n_5367)
);

INVx2_ASAP7_75t_SL g5368 ( 
.A(n_5000),
.Y(n_5368)
);

INVx2_ASAP7_75t_L g5369 ( 
.A(n_5019),
.Y(n_5369)
);

O2A1O1Ixp33_ASAP7_75t_SL g5370 ( 
.A1(n_5109),
.A2(n_4867),
.B(n_4972),
.C(n_4764),
.Y(n_5370)
);

O2A1O1Ixp33_ASAP7_75t_SL g5371 ( 
.A1(n_5193),
.A2(n_4777),
.B(n_4756),
.C(n_4545),
.Y(n_5371)
);

INVx2_ASAP7_75t_L g5372 ( 
.A(n_5055),
.Y(n_5372)
);

OAI21x1_ASAP7_75t_L g5373 ( 
.A1(n_5125),
.A2(n_4544),
.B(n_4519),
.Y(n_5373)
);

NAND2x1p5_ASAP7_75t_L g5374 ( 
.A(n_5210),
.B(n_4823),
.Y(n_5374)
);

NOR2x1_ASAP7_75t_SL g5375 ( 
.A(n_5092),
.B(n_4785),
.Y(n_5375)
);

O2A1O1Ixp33_ASAP7_75t_L g5376 ( 
.A1(n_5260),
.A2(n_4955),
.B(n_4978),
.C(n_4953),
.Y(n_5376)
);

AOI22xp33_ASAP7_75t_SL g5377 ( 
.A1(n_5169),
.A2(n_4670),
.B1(n_4875),
.B2(n_4548),
.Y(n_5377)
);

AO31x2_ASAP7_75t_L g5378 ( 
.A1(n_5039),
.A2(n_4585),
.A3(n_4738),
.B(n_4736),
.Y(n_5378)
);

OAI21xp5_ASAP7_75t_L g5379 ( 
.A1(n_5070),
.A2(n_4915),
.B(n_4709),
.Y(n_5379)
);

BUFx3_ASAP7_75t_L g5380 ( 
.A(n_5029),
.Y(n_5380)
);

HB1xp67_ASAP7_75t_L g5381 ( 
.A(n_5118),
.Y(n_5381)
);

A2O1A1Ixp33_ASAP7_75t_L g5382 ( 
.A1(n_5206),
.A2(n_4865),
.B(n_4891),
.C(n_4887),
.Y(n_5382)
);

NOR2xp33_ASAP7_75t_L g5383 ( 
.A(n_5067),
.B(n_4615),
.Y(n_5383)
);

OR2x6_ASAP7_75t_L g5384 ( 
.A(n_5136),
.B(n_4909),
.Y(n_5384)
);

A2O1A1Ixp33_ASAP7_75t_L g5385 ( 
.A1(n_5032),
.A2(n_4893),
.B(n_4732),
.C(n_4803),
.Y(n_5385)
);

INVx1_ASAP7_75t_SL g5386 ( 
.A(n_5016),
.Y(n_5386)
);

INVx2_ASAP7_75t_L g5387 ( 
.A(n_5095),
.Y(n_5387)
);

AOI21xp5_ASAP7_75t_L g5388 ( 
.A1(n_5123),
.A2(n_4573),
.B(n_4618),
.Y(n_5388)
);

AOI221x1_ASAP7_75t_L g5389 ( 
.A1(n_5241),
.A2(n_4740),
.B1(n_4623),
.B2(n_4636),
.C(n_4632),
.Y(n_5389)
);

AOI22xp33_ASAP7_75t_L g5390 ( 
.A1(n_5190),
.A2(n_4560),
.B1(n_4571),
.B2(n_4854),
.Y(n_5390)
);

CKINVDCx5p33_ASAP7_75t_R g5391 ( 
.A(n_5124),
.Y(n_5391)
);

A2O1A1Ixp33_ASAP7_75t_L g5392 ( 
.A1(n_5122),
.A2(n_4812),
.B(n_4816),
.C(n_4797),
.Y(n_5392)
);

NOR2xp33_ASAP7_75t_L g5393 ( 
.A(n_5016),
.B(n_4629),
.Y(n_5393)
);

OAI21xp5_ASAP7_75t_L g5394 ( 
.A1(n_4992),
.A2(n_4630),
.B(n_4835),
.Y(n_5394)
);

INVx2_ASAP7_75t_L g5395 ( 
.A(n_5113),
.Y(n_5395)
);

AOI21xp5_ASAP7_75t_L g5396 ( 
.A1(n_5026),
.A2(n_4646),
.B(n_4648),
.Y(n_5396)
);

AOI21xp5_ASAP7_75t_L g5397 ( 
.A1(n_5146),
.A2(n_4787),
.B(n_4860),
.Y(n_5397)
);

AOI21xp5_ASAP7_75t_L g5398 ( 
.A1(n_5218),
.A2(n_4959),
.B(n_4956),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5072),
.Y(n_5399)
);

AOI21xp5_ASAP7_75t_L g5400 ( 
.A1(n_5051),
.A2(n_4559),
.B(n_4516),
.Y(n_5400)
);

AO31x2_ASAP7_75t_L g5401 ( 
.A1(n_5231),
.A2(n_4651),
.A3(n_4724),
.B(n_4948),
.Y(n_5401)
);

NAND2xp5_ASAP7_75t_L g5402 ( 
.A(n_5138),
.B(n_4728),
.Y(n_5402)
);

NAND2xp33_ASAP7_75t_L g5403 ( 
.A(n_5169),
.B(n_4767),
.Y(n_5403)
);

INVx5_ASAP7_75t_L g5404 ( 
.A(n_5023),
.Y(n_5404)
);

AOI21xp5_ASAP7_75t_L g5405 ( 
.A1(n_5051),
.A2(n_4871),
.B(n_4975),
.Y(n_5405)
);

OAI221xp5_ASAP7_75t_L g5406 ( 
.A1(n_4998),
.A2(n_4808),
.B1(n_4905),
.B2(n_4843),
.C(n_4711),
.Y(n_5406)
);

OA21x2_ASAP7_75t_L g5407 ( 
.A1(n_5009),
.A2(n_5015),
.B(n_5236),
.Y(n_5407)
);

NAND2xp5_ASAP7_75t_L g5408 ( 
.A(n_5132),
.B(n_5227),
.Y(n_5408)
);

OAI22xp5_ASAP7_75t_L g5409 ( 
.A1(n_5122),
.A2(n_4920),
.B1(n_4926),
.B2(n_4907),
.Y(n_5409)
);

O2A1O1Ixp33_ASAP7_75t_SL g5410 ( 
.A1(n_5020),
.A2(n_4938),
.B(n_4941),
.C(n_4929),
.Y(n_5410)
);

AND2x2_ASAP7_75t_L g5411 ( 
.A(n_5045),
.B(n_4654),
.Y(n_5411)
);

INVx8_ASAP7_75t_L g5412 ( 
.A(n_5023),
.Y(n_5412)
);

OR2x6_ASAP7_75t_L g5413 ( 
.A(n_5136),
.B(n_4664),
.Y(n_5413)
);

AOI21x1_ASAP7_75t_L g5414 ( 
.A1(n_5137),
.A2(n_4696),
.B(n_4695),
.Y(n_5414)
);

INVx1_ASAP7_75t_SL g5415 ( 
.A(n_5102),
.Y(n_5415)
);

AOI22xp33_ASAP7_75t_L g5416 ( 
.A1(n_5244),
.A2(n_5238),
.B1(n_5179),
.B2(n_5005),
.Y(n_5416)
);

OAI21xp5_ASAP7_75t_L g5417 ( 
.A1(n_5172),
.A2(n_4587),
.B(n_386),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5077),
.Y(n_5418)
);

O2A1O1Ixp33_ASAP7_75t_SL g5419 ( 
.A1(n_5129),
.A2(n_5275),
.B(n_5213),
.C(n_5192),
.Y(n_5419)
);

OAI22xp5_ASAP7_75t_L g5420 ( 
.A1(n_5188),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_5420)
);

NOR2xp33_ASAP7_75t_L g5421 ( 
.A(n_5239),
.B(n_388),
.Y(n_5421)
);

AOI21xp5_ASAP7_75t_L g5422 ( 
.A1(n_4981),
.A2(n_389),
.B(n_390),
.Y(n_5422)
);

O2A1O1Ixp33_ASAP7_75t_L g5423 ( 
.A1(n_5246),
.A2(n_392),
.B(n_390),
.C(n_391),
.Y(n_5423)
);

AND2x4_ASAP7_75t_L g5424 ( 
.A(n_5063),
.B(n_4983),
.Y(n_5424)
);

O2A1O1Ixp33_ASAP7_75t_SL g5425 ( 
.A1(n_5027),
.A2(n_393),
.B(n_390),
.C(n_391),
.Y(n_5425)
);

INVx2_ASAP7_75t_L g5426 ( 
.A(n_5141),
.Y(n_5426)
);

AND2x4_ASAP7_75t_L g5427 ( 
.A(n_4999),
.B(n_393),
.Y(n_5427)
);

NOR2xp33_ASAP7_75t_L g5428 ( 
.A(n_5156),
.B(n_394),
.Y(n_5428)
);

NAND4xp25_ASAP7_75t_L g5429 ( 
.A(n_5262),
.B(n_396),
.C(n_394),
.D(n_395),
.Y(n_5429)
);

CKINVDCx5p33_ASAP7_75t_R g5430 ( 
.A(n_5134),
.Y(n_5430)
);

AOI31xp67_ASAP7_75t_L g5431 ( 
.A1(n_5277),
.A2(n_396),
.A3(n_394),
.B(n_395),
.Y(n_5431)
);

BUFx3_ASAP7_75t_L g5432 ( 
.A(n_5107),
.Y(n_5432)
);

CKINVDCx5p33_ASAP7_75t_R g5433 ( 
.A(n_5049),
.Y(n_5433)
);

O2A1O1Ixp33_ASAP7_75t_SL g5434 ( 
.A1(n_5143),
.A2(n_399),
.B(n_397),
.C(n_398),
.Y(n_5434)
);

BUFx8_ASAP7_75t_SL g5435 ( 
.A(n_5135),
.Y(n_5435)
);

AO31x2_ASAP7_75t_L g5436 ( 
.A1(n_5176),
.A2(n_399),
.A3(n_397),
.B(n_398),
.Y(n_5436)
);

BUFx2_ASAP7_75t_L g5437 ( 
.A(n_5160),
.Y(n_5437)
);

OAI21x1_ASAP7_75t_L g5438 ( 
.A1(n_5171),
.A2(n_858),
.B(n_857),
.Y(n_5438)
);

AND2x2_ASAP7_75t_L g5439 ( 
.A(n_4982),
.B(n_397),
.Y(n_5439)
);

INVx2_ASAP7_75t_L g5440 ( 
.A(n_5148),
.Y(n_5440)
);

OAI21x1_ASAP7_75t_L g5441 ( 
.A1(n_5233),
.A2(n_860),
.B(n_859),
.Y(n_5441)
);

NOR2xp33_ASAP7_75t_L g5442 ( 
.A(n_5268),
.B(n_398),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5082),
.Y(n_5443)
);

OAI22xp5_ASAP7_75t_L g5444 ( 
.A1(n_5164),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_5444)
);

AOI21xp33_ASAP7_75t_L g5445 ( 
.A1(n_5150),
.A2(n_400),
.B(n_401),
.Y(n_5445)
);

AOI21xp5_ASAP7_75t_L g5446 ( 
.A1(n_5137),
.A2(n_402),
.B(n_403),
.Y(n_5446)
);

AO21x1_ASAP7_75t_L g5447 ( 
.A1(n_5076),
.A2(n_402),
.B(n_404),
.Y(n_5447)
);

AO31x2_ASAP7_75t_L g5448 ( 
.A1(n_5021),
.A2(n_406),
.A3(n_404),
.B(n_405),
.Y(n_5448)
);

BUFx12f_ASAP7_75t_L g5449 ( 
.A(n_5158),
.Y(n_5449)
);

OAI21x1_ASAP7_75t_L g5450 ( 
.A1(n_5048),
.A2(n_862),
.B(n_861),
.Y(n_5450)
);

BUFx2_ASAP7_75t_L g5451 ( 
.A(n_5060),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_L g5452 ( 
.A(n_4985),
.B(n_404),
.Y(n_5452)
);

INVx4_ASAP7_75t_L g5453 ( 
.A(n_5210),
.Y(n_5453)
);

OAI22x1_ASAP7_75t_L g5454 ( 
.A1(n_5078),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_5454)
);

OAI21x1_ASAP7_75t_L g5455 ( 
.A1(n_5126),
.A2(n_863),
.B(n_862),
.Y(n_5455)
);

INVxp67_ASAP7_75t_L g5456 ( 
.A(n_5035),
.Y(n_5456)
);

AOI22xp33_ASAP7_75t_SL g5457 ( 
.A1(n_5169),
.A2(n_408),
.B1(n_405),
.B2(n_407),
.Y(n_5457)
);

AND2x6_ASAP7_75t_L g5458 ( 
.A(n_5168),
.B(n_5173),
.Y(n_5458)
);

AOI21xp5_ASAP7_75t_L g5459 ( 
.A1(n_5130),
.A2(n_408),
.B(n_409),
.Y(n_5459)
);

AOI22xp33_ASAP7_75t_L g5460 ( 
.A1(n_5279),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_5460)
);

AOI21xp5_ASAP7_75t_L g5461 ( 
.A1(n_5232),
.A2(n_409),
.B(n_410),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_5084),
.Y(n_5462)
);

OAI22xp5_ASAP7_75t_L g5463 ( 
.A1(n_5340),
.A2(n_5112),
.B1(n_5202),
.B2(n_5089),
.Y(n_5463)
);

BUFx2_ASAP7_75t_L g5464 ( 
.A(n_5451),
.Y(n_5464)
);

INVx2_ASAP7_75t_L g5465 ( 
.A(n_5320),
.Y(n_5465)
);

AND2x2_ASAP7_75t_L g5466 ( 
.A(n_5290),
.B(n_5104),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_5289),
.Y(n_5467)
);

AND2x2_ASAP7_75t_L g5468 ( 
.A(n_5356),
.B(n_5111),
.Y(n_5468)
);

BUFx3_ASAP7_75t_L g5469 ( 
.A(n_5301),
.Y(n_5469)
);

AO31x2_ASAP7_75t_L g5470 ( 
.A1(n_5331),
.A2(n_5087),
.A3(n_5088),
.B(n_5086),
.Y(n_5470)
);

AOI22xp33_ASAP7_75t_L g5471 ( 
.A1(n_5357),
.A2(n_5265),
.B1(n_5217),
.B2(n_5183),
.Y(n_5471)
);

O2A1O1Ixp33_ASAP7_75t_L g5472 ( 
.A1(n_5288),
.A2(n_5263),
.B(n_5267),
.C(n_5266),
.Y(n_5472)
);

OAI22xp5_ASAP7_75t_L g5473 ( 
.A1(n_5305),
.A2(n_5089),
.B1(n_5235),
.B2(n_5278),
.Y(n_5473)
);

OAI22xp33_ASAP7_75t_L g5474 ( 
.A1(n_5307),
.A2(n_5140),
.B1(n_5207),
.B2(n_5181),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_5294),
.Y(n_5475)
);

OAI22xp5_ASAP7_75t_L g5476 ( 
.A1(n_5354),
.A2(n_5083),
.B1(n_5036),
.B2(n_5219),
.Y(n_5476)
);

AOI22xp5_ASAP7_75t_L g5477 ( 
.A1(n_5429),
.A2(n_5075),
.B1(n_5013),
.B2(n_5091),
.Y(n_5477)
);

BUFx4f_ASAP7_75t_L g5478 ( 
.A(n_5322),
.Y(n_5478)
);

AND2x4_ASAP7_75t_L g5479 ( 
.A(n_5424),
.B(n_5229),
.Y(n_5479)
);

AOI22xp33_ASAP7_75t_L g5480 ( 
.A1(n_5400),
.A2(n_5237),
.B1(n_5251),
.B2(n_5226),
.Y(n_5480)
);

OAI22xp33_ASAP7_75t_L g5481 ( 
.A1(n_5384),
.A2(n_5194),
.B1(n_5187),
.B2(n_5152),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5300),
.Y(n_5482)
);

AND2x2_ASAP7_75t_L g5483 ( 
.A(n_5364),
.B(n_5071),
.Y(n_5483)
);

INVx3_ASAP7_75t_L g5484 ( 
.A(n_5412),
.Y(n_5484)
);

OR2x6_ASAP7_75t_L g5485 ( 
.A(n_5449),
.B(n_5024),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_5369),
.Y(n_5486)
);

INVx1_ASAP7_75t_L g5487 ( 
.A(n_5314),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_5319),
.Y(n_5488)
);

AO31x2_ASAP7_75t_L g5489 ( 
.A1(n_5295),
.A2(n_5099),
.A3(n_5101),
.B(n_5100),
.Y(n_5489)
);

AND3x2_ASAP7_75t_L g5490 ( 
.A(n_5437),
.B(n_5065),
.C(n_5034),
.Y(n_5490)
);

CKINVDCx16_ASAP7_75t_R g5491 ( 
.A(n_5283),
.Y(n_5491)
);

OAI22xp5_ASAP7_75t_L g5492 ( 
.A1(n_5358),
.A2(n_5220),
.B1(n_5157),
.B2(n_4996),
.Y(n_5492)
);

INVx2_ASAP7_75t_SL g5493 ( 
.A(n_5412),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_5372),
.Y(n_5494)
);

BUFx2_ASAP7_75t_L g5495 ( 
.A(n_5458),
.Y(n_5495)
);

INVx4_ASAP7_75t_L g5496 ( 
.A(n_5404),
.Y(n_5496)
);

OAI22xp33_ASAP7_75t_L g5497 ( 
.A1(n_5384),
.A2(n_5255),
.B1(n_5274),
.B2(n_5261),
.Y(n_5497)
);

NOR2xp33_ASAP7_75t_R g5498 ( 
.A(n_5347),
.B(n_5120),
.Y(n_5498)
);

AOI22xp33_ASAP7_75t_L g5499 ( 
.A1(n_5350),
.A2(n_5270),
.B1(n_5249),
.B2(n_5250),
.Y(n_5499)
);

NOR2xp33_ASAP7_75t_L g5500 ( 
.A(n_5336),
.B(n_5117),
.Y(n_5500)
);

AND2x2_ASAP7_75t_L g5501 ( 
.A(n_5381),
.B(n_5103),
.Y(n_5501)
);

OAI22xp5_ASAP7_75t_L g5502 ( 
.A1(n_5358),
.A2(n_5081),
.B1(n_5127),
.B2(n_5204),
.Y(n_5502)
);

INVx4_ASAP7_75t_L g5503 ( 
.A(n_5404),
.Y(n_5503)
);

AOI21xp5_ASAP7_75t_L g5504 ( 
.A1(n_5375),
.A2(n_5240),
.B(n_5230),
.Y(n_5504)
);

INVx2_ASAP7_75t_L g5505 ( 
.A(n_5387),
.Y(n_5505)
);

OAI221xp5_ASAP7_75t_L g5506 ( 
.A1(n_5416),
.A2(n_5271),
.B1(n_5273),
.B2(n_5252),
.C(n_5253),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5334),
.Y(n_5507)
);

AND2x2_ASAP7_75t_L g5508 ( 
.A(n_5361),
.B(n_5105),
.Y(n_5508)
);

INVxp67_ASAP7_75t_SL g5509 ( 
.A(n_5321),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_5395),
.Y(n_5510)
);

INVx2_ASAP7_75t_L g5511 ( 
.A(n_5426),
.Y(n_5511)
);

NOR2x1_ASAP7_75t_L g5512 ( 
.A(n_5380),
.B(n_5247),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5362),
.Y(n_5513)
);

AND2x4_ASAP7_75t_L g5514 ( 
.A(n_5458),
.B(n_5180),
.Y(n_5514)
);

OR2x6_ASAP7_75t_L g5515 ( 
.A(n_5368),
.B(n_5098),
.Y(n_5515)
);

AOI221xp5_ASAP7_75t_L g5516 ( 
.A1(n_5454),
.A2(n_5221),
.B1(n_5264),
.B2(n_4986),
.C(n_5011),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5399),
.Y(n_5517)
);

INVx2_ASAP7_75t_L g5518 ( 
.A(n_5440),
.Y(n_5518)
);

BUFx12f_ASAP7_75t_L g5519 ( 
.A(n_5287),
.Y(n_5519)
);

INVx6_ASAP7_75t_L g5520 ( 
.A(n_5345),
.Y(n_5520)
);

OR2x6_ASAP7_75t_L g5521 ( 
.A(n_5353),
.B(n_5453),
.Y(n_5521)
);

AND2x4_ASAP7_75t_L g5522 ( 
.A(n_5458),
.B(n_5198),
.Y(n_5522)
);

CKINVDCx5p33_ASAP7_75t_R g5523 ( 
.A(n_5435),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_5292),
.Y(n_5524)
);

AND2x2_ASAP7_75t_L g5525 ( 
.A(n_5333),
.B(n_5114),
.Y(n_5525)
);

NAND2xp5_ASAP7_75t_L g5526 ( 
.A(n_5408),
.B(n_5119),
.Y(n_5526)
);

OA21x2_ASAP7_75t_L g5527 ( 
.A1(n_5308),
.A2(n_5324),
.B(n_5373),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5418),
.Y(n_5528)
);

OAI22xp33_ASAP7_75t_L g5529 ( 
.A1(n_5367),
.A2(n_4995),
.B1(n_5259),
.B2(n_5282),
.Y(n_5529)
);

AOI221xp5_ASAP7_75t_L g5530 ( 
.A1(n_5299),
.A2(n_5131),
.B1(n_5254),
.B2(n_5258),
.C(n_5212),
.Y(n_5530)
);

NOR2xp33_ASAP7_75t_L g5531 ( 
.A(n_5336),
.B(n_5128),
.Y(n_5531)
);

AOI22xp33_ASAP7_75t_L g5532 ( 
.A1(n_5403),
.A2(n_5447),
.B1(n_5293),
.B2(n_5411),
.Y(n_5532)
);

NAND2xp33_ASAP7_75t_L g5533 ( 
.A(n_5330),
.B(n_5151),
.Y(n_5533)
);

AOI22xp5_ASAP7_75t_L g5534 ( 
.A1(n_5323),
.A2(n_5200),
.B1(n_5203),
.B2(n_5199),
.Y(n_5534)
);

CKINVDCx20_ASAP7_75t_R g5535 ( 
.A(n_5391),
.Y(n_5535)
);

INVx2_ASAP7_75t_L g5536 ( 
.A(n_5443),
.Y(n_5536)
);

BUFx2_ASAP7_75t_R g5537 ( 
.A(n_5433),
.Y(n_5537)
);

AOI22xp5_ASAP7_75t_L g5538 ( 
.A1(n_5343),
.A2(n_5209),
.B1(n_5166),
.B2(n_5174),
.Y(n_5538)
);

INVx1_ASAP7_75t_SL g5539 ( 
.A(n_5415),
.Y(n_5539)
);

AOI22xp33_ASAP7_75t_L g5540 ( 
.A1(n_5367),
.A2(n_5197),
.B1(n_5211),
.B2(n_5155),
.Y(n_5540)
);

OA21x2_ASAP7_75t_L g5541 ( 
.A1(n_5297),
.A2(n_5318),
.B(n_5339),
.Y(n_5541)
);

AOI22xp33_ASAP7_75t_L g5542 ( 
.A1(n_5390),
.A2(n_5154),
.B1(n_5182),
.B2(n_5149),
.Y(n_5542)
);

INVx2_ASAP7_75t_L g5543 ( 
.A(n_5462),
.Y(n_5543)
);

INVx2_ASAP7_75t_L g5544 ( 
.A(n_5298),
.Y(n_5544)
);

CKINVDCx9p33_ASAP7_75t_R g5545 ( 
.A(n_5421),
.Y(n_5545)
);

BUFx3_ASAP7_75t_L g5546 ( 
.A(n_5330),
.Y(n_5546)
);

AOI21xp5_ASAP7_75t_L g5547 ( 
.A1(n_5337),
.A2(n_5195),
.B(n_5185),
.Y(n_5547)
);

INVx3_ASAP7_75t_L g5548 ( 
.A(n_5296),
.Y(n_5548)
);

NAND2xp5_ASAP7_75t_L g5549 ( 
.A(n_5365),
.B(n_5201),
.Y(n_5549)
);

OAI21xp5_ASAP7_75t_SL g5550 ( 
.A1(n_5325),
.A2(n_5377),
.B(n_5457),
.Y(n_5550)
);

AND2x2_ASAP7_75t_L g5551 ( 
.A(n_5355),
.B(n_5214),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5338),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5302),
.Y(n_5553)
);

INVx2_ASAP7_75t_L g5554 ( 
.A(n_5378),
.Y(n_5554)
);

BUFx2_ASAP7_75t_L g5555 ( 
.A(n_5286),
.Y(n_5555)
);

OAI22xp5_ASAP7_75t_L g5556 ( 
.A1(n_5349),
.A2(n_5216),
.B1(n_5147),
.B2(n_5163),
.Y(n_5556)
);

AOI22xp33_ASAP7_75t_L g5557 ( 
.A1(n_5315),
.A2(n_5422),
.B1(n_5406),
.B2(n_5379),
.Y(n_5557)
);

AND2x2_ASAP7_75t_L g5558 ( 
.A(n_5407),
.B(n_5133),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5303),
.Y(n_5559)
);

HB1xp67_ASAP7_75t_L g5560 ( 
.A(n_5386),
.Y(n_5560)
);

INVx8_ASAP7_75t_L g5561 ( 
.A(n_5430),
.Y(n_5561)
);

AOI222xp33_ASAP7_75t_L g5562 ( 
.A1(n_5444),
.A2(n_5165),
.B1(n_5147),
.B2(n_5170),
.C1(n_5163),
.C2(n_5133),
.Y(n_5562)
);

AOI22xp33_ASAP7_75t_L g5563 ( 
.A1(n_5313),
.A2(n_5170),
.B1(n_5223),
.B2(n_5165),
.Y(n_5563)
);

INVx2_ASAP7_75t_L g5564 ( 
.A(n_5378),
.Y(n_5564)
);

OAI22xp33_ASAP7_75t_L g5565 ( 
.A1(n_5413),
.A2(n_5243),
.B1(n_5245),
.B2(n_5223),
.Y(n_5565)
);

AND2x4_ASAP7_75t_L g5566 ( 
.A(n_5360),
.B(n_5243),
.Y(n_5566)
);

OAI222xp33_ASAP7_75t_L g5567 ( 
.A1(n_5413),
.A2(n_412),
.B1(n_414),
.B2(n_410),
.C1(n_411),
.C2(n_413),
.Y(n_5567)
);

OAI22xp33_ASAP7_75t_L g5568 ( 
.A1(n_5405),
.A2(n_5248),
.B1(n_5280),
.B2(n_5245),
.Y(n_5568)
);

OR2x6_ASAP7_75t_L g5569 ( 
.A(n_5432),
.B(n_5248),
.Y(n_5569)
);

A2O1A1Ixp33_ASAP7_75t_L g5570 ( 
.A1(n_5310),
.A2(n_5285),
.B(n_5423),
.C(n_5446),
.Y(n_5570)
);

INVx5_ASAP7_75t_L g5571 ( 
.A(n_5296),
.Y(n_5571)
);

BUFx6f_ASAP7_75t_L g5572 ( 
.A(n_5427),
.Y(n_5572)
);

O2A1O1Ixp33_ASAP7_75t_SL g5573 ( 
.A1(n_5385),
.A2(n_414),
.B(n_411),
.C(n_412),
.Y(n_5573)
);

AOI21xp33_ASAP7_75t_L g5574 ( 
.A1(n_5309),
.A2(n_5280),
.B(n_411),
.Y(n_5574)
);

AND2x4_ASAP7_75t_L g5575 ( 
.A(n_5348),
.B(n_412),
.Y(n_5575)
);

CKINVDCx6p67_ASAP7_75t_R g5576 ( 
.A(n_5439),
.Y(n_5576)
);

OAI22xp5_ASAP7_75t_L g5577 ( 
.A1(n_5284),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_5577)
);

OAI221xp5_ASAP7_75t_L g5578 ( 
.A1(n_5291),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.C(n_418),
.Y(n_5578)
);

NOR2xp33_ASAP7_75t_L g5579 ( 
.A(n_5419),
.B(n_415),
.Y(n_5579)
);

BUFx2_ASAP7_75t_L g5580 ( 
.A(n_5456),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_5306),
.Y(n_5581)
);

AOI22xp5_ASAP7_75t_L g5582 ( 
.A1(n_5317),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_5582)
);

BUFx12f_ASAP7_75t_L g5583 ( 
.A(n_5316),
.Y(n_5583)
);

AOI22xp33_ASAP7_75t_L g5584 ( 
.A1(n_5394),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_5584)
);

NOR2xp67_ASAP7_75t_L g5585 ( 
.A(n_5304),
.B(n_420),
.Y(n_5585)
);

AOI22xp33_ASAP7_75t_L g5586 ( 
.A1(n_5398),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_5586)
);

AOI22xp33_ASAP7_75t_L g5587 ( 
.A1(n_5409),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5342),
.Y(n_5588)
);

OR2x2_ASAP7_75t_L g5589 ( 
.A(n_5342),
.B(n_421),
.Y(n_5589)
);

INVx2_ASAP7_75t_SL g5590 ( 
.A(n_5351),
.Y(n_5590)
);

INVx1_ASAP7_75t_SL g5591 ( 
.A(n_5393),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5346),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5346),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_5383),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5452),
.Y(n_5595)
);

AO31x2_ASAP7_75t_L g5596 ( 
.A1(n_5588),
.A2(n_5389),
.A3(n_5396),
.B(n_5388),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_5536),
.Y(n_5597)
);

NAND2xp5_ASAP7_75t_SL g5598 ( 
.A(n_5495),
.B(n_5374),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5543),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_5467),
.Y(n_5600)
);

AOI22xp33_ASAP7_75t_SL g5601 ( 
.A1(n_5463),
.A2(n_5464),
.B1(n_5473),
.B2(n_5492),
.Y(n_5601)
);

BUFx2_ASAP7_75t_L g5602 ( 
.A(n_5490),
.Y(n_5602)
);

AND2x2_ASAP7_75t_L g5603 ( 
.A(n_5466),
.B(n_5327),
.Y(n_5603)
);

CKINVDCx14_ASAP7_75t_R g5604 ( 
.A(n_5498),
.Y(n_5604)
);

HB1xp67_ASAP7_75t_L g5605 ( 
.A(n_5580),
.Y(n_5605)
);

NAND2xp5_ASAP7_75t_L g5606 ( 
.A(n_5559),
.B(n_5402),
.Y(n_5606)
);

INVxp67_ASAP7_75t_L g5607 ( 
.A(n_5560),
.Y(n_5607)
);

AOI22xp33_ASAP7_75t_L g5608 ( 
.A1(n_5557),
.A2(n_5420),
.B1(n_5442),
.B2(n_5428),
.Y(n_5608)
);

AO21x2_ASAP7_75t_L g5609 ( 
.A1(n_5592),
.A2(n_5593),
.B(n_5564),
.Y(n_5609)
);

INVx1_ASAP7_75t_L g5610 ( 
.A(n_5475),
.Y(n_5610)
);

OAI21xp5_ASAP7_75t_L g5611 ( 
.A1(n_5472),
.A2(n_5550),
.B(n_5570),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5470),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5482),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5487),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5488),
.Y(n_5615)
);

INVx2_ASAP7_75t_L g5616 ( 
.A(n_5470),
.Y(n_5616)
);

CKINVDCx14_ASAP7_75t_R g5617 ( 
.A(n_5478),
.Y(n_5617)
);

CKINVDCx8_ASAP7_75t_R g5618 ( 
.A(n_5523),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_5507),
.Y(n_5619)
);

BUFx2_ASAP7_75t_L g5620 ( 
.A(n_5521),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_L g5621 ( 
.A(n_5581),
.B(n_5327),
.Y(n_5621)
);

INVxp67_ASAP7_75t_L g5622 ( 
.A(n_5469),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_5513),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5517),
.Y(n_5624)
);

OAI21x1_ASAP7_75t_L g5625 ( 
.A1(n_5558),
.A2(n_5397),
.B(n_5414),
.Y(n_5625)
);

AND2x2_ASAP7_75t_L g5626 ( 
.A(n_5483),
.B(n_5366),
.Y(n_5626)
);

INVx2_ASAP7_75t_L g5627 ( 
.A(n_5486),
.Y(n_5627)
);

OAI21xp5_ASAP7_75t_L g5628 ( 
.A1(n_5532),
.A2(n_5425),
.B(n_5371),
.Y(n_5628)
);

AO21x1_ASAP7_75t_L g5629 ( 
.A1(n_5476),
.A2(n_5461),
.B(n_5311),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_5528),
.Y(n_5630)
);

CKINVDCx5p33_ASAP7_75t_R g5631 ( 
.A(n_5519),
.Y(n_5631)
);

INVx1_ASAP7_75t_L g5632 ( 
.A(n_5552),
.Y(n_5632)
);

BUFx2_ASAP7_75t_L g5633 ( 
.A(n_5521),
.Y(n_5633)
);

BUFx2_ASAP7_75t_L g5634 ( 
.A(n_5515),
.Y(n_5634)
);

HB1xp67_ASAP7_75t_L g5635 ( 
.A(n_5539),
.Y(n_5635)
);

INVx2_ASAP7_75t_SL g5636 ( 
.A(n_5520),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_L g5637 ( 
.A(n_5553),
.B(n_5501),
.Y(n_5637)
);

INVx1_ASAP7_75t_L g5638 ( 
.A(n_5549),
.Y(n_5638)
);

INVx2_ASAP7_75t_L g5639 ( 
.A(n_5494),
.Y(n_5639)
);

INVx2_ASAP7_75t_L g5640 ( 
.A(n_5505),
.Y(n_5640)
);

INVxp67_ASAP7_75t_SL g5641 ( 
.A(n_5533),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_5508),
.Y(n_5642)
);

BUFx4f_ASAP7_75t_SL g5643 ( 
.A(n_5535),
.Y(n_5643)
);

INVx2_ASAP7_75t_L g5644 ( 
.A(n_5510),
.Y(n_5644)
);

OR2x6_ASAP7_75t_L g5645 ( 
.A(n_5485),
.B(n_5341),
.Y(n_5645)
);

INVx1_ASAP7_75t_L g5646 ( 
.A(n_5551),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5525),
.Y(n_5647)
);

INVx3_ASAP7_75t_L g5648 ( 
.A(n_5515),
.Y(n_5648)
);

INVx1_ASAP7_75t_L g5649 ( 
.A(n_5526),
.Y(n_5649)
);

INVx1_ASAP7_75t_L g5650 ( 
.A(n_5524),
.Y(n_5650)
);

HB1xp67_ASAP7_75t_L g5651 ( 
.A(n_5465),
.Y(n_5651)
);

INVx1_ASAP7_75t_L g5652 ( 
.A(n_5511),
.Y(n_5652)
);

BUFx2_ASAP7_75t_L g5653 ( 
.A(n_5569),
.Y(n_5653)
);

INVx3_ASAP7_75t_L g5654 ( 
.A(n_5485),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_5518),
.Y(n_5655)
);

AOI222xp33_ASAP7_75t_L g5656 ( 
.A1(n_5516),
.A2(n_5417),
.B1(n_5460),
.B2(n_5359),
.C1(n_5363),
.C2(n_5366),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_5468),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5544),
.B(n_5328),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_5509),
.Y(n_5659)
);

OR2x2_ASAP7_75t_L g5660 ( 
.A(n_5594),
.B(n_5436),
.Y(n_5660)
);

AO21x2_ASAP7_75t_L g5661 ( 
.A1(n_5554),
.A2(n_5352),
.B(n_5445),
.Y(n_5661)
);

HB1xp67_ASAP7_75t_L g5662 ( 
.A(n_5555),
.Y(n_5662)
);

INVx2_ASAP7_75t_L g5663 ( 
.A(n_5489),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5489),
.Y(n_5664)
);

OAI21x1_ASAP7_75t_L g5665 ( 
.A1(n_5547),
.A2(n_5455),
.B(n_5450),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_5522),
.Y(n_5666)
);

INVx2_ASAP7_75t_L g5667 ( 
.A(n_5541),
.Y(n_5667)
);

INVx2_ASAP7_75t_SL g5668 ( 
.A(n_5520),
.Y(n_5668)
);

INVx3_ASAP7_75t_L g5669 ( 
.A(n_5496),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_5589),
.Y(n_5670)
);

AND2x2_ASAP7_75t_L g5671 ( 
.A(n_5590),
.B(n_5328),
.Y(n_5671)
);

AND2x4_ASAP7_75t_SL g5672 ( 
.A(n_5503),
.B(n_5329),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_5595),
.Y(n_5673)
);

OR2x6_ASAP7_75t_L g5674 ( 
.A(n_5569),
.B(n_5459),
.Y(n_5674)
);

INVx2_ASAP7_75t_L g5675 ( 
.A(n_5479),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5538),
.Y(n_5676)
);

INVx4_ASAP7_75t_L g5677 ( 
.A(n_5571),
.Y(n_5677)
);

INVx2_ASAP7_75t_L g5678 ( 
.A(n_5512),
.Y(n_5678)
);

BUFx3_ASAP7_75t_L g5679 ( 
.A(n_5546),
.Y(n_5679)
);

INVx5_ASAP7_75t_L g5680 ( 
.A(n_5571),
.Y(n_5680)
);

AO21x2_ASAP7_75t_L g5681 ( 
.A1(n_5497),
.A2(n_5434),
.B(n_5332),
.Y(n_5681)
);

NOR2xp33_ASAP7_75t_L g5682 ( 
.A(n_5491),
.B(n_5583),
.Y(n_5682)
);

BUFx3_ASAP7_75t_L g5683 ( 
.A(n_5561),
.Y(n_5683)
);

INVx2_ASAP7_75t_L g5684 ( 
.A(n_5514),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_5534),
.Y(n_5685)
);

INVx2_ASAP7_75t_L g5686 ( 
.A(n_5566),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5502),
.Y(n_5687)
);

OAI21x1_ASAP7_75t_L g5688 ( 
.A1(n_5527),
.A2(n_5441),
.B(n_5438),
.Y(n_5688)
);

INVx2_ASAP7_75t_SL g5689 ( 
.A(n_5493),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_5556),
.Y(n_5690)
);

OAI21x1_ASAP7_75t_L g5691 ( 
.A1(n_5540),
.A2(n_5326),
.B(n_5376),
.Y(n_5691)
);

INVxp67_ASAP7_75t_SL g5692 ( 
.A(n_5585),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5591),
.Y(n_5693)
);

INVx2_ASAP7_75t_SL g5694 ( 
.A(n_5561),
.Y(n_5694)
);

INVx2_ASAP7_75t_L g5695 ( 
.A(n_5572),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_5542),
.Y(n_5696)
);

OA21x2_ASAP7_75t_L g5697 ( 
.A1(n_5480),
.A2(n_5382),
.B(n_5392),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5481),
.Y(n_5698)
);

INVx2_ASAP7_75t_L g5699 ( 
.A(n_5572),
.Y(n_5699)
);

INVx3_ASAP7_75t_L g5700 ( 
.A(n_5484),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_5576),
.Y(n_5701)
);

INVx2_ASAP7_75t_L g5702 ( 
.A(n_5575),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5531),
.Y(n_5703)
);

HB1xp67_ASAP7_75t_L g5704 ( 
.A(n_5548),
.Y(n_5704)
);

OAI21x1_ASAP7_75t_L g5705 ( 
.A1(n_5504),
.A2(n_5312),
.B(n_5431),
.Y(n_5705)
);

AND2x2_ASAP7_75t_L g5706 ( 
.A(n_5471),
.B(n_5563),
.Y(n_5706)
);

INVx8_ASAP7_75t_L g5707 ( 
.A(n_5537),
.Y(n_5707)
);

INVx3_ASAP7_75t_L g5708 ( 
.A(n_5565),
.Y(n_5708)
);

AND2x2_ASAP7_75t_L g5709 ( 
.A(n_5634),
.B(n_5500),
.Y(n_5709)
);

INVx1_ASAP7_75t_L g5710 ( 
.A(n_5605),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5597),
.Y(n_5711)
);

AOI211xp5_ASAP7_75t_L g5712 ( 
.A1(n_5611),
.A2(n_5629),
.B(n_5602),
.C(n_5628),
.Y(n_5712)
);

AND2x4_ASAP7_75t_L g5713 ( 
.A(n_5634),
.B(n_5477),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_5648),
.B(n_5562),
.Y(n_5714)
);

INVx1_ASAP7_75t_L g5715 ( 
.A(n_5599),
.Y(n_5715)
);

AOI22xp33_ASAP7_75t_SL g5716 ( 
.A1(n_5602),
.A2(n_5579),
.B1(n_5506),
.B2(n_5577),
.Y(n_5716)
);

AND2x2_ASAP7_75t_L g5717 ( 
.A(n_5648),
.B(n_5499),
.Y(n_5717)
);

INVx8_ASAP7_75t_L g5718 ( 
.A(n_5680),
.Y(n_5718)
);

INVx5_ASAP7_75t_SL g5719 ( 
.A(n_5617),
.Y(n_5719)
);

OAI22xp5_ASAP7_75t_L g5720 ( 
.A1(n_5601),
.A2(n_5529),
.B1(n_5474),
.B2(n_5568),
.Y(n_5720)
);

AOI21x1_ASAP7_75t_L g5721 ( 
.A1(n_5645),
.A2(n_5545),
.B(n_5567),
.Y(n_5721)
);

INVx1_ASAP7_75t_L g5722 ( 
.A(n_5600),
.Y(n_5722)
);

AOI22xp33_ASAP7_75t_L g5723 ( 
.A1(n_5626),
.A2(n_5574),
.B1(n_5578),
.B2(n_5530),
.Y(n_5723)
);

AND2x2_ASAP7_75t_L g5724 ( 
.A(n_5698),
.B(n_5401),
.Y(n_5724)
);

AOI31xp33_ASAP7_75t_L g5725 ( 
.A1(n_5604),
.A2(n_5573),
.A3(n_5584),
.B(n_5344),
.Y(n_5725)
);

OAI221xp5_ASAP7_75t_L g5726 ( 
.A1(n_5645),
.A2(n_5656),
.B1(n_5692),
.B2(n_5633),
.C(n_5620),
.Y(n_5726)
);

AOI22xp33_ASAP7_75t_L g5727 ( 
.A1(n_5687),
.A2(n_5587),
.B1(n_5586),
.B2(n_5582),
.Y(n_5727)
);

AOI21xp33_ASAP7_75t_L g5728 ( 
.A1(n_5674),
.A2(n_5681),
.B(n_5661),
.Y(n_5728)
);

AOI22xp33_ASAP7_75t_SL g5729 ( 
.A1(n_5620),
.A2(n_5370),
.B1(n_5436),
.B2(n_5448),
.Y(n_5729)
);

OR2x6_ASAP7_75t_L g5730 ( 
.A(n_5677),
.B(n_5448),
.Y(n_5730)
);

NAND2x1_ASAP7_75t_L g5731 ( 
.A(n_5633),
.B(n_5410),
.Y(n_5731)
);

INVx4_ASAP7_75t_L g5732 ( 
.A(n_5680),
.Y(n_5732)
);

AOI211xp5_ASAP7_75t_L g5733 ( 
.A1(n_5682),
.A2(n_5335),
.B(n_5401),
.C(n_425),
.Y(n_5733)
);

OAI22xp5_ASAP7_75t_L g5734 ( 
.A1(n_5653),
.A2(n_5335),
.B1(n_425),
.B2(n_423),
.Y(n_5734)
);

AOI22xp33_ASAP7_75t_SL g5735 ( 
.A1(n_5641),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_5735)
);

BUFx6f_ASAP7_75t_L g5736 ( 
.A(n_5618),
.Y(n_5736)
);

NAND2xp5_ASAP7_75t_L g5737 ( 
.A(n_5696),
.B(n_424),
.Y(n_5737)
);

BUFx2_ASAP7_75t_L g5738 ( 
.A(n_5679),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_5610),
.Y(n_5739)
);

NOR2x1_ASAP7_75t_L g5740 ( 
.A(n_5677),
.B(n_424),
.Y(n_5740)
);

HB1xp67_ASAP7_75t_L g5741 ( 
.A(n_5651),
.Y(n_5741)
);

AND2x2_ASAP7_75t_SL g5742 ( 
.A(n_5653),
.B(n_426),
.Y(n_5742)
);

NAND2xp5_ASAP7_75t_L g5743 ( 
.A(n_5670),
.B(n_426),
.Y(n_5743)
);

AOI222xp33_ASAP7_75t_L g5744 ( 
.A1(n_5608),
.A2(n_429),
.B1(n_431),
.B2(n_427),
.C1(n_428),
.C2(n_430),
.Y(n_5744)
);

CKINVDCx8_ASAP7_75t_R g5745 ( 
.A(n_5707),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5613),
.Y(n_5746)
);

AND2x2_ASAP7_75t_L g5747 ( 
.A(n_5690),
.B(n_427),
.Y(n_5747)
);

AOI21xp5_ASAP7_75t_L g5748 ( 
.A1(n_5598),
.A2(n_427),
.B(n_428),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5614),
.Y(n_5749)
);

AOI22xp33_ASAP7_75t_SL g5750 ( 
.A1(n_5697),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_5750)
);

INVx1_ASAP7_75t_L g5751 ( 
.A(n_5615),
.Y(n_5751)
);

OAI22xp5_ASAP7_75t_L g5752 ( 
.A1(n_5654),
.A2(n_434),
.B1(n_431),
.B2(n_432),
.Y(n_5752)
);

OAI22xp5_ASAP7_75t_L g5753 ( 
.A1(n_5662),
.A2(n_435),
.B1(n_432),
.B2(n_434),
.Y(n_5753)
);

AOI222xp33_ASAP7_75t_L g5754 ( 
.A1(n_5685),
.A2(n_435),
.B1(n_437),
.B2(n_432),
.C1(n_434),
.C2(n_436),
.Y(n_5754)
);

AOI222xp33_ASAP7_75t_L g5755 ( 
.A1(n_5707),
.A2(n_437),
.B1(n_439),
.B2(n_435),
.C1(n_436),
.C2(n_438),
.Y(n_5755)
);

OAI21xp5_ASAP7_75t_L g5756 ( 
.A1(n_5691),
.A2(n_437),
.B(n_438),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5619),
.Y(n_5757)
);

NAND2xp5_ASAP7_75t_L g5758 ( 
.A(n_5676),
.B(n_438),
.Y(n_5758)
);

AOI22xp33_ASAP7_75t_SL g5759 ( 
.A1(n_5697),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_5759)
);

AND2x4_ASAP7_75t_L g5760 ( 
.A(n_5678),
.B(n_439),
.Y(n_5760)
);

AOI22xp33_ASAP7_75t_L g5761 ( 
.A1(n_5674),
.A2(n_443),
.B1(n_440),
.B2(n_442),
.Y(n_5761)
);

AND2x2_ASAP7_75t_L g5762 ( 
.A(n_5706),
.B(n_443),
.Y(n_5762)
);

AO21x2_ASAP7_75t_L g5763 ( 
.A1(n_5667),
.A2(n_443),
.B(n_444),
.Y(n_5763)
);

INVx2_ASAP7_75t_SL g5764 ( 
.A(n_5683),
.Y(n_5764)
);

INVx2_ASAP7_75t_L g5765 ( 
.A(n_5627),
.Y(n_5765)
);

OAI22xp5_ASAP7_75t_L g5766 ( 
.A1(n_5622),
.A2(n_5708),
.B1(n_5669),
.B2(n_5680),
.Y(n_5766)
);

AOI22xp33_ASAP7_75t_L g5767 ( 
.A1(n_5603),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_5767)
);

INVx1_ASAP7_75t_L g5768 ( 
.A(n_5623),
.Y(n_5768)
);

OAI22xp5_ASAP7_75t_L g5769 ( 
.A1(n_5708),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_5769)
);

OAI22xp5_ASAP7_75t_L g5770 ( 
.A1(n_5635),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_5770)
);

OAI221xp5_ASAP7_75t_L g5771 ( 
.A1(n_5621),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.C(n_450),
.Y(n_5771)
);

AOI22xp33_ASAP7_75t_L g5772 ( 
.A1(n_5671),
.A2(n_450),
.B1(n_447),
.B2(n_449),
.Y(n_5772)
);

OAI221xp5_ASAP7_75t_L g5773 ( 
.A1(n_5607),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.C(n_452),
.Y(n_5773)
);

OAI22xp5_ASAP7_75t_L g5774 ( 
.A1(n_5689),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5624),
.Y(n_5775)
);

NAND3xp33_ASAP7_75t_L g5776 ( 
.A(n_5664),
.B(n_452),
.C(n_453),
.Y(n_5776)
);

CKINVDCx11_ASAP7_75t_R g5777 ( 
.A(n_5701),
.Y(n_5777)
);

AOI22xp5_ASAP7_75t_L g5778 ( 
.A1(n_5693),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_5778)
);

OR2x2_ASAP7_75t_L g5779 ( 
.A(n_5606),
.B(n_455),
.Y(n_5779)
);

OAI22xp5_ASAP7_75t_L g5780 ( 
.A1(n_5700),
.A2(n_458),
.B1(n_455),
.B2(n_456),
.Y(n_5780)
);

A2O1A1Ixp33_ASAP7_75t_L g5781 ( 
.A1(n_5672),
.A2(n_5694),
.B(n_5636),
.C(n_5668),
.Y(n_5781)
);

AOI22xp33_ASAP7_75t_L g5782 ( 
.A1(n_5647),
.A2(n_459),
.B1(n_456),
.B2(n_458),
.Y(n_5782)
);

INVx2_ASAP7_75t_L g5783 ( 
.A(n_5639),
.Y(n_5783)
);

AOI22xp33_ASAP7_75t_L g5784 ( 
.A1(n_5642),
.A2(n_460),
.B1(n_456),
.B2(n_459),
.Y(n_5784)
);

INVx2_ASAP7_75t_L g5785 ( 
.A(n_5640),
.Y(n_5785)
);

HB1xp67_ASAP7_75t_L g5786 ( 
.A(n_5659),
.Y(n_5786)
);

INVx2_ASAP7_75t_L g5787 ( 
.A(n_5644),
.Y(n_5787)
);

AOI22xp33_ASAP7_75t_L g5788 ( 
.A1(n_5703),
.A2(n_5702),
.B1(n_5658),
.B2(n_5705),
.Y(n_5788)
);

CKINVDCx20_ASAP7_75t_R g5789 ( 
.A(n_5643),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_5630),
.Y(n_5790)
);

HB1xp67_ASAP7_75t_L g5791 ( 
.A(n_5650),
.Y(n_5791)
);

OAI33xp33_ASAP7_75t_L g5792 ( 
.A1(n_5660),
.A2(n_5649),
.A3(n_5673),
.B1(n_5632),
.B2(n_5638),
.B3(n_5637),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_5652),
.Y(n_5793)
);

INVx2_ASAP7_75t_L g5794 ( 
.A(n_5741),
.Y(n_5794)
);

OR2x2_ASAP7_75t_L g5795 ( 
.A(n_5710),
.B(n_5596),
.Y(n_5795)
);

BUFx6f_ASAP7_75t_L g5796 ( 
.A(n_5736),
.Y(n_5796)
);

AND2x4_ASAP7_75t_L g5797 ( 
.A(n_5781),
.B(n_5704),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5786),
.Y(n_5798)
);

INVx2_ASAP7_75t_L g5799 ( 
.A(n_5791),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_5722),
.Y(n_5800)
);

AND2x2_ASAP7_75t_L g5801 ( 
.A(n_5714),
.B(n_5666),
.Y(n_5801)
);

INVx2_ASAP7_75t_L g5802 ( 
.A(n_5738),
.Y(n_5802)
);

AND2x2_ASAP7_75t_L g5803 ( 
.A(n_5709),
.B(n_5684),
.Y(n_5803)
);

BUFx2_ASAP7_75t_L g5804 ( 
.A(n_5732),
.Y(n_5804)
);

INVx1_ASAP7_75t_L g5805 ( 
.A(n_5739),
.Y(n_5805)
);

INVx1_ASAP7_75t_L g5806 ( 
.A(n_5746),
.Y(n_5806)
);

HB1xp67_ASAP7_75t_L g5807 ( 
.A(n_5793),
.Y(n_5807)
);

HB1xp67_ASAP7_75t_L g5808 ( 
.A(n_5711),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5749),
.Y(n_5809)
);

AND2x4_ASAP7_75t_L g5810 ( 
.A(n_5764),
.B(n_5695),
.Y(n_5810)
);

AND2x2_ASAP7_75t_L g5811 ( 
.A(n_5717),
.B(n_5699),
.Y(n_5811)
);

OR2x2_ASAP7_75t_L g5812 ( 
.A(n_5713),
.B(n_5596),
.Y(n_5812)
);

AND2x2_ASAP7_75t_L g5813 ( 
.A(n_5766),
.B(n_5625),
.Y(n_5813)
);

INVx1_ASAP7_75t_SL g5814 ( 
.A(n_5777),
.Y(n_5814)
);

HB1xp67_ASAP7_75t_L g5815 ( 
.A(n_5715),
.Y(n_5815)
);

NOR2xp33_ASAP7_75t_L g5816 ( 
.A(n_5745),
.B(n_5631),
.Y(n_5816)
);

AOI22xp33_ASAP7_75t_L g5817 ( 
.A1(n_5726),
.A2(n_5686),
.B1(n_5675),
.B2(n_5657),
.Y(n_5817)
);

OAI221xp5_ASAP7_75t_L g5818 ( 
.A1(n_5712),
.A2(n_5612),
.B1(n_5616),
.B2(n_5663),
.C(n_5646),
.Y(n_5818)
);

INVx1_ASAP7_75t_L g5819 ( 
.A(n_5751),
.Y(n_5819)
);

INVx3_ASAP7_75t_L g5820 ( 
.A(n_5719),
.Y(n_5820)
);

AND2x2_ASAP7_75t_L g5821 ( 
.A(n_5724),
.B(n_5788),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5757),
.Y(n_5822)
);

HB1xp67_ASAP7_75t_L g5823 ( 
.A(n_5763),
.Y(n_5823)
);

AND2x2_ASAP7_75t_L g5824 ( 
.A(n_5747),
.B(n_5596),
.Y(n_5824)
);

AND2x2_ASAP7_75t_L g5825 ( 
.A(n_5721),
.B(n_5609),
.Y(n_5825)
);

OR2x2_ASAP7_75t_L g5826 ( 
.A(n_5737),
.B(n_5655),
.Y(n_5826)
);

AND2x4_ASAP7_75t_L g5827 ( 
.A(n_5736),
.B(n_5688),
.Y(n_5827)
);

AO21x2_ASAP7_75t_L g5828 ( 
.A1(n_5728),
.A2(n_5665),
.B(n_459),
.Y(n_5828)
);

BUFx4f_ASAP7_75t_L g5829 ( 
.A(n_5718),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5768),
.Y(n_5830)
);

AO21x2_ASAP7_75t_L g5831 ( 
.A1(n_5756),
.A2(n_461),
.B(n_462),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5775),
.Y(n_5832)
);

NAND2xp5_ASAP7_75t_L g5833 ( 
.A(n_5723),
.B(n_461),
.Y(n_5833)
);

NAND2xp5_ASAP7_75t_L g5834 ( 
.A(n_5729),
.B(n_461),
.Y(n_5834)
);

BUFx2_ASAP7_75t_L g5835 ( 
.A(n_5718),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5790),
.Y(n_5836)
);

INVx3_ASAP7_75t_L g5837 ( 
.A(n_5719),
.Y(n_5837)
);

INVx2_ASAP7_75t_SL g5838 ( 
.A(n_5789),
.Y(n_5838)
);

NAND2x1p5_ASAP7_75t_L g5839 ( 
.A(n_5740),
.B(n_463),
.Y(n_5839)
);

AND2x2_ASAP7_75t_L g5840 ( 
.A(n_5762),
.B(n_462),
.Y(n_5840)
);

INVx2_ASAP7_75t_L g5841 ( 
.A(n_5765),
.Y(n_5841)
);

BUFx2_ASAP7_75t_L g5842 ( 
.A(n_5760),
.Y(n_5842)
);

INVx2_ASAP7_75t_L g5843 ( 
.A(n_5783),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5758),
.Y(n_5844)
);

NAND2xp5_ASAP7_75t_L g5845 ( 
.A(n_5716),
.B(n_463),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_5760),
.Y(n_5846)
);

BUFx6f_ASAP7_75t_L g5847 ( 
.A(n_5742),
.Y(n_5847)
);

BUFx3_ASAP7_75t_L g5848 ( 
.A(n_5743),
.Y(n_5848)
);

INVx1_ASAP7_75t_SL g5849 ( 
.A(n_5779),
.Y(n_5849)
);

OR2x2_ASAP7_75t_L g5850 ( 
.A(n_5785),
.B(n_463),
.Y(n_5850)
);

INVx2_ASAP7_75t_L g5851 ( 
.A(n_5787),
.Y(n_5851)
);

AND2x4_ASAP7_75t_L g5852 ( 
.A(n_5730),
.B(n_464),
.Y(n_5852)
);

HB1xp67_ASAP7_75t_L g5853 ( 
.A(n_5769),
.Y(n_5853)
);

NOR2xp33_ASAP7_75t_L g5854 ( 
.A(n_5792),
.B(n_464),
.Y(n_5854)
);

BUFx3_ASAP7_75t_L g5855 ( 
.A(n_5730),
.Y(n_5855)
);

BUFx3_ASAP7_75t_L g5856 ( 
.A(n_5731),
.Y(n_5856)
);

INVx2_ASAP7_75t_L g5857 ( 
.A(n_5776),
.Y(n_5857)
);

HB1xp67_ASAP7_75t_L g5858 ( 
.A(n_5720),
.Y(n_5858)
);

INVx2_ASAP7_75t_L g5859 ( 
.A(n_5771),
.Y(n_5859)
);

OR2x2_ASAP7_75t_L g5860 ( 
.A(n_5772),
.B(n_464),
.Y(n_5860)
);

NAND2x1p5_ASAP7_75t_L g5861 ( 
.A(n_5748),
.B(n_5778),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_5734),
.Y(n_5862)
);

HB1xp67_ASAP7_75t_L g5863 ( 
.A(n_5774),
.Y(n_5863)
);

AND2x2_ASAP7_75t_L g5864 ( 
.A(n_5761),
.B(n_465),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5753),
.Y(n_5865)
);

NAND2xp5_ASAP7_75t_L g5866 ( 
.A(n_5733),
.B(n_465),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5727),
.Y(n_5867)
);

AOI21xp33_ASAP7_75t_L g5868 ( 
.A1(n_5725),
.A2(n_466),
.B(n_467),
.Y(n_5868)
);

AND2x4_ASAP7_75t_L g5869 ( 
.A(n_5767),
.B(n_466),
.Y(n_5869)
);

NAND2xp5_ASAP7_75t_L g5870 ( 
.A(n_5750),
.B(n_466),
.Y(n_5870)
);

AND2x4_ASAP7_75t_L g5871 ( 
.A(n_5784),
.B(n_467),
.Y(n_5871)
);

OR2x2_ASAP7_75t_SL g5872 ( 
.A(n_5759),
.B(n_467),
.Y(n_5872)
);

OR2x2_ASAP7_75t_L g5873 ( 
.A(n_5770),
.B(n_468),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5752),
.Y(n_5874)
);

NAND2xp5_ASAP7_75t_L g5875 ( 
.A(n_5754),
.B(n_469),
.Y(n_5875)
);

OR2x2_ASAP7_75t_L g5876 ( 
.A(n_5780),
.B(n_469),
.Y(n_5876)
);

INVx1_ASAP7_75t_L g5877 ( 
.A(n_5735),
.Y(n_5877)
);

AND2x4_ASAP7_75t_L g5878 ( 
.A(n_5782),
.B(n_469),
.Y(n_5878)
);

NAND2xp5_ASAP7_75t_L g5879 ( 
.A(n_5755),
.B(n_470),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5773),
.Y(n_5880)
);

HB1xp67_ASAP7_75t_L g5881 ( 
.A(n_5744),
.Y(n_5881)
);

HB1xp67_ASAP7_75t_L g5882 ( 
.A(n_5741),
.Y(n_5882)
);

OAI21x1_ASAP7_75t_L g5883 ( 
.A1(n_5766),
.A2(n_470),
.B(n_471),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5786),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5786),
.Y(n_5885)
);

AND2x2_ASAP7_75t_L g5886 ( 
.A(n_5797),
.B(n_471),
.Y(n_5886)
);

INVx2_ASAP7_75t_L g5887 ( 
.A(n_5802),
.Y(n_5887)
);

AOI22xp33_ASAP7_75t_L g5888 ( 
.A1(n_5858),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_5888)
);

AOI221xp5_ASAP7_75t_L g5889 ( 
.A1(n_5868),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.C(n_475),
.Y(n_5889)
);

AOI33xp33_ASAP7_75t_L g5890 ( 
.A1(n_5867),
.A2(n_475),
.A3(n_477),
.B1(n_473),
.B2(n_474),
.B3(n_476),
.Y(n_5890)
);

NAND3xp33_ASAP7_75t_L g5891 ( 
.A(n_5854),
.B(n_476),
.C(n_477),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5882),
.Y(n_5892)
);

INVx2_ASAP7_75t_L g5893 ( 
.A(n_5794),
.Y(n_5893)
);

INVx1_ASAP7_75t_L g5894 ( 
.A(n_5826),
.Y(n_5894)
);

AOI221xp5_ASAP7_75t_L g5895 ( 
.A1(n_5881),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.C(n_479),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_5798),
.Y(n_5896)
);

OAI21xp5_ASAP7_75t_L g5897 ( 
.A1(n_5852),
.A2(n_478),
.B(n_479),
.Y(n_5897)
);

INVx2_ASAP7_75t_L g5898 ( 
.A(n_5804),
.Y(n_5898)
);

INVx1_ASAP7_75t_SL g5899 ( 
.A(n_5814),
.Y(n_5899)
);

AOI21xp5_ASAP7_75t_L g5900 ( 
.A1(n_5829),
.A2(n_479),
.B(n_480),
.Y(n_5900)
);

OAI22xp33_ASAP7_75t_L g5901 ( 
.A1(n_5856),
.A2(n_5855),
.B1(n_5842),
.B2(n_5812),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5884),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5885),
.Y(n_5903)
);

AOI22xp33_ASAP7_75t_SL g5904 ( 
.A1(n_5797),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_5904)
);

NOR2x1p5_ASAP7_75t_L g5905 ( 
.A(n_5820),
.B(n_480),
.Y(n_5905)
);

AOI22xp33_ASAP7_75t_L g5906 ( 
.A1(n_5821),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_5906)
);

AOI31xp33_ASAP7_75t_L g5907 ( 
.A1(n_5839),
.A2(n_485),
.A3(n_483),
.B(n_484),
.Y(n_5907)
);

AND2x2_ASAP7_75t_L g5908 ( 
.A(n_5835),
.B(n_483),
.Y(n_5908)
);

OAI322xp33_ASAP7_75t_L g5909 ( 
.A1(n_5845),
.A2(n_5834),
.A3(n_5862),
.B1(n_5877),
.B2(n_5853),
.C1(n_5865),
.C2(n_5833),
.Y(n_5909)
);

NAND4xp25_ASAP7_75t_SL g5910 ( 
.A(n_5817),
.B(n_5825),
.C(n_5813),
.D(n_5874),
.Y(n_5910)
);

AOI22xp33_ASAP7_75t_L g5911 ( 
.A1(n_5863),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_5911)
);

NAND2xp5_ASAP7_75t_L g5912 ( 
.A(n_5824),
.B(n_484),
.Y(n_5912)
);

AND2x2_ASAP7_75t_L g5913 ( 
.A(n_5835),
.B(n_485),
.Y(n_5913)
);

AND2x2_ASAP7_75t_L g5914 ( 
.A(n_5801),
.B(n_487),
.Y(n_5914)
);

AOI221xp5_ASAP7_75t_SL g5915 ( 
.A1(n_5872),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.C(n_490),
.Y(n_5915)
);

AND2x2_ASAP7_75t_L g5916 ( 
.A(n_5804),
.B(n_488),
.Y(n_5916)
);

CKINVDCx5p33_ASAP7_75t_R g5917 ( 
.A(n_5816),
.Y(n_5917)
);

OAI222xp33_ASAP7_75t_L g5918 ( 
.A1(n_5818),
.A2(n_490),
.B1(n_492),
.B2(n_488),
.C1(n_489),
.C2(n_491),
.Y(n_5918)
);

HB1xp67_ASAP7_75t_L g5919 ( 
.A(n_5807),
.Y(n_5919)
);

OAI33xp33_ASAP7_75t_L g5920 ( 
.A1(n_5880),
.A2(n_492),
.A3(n_494),
.B1(n_490),
.B2(n_491),
.B3(n_493),
.Y(n_5920)
);

OAI31xp33_ASAP7_75t_SL g5921 ( 
.A1(n_5852),
.A2(n_493),
.A3(n_491),
.B(n_492),
.Y(n_5921)
);

AOI22xp33_ASAP7_75t_L g5922 ( 
.A1(n_5847),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_5922)
);

AND2x2_ASAP7_75t_L g5923 ( 
.A(n_5811),
.B(n_494),
.Y(n_5923)
);

OAI33xp33_ASAP7_75t_L g5924 ( 
.A1(n_5879),
.A2(n_497),
.A3(n_499),
.B1(n_495),
.B2(n_496),
.B3(n_498),
.Y(n_5924)
);

INVx2_ASAP7_75t_SL g5925 ( 
.A(n_5837),
.Y(n_5925)
);

AOI22xp5_ASAP7_75t_L g5926 ( 
.A1(n_5847),
.A2(n_497),
.B1(n_495),
.B2(n_496),
.Y(n_5926)
);

AOI22xp33_ASAP7_75t_L g5927 ( 
.A1(n_5859),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.Y(n_5927)
);

AO31x2_ASAP7_75t_L g5928 ( 
.A1(n_5857),
.A2(n_5842),
.A3(n_5844),
.B(n_5799),
.Y(n_5928)
);

NAND2xp5_ASAP7_75t_SL g5929 ( 
.A(n_5827),
.B(n_498),
.Y(n_5929)
);

INVx4_ASAP7_75t_L g5930 ( 
.A(n_5796),
.Y(n_5930)
);

AND2x2_ASAP7_75t_L g5931 ( 
.A(n_5810),
.B(n_5803),
.Y(n_5931)
);

AOI22xp33_ASAP7_75t_L g5932 ( 
.A1(n_5848),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_5932)
);

OA222x2_ASAP7_75t_L g5933 ( 
.A1(n_5846),
.A2(n_503),
.B1(n_505),
.B2(n_501),
.C1(n_502),
.C2(n_504),
.Y(n_5933)
);

AOI22xp33_ASAP7_75t_L g5934 ( 
.A1(n_5828),
.A2(n_504),
.B1(n_501),
.B2(n_503),
.Y(n_5934)
);

AOI22xp33_ASAP7_75t_SL g5935 ( 
.A1(n_5823),
.A2(n_506),
.B1(n_503),
.B2(n_505),
.Y(n_5935)
);

BUFx2_ASAP7_75t_L g5936 ( 
.A(n_5796),
.Y(n_5936)
);

AOI31xp33_ASAP7_75t_L g5937 ( 
.A1(n_5861),
.A2(n_508),
.A3(n_505),
.B(n_507),
.Y(n_5937)
);

AOI22xp33_ASAP7_75t_L g5938 ( 
.A1(n_5849),
.A2(n_5838),
.B1(n_5869),
.B2(n_5808),
.Y(n_5938)
);

AOI22xp33_ASAP7_75t_L g5939 ( 
.A1(n_5869),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.Y(n_5939)
);

HB1xp67_ASAP7_75t_L g5940 ( 
.A(n_5815),
.Y(n_5940)
);

NOR2xp33_ASAP7_75t_L g5941 ( 
.A(n_5866),
.B(n_507),
.Y(n_5941)
);

OR2x2_ASAP7_75t_L g5942 ( 
.A(n_5795),
.B(n_508),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5800),
.Y(n_5943)
);

OAI211xp5_ASAP7_75t_SL g5944 ( 
.A1(n_5875),
.A2(n_512),
.B(n_510),
.C(n_511),
.Y(n_5944)
);

OAI22xp5_ASAP7_75t_L g5945 ( 
.A1(n_5850),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_5945)
);

AOI21xp5_ASAP7_75t_SL g5946 ( 
.A1(n_5831),
.A2(n_510),
.B(n_511),
.Y(n_5946)
);

AND2x2_ASAP7_75t_L g5947 ( 
.A(n_5841),
.B(n_513),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_5805),
.Y(n_5948)
);

INVx5_ASAP7_75t_L g5949 ( 
.A(n_5864),
.Y(n_5949)
);

AOI322xp5_ASAP7_75t_L g5950 ( 
.A1(n_5840),
.A2(n_518),
.A3(n_517),
.B1(n_515),
.B2(n_513),
.C1(n_514),
.C2(n_516),
.Y(n_5950)
);

OAI21xp33_ASAP7_75t_L g5951 ( 
.A1(n_5870),
.A2(n_513),
.B(n_514),
.Y(n_5951)
);

OAI22xp33_ASAP7_75t_L g5952 ( 
.A1(n_5843),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_5952)
);

INVx2_ASAP7_75t_L g5953 ( 
.A(n_5851),
.Y(n_5953)
);

AOI22xp33_ASAP7_75t_L g5954 ( 
.A1(n_5871),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_5954)
);

AOI22xp33_ASAP7_75t_L g5955 ( 
.A1(n_5871),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_5955)
);

AOI221xp5_ASAP7_75t_L g5956 ( 
.A1(n_5806),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.C(n_522),
.Y(n_5956)
);

AOI22xp33_ASAP7_75t_L g5957 ( 
.A1(n_5878),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.Y(n_5957)
);

AOI21xp5_ASAP7_75t_L g5958 ( 
.A1(n_5883),
.A2(n_522),
.B(n_523),
.Y(n_5958)
);

AOI22xp33_ASAP7_75t_L g5959 ( 
.A1(n_5878),
.A2(n_525),
.B1(n_523),
.B2(n_524),
.Y(n_5959)
);

OAI221xp5_ASAP7_75t_L g5960 ( 
.A1(n_5873),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.C(n_527),
.Y(n_5960)
);

INVx2_ASAP7_75t_L g5961 ( 
.A(n_5809),
.Y(n_5961)
);

OR2x2_ASAP7_75t_L g5962 ( 
.A(n_5819),
.B(n_525),
.Y(n_5962)
);

INVx4_ASAP7_75t_L g5963 ( 
.A(n_5876),
.Y(n_5963)
);

OAI31xp33_ASAP7_75t_L g5964 ( 
.A1(n_5822),
.A2(n_528),
.A3(n_526),
.B(n_527),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5830),
.Y(n_5965)
);

BUFx6f_ASAP7_75t_L g5966 ( 
.A(n_5860),
.Y(n_5966)
);

AOI221xp5_ASAP7_75t_SL g5967 ( 
.A1(n_5832),
.A2(n_528),
.B1(n_526),
.B2(n_527),
.C(n_529),
.Y(n_5967)
);

HB1xp67_ASAP7_75t_L g5968 ( 
.A(n_5836),
.Y(n_5968)
);

OAI22xp5_ASAP7_75t_L g5969 ( 
.A1(n_5817),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.Y(n_5969)
);

AOI22xp33_ASAP7_75t_L g5970 ( 
.A1(n_5858),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_5970)
);

AOI33xp33_ASAP7_75t_L g5971 ( 
.A1(n_5867),
.A2(n_533),
.A3(n_535),
.B1(n_531),
.B2(n_532),
.B3(n_534),
.Y(n_5971)
);

INVx2_ASAP7_75t_L g5972 ( 
.A(n_5802),
.Y(n_5972)
);

OAI222xp33_ASAP7_75t_L g5973 ( 
.A1(n_5858),
.A2(n_535),
.B1(n_537),
.B2(n_533),
.C1(n_534),
.C2(n_536),
.Y(n_5973)
);

INVx2_ASAP7_75t_L g5974 ( 
.A(n_5802),
.Y(n_5974)
);

INVx1_ASAP7_75t_L g5975 ( 
.A(n_5882),
.Y(n_5975)
);

OAI321xp33_ASAP7_75t_L g5976 ( 
.A1(n_5817),
.A2(n_536),
.A3(n_538),
.B1(n_533),
.B2(n_535),
.C(n_537),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5882),
.Y(n_5977)
);

NAND3xp33_ASAP7_75t_L g5978 ( 
.A(n_5858),
.B(n_536),
.C(n_538),
.Y(n_5978)
);

OAI21xp5_ASAP7_75t_SL g5979 ( 
.A1(n_5858),
.A2(n_538),
.B(n_539),
.Y(n_5979)
);

AOI221xp5_ASAP7_75t_L g5980 ( 
.A1(n_5858),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.C(n_542),
.Y(n_5980)
);

INVx2_ASAP7_75t_L g5981 ( 
.A(n_5802),
.Y(n_5981)
);

AOI211xp5_ASAP7_75t_SL g5982 ( 
.A1(n_5868),
.A2(n_541),
.B(n_539),
.C(n_540),
.Y(n_5982)
);

OA21x2_ASAP7_75t_L g5983 ( 
.A1(n_5804),
.A2(n_541),
.B(n_542),
.Y(n_5983)
);

INVx2_ASAP7_75t_L g5984 ( 
.A(n_5802),
.Y(n_5984)
);

AOI33xp33_ASAP7_75t_L g5985 ( 
.A1(n_5867),
.A2(n_545),
.A3(n_547),
.B1(n_543),
.B2(n_544),
.B3(n_546),
.Y(n_5985)
);

OAI22xp5_ASAP7_75t_L g5986 ( 
.A1(n_5817),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5882),
.Y(n_5987)
);

OAI221xp5_ASAP7_75t_L g5988 ( 
.A1(n_5817),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.C(n_546),
.Y(n_5988)
);

OAI33xp33_ASAP7_75t_L g5989 ( 
.A1(n_5867),
.A2(n_548),
.A3(n_550),
.B1(n_546),
.B2(n_547),
.B3(n_549),
.Y(n_5989)
);

INVxp67_ASAP7_75t_SL g5990 ( 
.A(n_5839),
.Y(n_5990)
);

OR2x2_ASAP7_75t_L g5991 ( 
.A(n_5867),
.B(n_548),
.Y(n_5991)
);

OAI221xp5_ASAP7_75t_L g5992 ( 
.A1(n_5817),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.C(n_551),
.Y(n_5992)
);

AND2x2_ASAP7_75t_L g5993 ( 
.A(n_5797),
.B(n_549),
.Y(n_5993)
);

AND2x2_ASAP7_75t_L g5994 ( 
.A(n_5797),
.B(n_550),
.Y(n_5994)
);

OAI221xp5_ASAP7_75t_L g5995 ( 
.A1(n_5817),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.C(n_554),
.Y(n_5995)
);

NAND3xp33_ASAP7_75t_L g5996 ( 
.A(n_5858),
.B(n_553),
.C(n_554),
.Y(n_5996)
);

AOI22xp5_ASAP7_75t_L g5997 ( 
.A1(n_5858),
.A2(n_557),
.B1(n_553),
.B2(n_556),
.Y(n_5997)
);

AOI221xp5_ASAP7_75t_L g5998 ( 
.A1(n_5858),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.C(n_560),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5882),
.Y(n_5999)
);

AND2x2_ASAP7_75t_L g6000 ( 
.A(n_5797),
.B(n_558),
.Y(n_6000)
);

OAI321xp33_ASAP7_75t_L g6001 ( 
.A1(n_5817),
.A2(n_560),
.A3(n_562),
.B1(n_558),
.B2(n_559),
.C(n_561),
.Y(n_6001)
);

AOI22xp33_ASAP7_75t_L g6002 ( 
.A1(n_5858),
.A2(n_561),
.B1(n_559),
.B2(n_560),
.Y(n_6002)
);

INVx2_ASAP7_75t_L g6003 ( 
.A(n_5802),
.Y(n_6003)
);

INVxp67_ASAP7_75t_SL g6004 ( 
.A(n_5839),
.Y(n_6004)
);

BUFx6f_ASAP7_75t_L g6005 ( 
.A(n_5796),
.Y(n_6005)
);

AOI222xp33_ASAP7_75t_L g6006 ( 
.A1(n_5858),
.A2(n_563),
.B1(n_565),
.B2(n_561),
.C1(n_562),
.C2(n_564),
.Y(n_6006)
);

AOI22xp33_ASAP7_75t_SL g6007 ( 
.A1(n_5858),
.A2(n_564),
.B1(n_562),
.B2(n_563),
.Y(n_6007)
);

OAI221xp5_ASAP7_75t_L g6008 ( 
.A1(n_5817),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.C(n_566),
.Y(n_6008)
);

INVxp67_ASAP7_75t_SL g6009 ( 
.A(n_5839),
.Y(n_6009)
);

AOI22xp33_ASAP7_75t_L g6010 ( 
.A1(n_5858),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.Y(n_6010)
);

AOI22xp33_ASAP7_75t_L g6011 ( 
.A1(n_5858),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_6011)
);

NOR3xp33_ASAP7_75t_SL g6012 ( 
.A(n_5868),
.B(n_567),
.C(n_568),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_5882),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5916),
.Y(n_6014)
);

AND2x2_ASAP7_75t_L g6015 ( 
.A(n_5925),
.B(n_569),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5908),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5913),
.Y(n_6017)
);

BUFx3_ASAP7_75t_L g6018 ( 
.A(n_6005),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_5898),
.Y(n_6019)
);

OR2x2_ASAP7_75t_L g6020 ( 
.A(n_5991),
.B(n_569),
.Y(n_6020)
);

INVx5_ASAP7_75t_L g6021 ( 
.A(n_6005),
.Y(n_6021)
);

INVx2_ASAP7_75t_L g6022 ( 
.A(n_5887),
.Y(n_6022)
);

INVx2_ASAP7_75t_L g6023 ( 
.A(n_5972),
.Y(n_6023)
);

OR2x2_ASAP7_75t_L g6024 ( 
.A(n_5912),
.B(n_570),
.Y(n_6024)
);

INVx3_ASAP7_75t_L g6025 ( 
.A(n_5930),
.Y(n_6025)
);

NAND2xp5_ASAP7_75t_L g6026 ( 
.A(n_6007),
.B(n_570),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5936),
.B(n_5931),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5919),
.Y(n_6028)
);

INVx2_ASAP7_75t_L g6029 ( 
.A(n_5974),
.Y(n_6029)
);

AND2x2_ASAP7_75t_L g6030 ( 
.A(n_5899),
.B(n_571),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5940),
.Y(n_6031)
);

OR2x6_ASAP7_75t_SL g6032 ( 
.A(n_5917),
.B(n_571),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5892),
.Y(n_6033)
);

AND2x2_ASAP7_75t_L g6034 ( 
.A(n_5990),
.B(n_572),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5975),
.Y(n_6035)
);

AND2x2_ASAP7_75t_L g6036 ( 
.A(n_6004),
.B(n_572),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5977),
.Y(n_6037)
);

AND2x2_ASAP7_75t_L g6038 ( 
.A(n_6009),
.B(n_572),
.Y(n_6038)
);

INVx2_ASAP7_75t_L g6039 ( 
.A(n_5981),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5987),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5949),
.B(n_573),
.Y(n_6041)
);

OR2x2_ASAP7_75t_L g6042 ( 
.A(n_5999),
.B(n_573),
.Y(n_6042)
);

INVx2_ASAP7_75t_L g6043 ( 
.A(n_5984),
.Y(n_6043)
);

AND2x4_ASAP7_75t_L g6044 ( 
.A(n_6005),
.B(n_573),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_6013),
.Y(n_6045)
);

INVx2_ASAP7_75t_L g6046 ( 
.A(n_6003),
.Y(n_6046)
);

AND2x2_ASAP7_75t_L g6047 ( 
.A(n_5949),
.B(n_574),
.Y(n_6047)
);

INVx2_ASAP7_75t_L g6048 ( 
.A(n_5893),
.Y(n_6048)
);

NOR2xp33_ASAP7_75t_L g6049 ( 
.A(n_5909),
.B(n_5973),
.Y(n_6049)
);

AND2x2_ASAP7_75t_L g6050 ( 
.A(n_5949),
.B(n_574),
.Y(n_6050)
);

INVx2_ASAP7_75t_L g6051 ( 
.A(n_5953),
.Y(n_6051)
);

AND2x2_ASAP7_75t_L g6052 ( 
.A(n_5938),
.B(n_575),
.Y(n_6052)
);

INVx2_ASAP7_75t_L g6053 ( 
.A(n_5983),
.Y(n_6053)
);

AND2x2_ASAP7_75t_L g6054 ( 
.A(n_5963),
.B(n_575),
.Y(n_6054)
);

INVx2_ASAP7_75t_L g6055 ( 
.A(n_5983),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5894),
.Y(n_6056)
);

INVx5_ASAP7_75t_SL g6057 ( 
.A(n_5966),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_5928),
.Y(n_6058)
);

AND2x2_ASAP7_75t_L g6059 ( 
.A(n_5886),
.B(n_576),
.Y(n_6059)
);

AND2x2_ASAP7_75t_L g6060 ( 
.A(n_5993),
.B(n_576),
.Y(n_6060)
);

INVx2_ASAP7_75t_L g6061 ( 
.A(n_5928),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5968),
.Y(n_6062)
);

INVx1_ASAP7_75t_L g6063 ( 
.A(n_5942),
.Y(n_6063)
);

NAND2xp5_ASAP7_75t_L g6064 ( 
.A(n_6006),
.B(n_576),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5928),
.Y(n_6065)
);

BUFx3_ASAP7_75t_L g6066 ( 
.A(n_5966),
.Y(n_6066)
);

AND2x2_ASAP7_75t_L g6067 ( 
.A(n_5994),
.B(n_577),
.Y(n_6067)
);

AND2x2_ASAP7_75t_L g6068 ( 
.A(n_6000),
.B(n_577),
.Y(n_6068)
);

AND2x2_ASAP7_75t_L g6069 ( 
.A(n_5914),
.B(n_5923),
.Y(n_6069)
);

HB1xp67_ASAP7_75t_L g6070 ( 
.A(n_5896),
.Y(n_6070)
);

INVx2_ASAP7_75t_L g6071 ( 
.A(n_5961),
.Y(n_6071)
);

AND2x2_ASAP7_75t_L g6072 ( 
.A(n_5888),
.B(n_577),
.Y(n_6072)
);

OR2x2_ASAP7_75t_L g6073 ( 
.A(n_5978),
.B(n_578),
.Y(n_6073)
);

NAND2xp5_ASAP7_75t_L g6074 ( 
.A(n_5979),
.B(n_5970),
.Y(n_6074)
);

AND2x2_ASAP7_75t_L g6075 ( 
.A(n_6002),
.B(n_578),
.Y(n_6075)
);

INVx1_ASAP7_75t_L g6076 ( 
.A(n_5902),
.Y(n_6076)
);

NAND2xp5_ASAP7_75t_L g6077 ( 
.A(n_6010),
.B(n_578),
.Y(n_6077)
);

INVx2_ASAP7_75t_L g6078 ( 
.A(n_5947),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5903),
.Y(n_6079)
);

AND2x2_ASAP7_75t_L g6080 ( 
.A(n_6011),
.B(n_579),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5943),
.Y(n_6081)
);

NAND2xp5_ASAP7_75t_L g6082 ( 
.A(n_5980),
.B(n_579),
.Y(n_6082)
);

NAND2xp5_ASAP7_75t_L g6083 ( 
.A(n_5998),
.B(n_580),
.Y(n_6083)
);

AND2x2_ASAP7_75t_L g6084 ( 
.A(n_5997),
.B(n_580),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_5948),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_5906),
.B(n_581),
.Y(n_6086)
);

INVx1_ASAP7_75t_L g6087 ( 
.A(n_5965),
.Y(n_6087)
);

NAND2xp5_ASAP7_75t_L g6088 ( 
.A(n_5934),
.B(n_581),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5962),
.Y(n_6089)
);

HB1xp67_ASAP7_75t_L g6090 ( 
.A(n_5996),
.Y(n_6090)
);

AND2x2_ASAP7_75t_L g6091 ( 
.A(n_5905),
.B(n_581),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_5952),
.Y(n_6092)
);

AND2x4_ASAP7_75t_SL g6093 ( 
.A(n_6012),
.B(n_582),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_5904),
.B(n_582),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_5941),
.Y(n_6095)
);

HB1xp67_ASAP7_75t_L g6096 ( 
.A(n_5929),
.Y(n_6096)
);

INVx1_ASAP7_75t_L g6097 ( 
.A(n_5945),
.Y(n_6097)
);

AND2x2_ASAP7_75t_L g6098 ( 
.A(n_5911),
.B(n_5933),
.Y(n_6098)
);

AND2x2_ASAP7_75t_L g6099 ( 
.A(n_5969),
.B(n_582),
.Y(n_6099)
);

INVx2_ASAP7_75t_L g6100 ( 
.A(n_5946),
.Y(n_6100)
);

OR2x2_ASAP7_75t_L g6101 ( 
.A(n_5986),
.B(n_583),
.Y(n_6101)
);

INVx2_ASAP7_75t_L g6102 ( 
.A(n_6008),
.Y(n_6102)
);

NOR2xp33_ASAP7_75t_L g6103 ( 
.A(n_5910),
.B(n_583),
.Y(n_6103)
);

AND2x4_ASAP7_75t_L g6104 ( 
.A(n_5891),
.B(n_583),
.Y(n_6104)
);

INVx1_ASAP7_75t_L g6105 ( 
.A(n_5901),
.Y(n_6105)
);

NAND2xp5_ASAP7_75t_L g6106 ( 
.A(n_5935),
.B(n_585),
.Y(n_6106)
);

AND2x2_ASAP7_75t_L g6107 ( 
.A(n_5895),
.B(n_585),
.Y(n_6107)
);

INVx2_ASAP7_75t_L g6108 ( 
.A(n_5988),
.Y(n_6108)
);

AND2x2_ASAP7_75t_L g6109 ( 
.A(n_5897),
.B(n_585),
.Y(n_6109)
);

INVx2_ASAP7_75t_L g6110 ( 
.A(n_5992),
.Y(n_6110)
);

AND2x4_ASAP7_75t_L g6111 ( 
.A(n_5926),
.B(n_586),
.Y(n_6111)
);

INVx2_ASAP7_75t_L g6112 ( 
.A(n_5995),
.Y(n_6112)
);

INVx1_ASAP7_75t_L g6113 ( 
.A(n_5960),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_5937),
.Y(n_6114)
);

AND2x2_ASAP7_75t_L g6115 ( 
.A(n_5927),
.B(n_586),
.Y(n_6115)
);

AND2x2_ASAP7_75t_L g6116 ( 
.A(n_5951),
.B(n_586),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5890),
.Y(n_6117)
);

BUFx2_ASAP7_75t_L g6118 ( 
.A(n_5889),
.Y(n_6118)
);

AND2x2_ASAP7_75t_L g6119 ( 
.A(n_5915),
.B(n_587),
.Y(n_6119)
);

OR2x2_ASAP7_75t_L g6120 ( 
.A(n_5964),
.B(n_588),
.Y(n_6120)
);

INVx1_ASAP7_75t_L g6121 ( 
.A(n_5971),
.Y(n_6121)
);

A2O1A1Ixp33_ASAP7_75t_L g6122 ( 
.A1(n_6049),
.A2(n_5900),
.B(n_5982),
.C(n_6001),
.Y(n_6122)
);

INVx4_ASAP7_75t_L g6123 ( 
.A(n_6025),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_6030),
.Y(n_6124)
);

OR2x2_ASAP7_75t_L g6125 ( 
.A(n_6019),
.B(n_5932),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_6034),
.Y(n_6126)
);

AOI22xp5_ASAP7_75t_L g6127 ( 
.A1(n_6105),
.A2(n_5924),
.B1(n_5944),
.B2(n_5920),
.Y(n_6127)
);

AOI22xp33_ASAP7_75t_L g6128 ( 
.A1(n_6066),
.A2(n_5989),
.B1(n_5956),
.B2(n_5958),
.Y(n_6128)
);

AOI22xp5_ASAP7_75t_L g6129 ( 
.A1(n_6103),
.A2(n_5967),
.B1(n_5939),
.B2(n_5955),
.Y(n_6129)
);

AND2x4_ASAP7_75t_SL g6130 ( 
.A(n_6025),
.B(n_5922),
.Y(n_6130)
);

AND2x2_ASAP7_75t_L g6131 ( 
.A(n_6027),
.B(n_5921),
.Y(n_6131)
);

AND2x2_ASAP7_75t_SL g6132 ( 
.A(n_6053),
.B(n_5985),
.Y(n_6132)
);

AOI31xp33_ASAP7_75t_L g6133 ( 
.A1(n_6114),
.A2(n_5954),
.A3(n_5959),
.B(n_5957),
.Y(n_6133)
);

HB1xp67_ASAP7_75t_L g6134 ( 
.A(n_6028),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_6057),
.B(n_5950),
.Y(n_6135)
);

AOI22xp33_ASAP7_75t_L g6136 ( 
.A1(n_6018),
.A2(n_5918),
.B1(n_5976),
.B2(n_5907),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_6036),
.Y(n_6137)
);

NAND2xp5_ASAP7_75t_L g6138 ( 
.A(n_6052),
.B(n_589),
.Y(n_6138)
);

NOR2xp33_ASAP7_75t_L g6139 ( 
.A(n_6021),
.B(n_589),
.Y(n_6139)
);

AND2x2_ASAP7_75t_L g6140 ( 
.A(n_6057),
.B(n_589),
.Y(n_6140)
);

AND2x2_ASAP7_75t_L g6141 ( 
.A(n_6114),
.B(n_590),
.Y(n_6141)
);

NAND2xp5_ASAP7_75t_L g6142 ( 
.A(n_6117),
.B(n_590),
.Y(n_6142)
);

INVx3_ASAP7_75t_L g6143 ( 
.A(n_6021),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_6038),
.Y(n_6144)
);

AO22x1_ASAP7_75t_L g6145 ( 
.A1(n_6055),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.Y(n_6145)
);

AND2x2_ASAP7_75t_L g6146 ( 
.A(n_6069),
.B(n_591),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_6015),
.Y(n_6147)
);

AOI33xp33_ASAP7_75t_L g6148 ( 
.A1(n_6098),
.A2(n_593),
.A3(n_595),
.B1(n_591),
.B2(n_592),
.B3(n_594),
.Y(n_6148)
);

AND2x2_ASAP7_75t_L g6149 ( 
.A(n_6016),
.B(n_593),
.Y(n_6149)
);

AND2x2_ASAP7_75t_L g6150 ( 
.A(n_6016),
.B(n_593),
.Y(n_6150)
);

OR2x2_ASAP7_75t_L g6151 ( 
.A(n_6017),
.B(n_594),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_6065),
.Y(n_6152)
);

INVx1_ASAP7_75t_L g6153 ( 
.A(n_6058),
.Y(n_6153)
);

AND2x2_ASAP7_75t_L g6154 ( 
.A(n_6017),
.B(n_6092),
.Y(n_6154)
);

OAI31xp33_ASAP7_75t_L g6155 ( 
.A1(n_6090),
.A2(n_597),
.A3(n_595),
.B(n_596),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_6061),
.Y(n_6156)
);

NAND3xp33_ASAP7_75t_L g6157 ( 
.A(n_6021),
.B(n_595),
.C(n_596),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_6054),
.Y(n_6158)
);

AND2x6_ASAP7_75t_SL g6159 ( 
.A(n_6064),
.B(n_598),
.Y(n_6159)
);

NAND2xp5_ASAP7_75t_SL g6160 ( 
.A(n_6102),
.B(n_598),
.Y(n_6160)
);

OAI22xp5_ASAP7_75t_L g6161 ( 
.A1(n_6097),
.A2(n_600),
.B1(n_598),
.B2(n_599),
.Y(n_6161)
);

BUFx6f_ASAP7_75t_L g6162 ( 
.A(n_6044),
.Y(n_6162)
);

AND2x2_ASAP7_75t_L g6163 ( 
.A(n_6100),
.B(n_599),
.Y(n_6163)
);

NAND2xp5_ASAP7_75t_L g6164 ( 
.A(n_6117),
.B(n_600),
.Y(n_6164)
);

OR2x2_ASAP7_75t_L g6165 ( 
.A(n_6031),
.B(n_601),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_6041),
.Y(n_6166)
);

INVx3_ASAP7_75t_L g6167 ( 
.A(n_6022),
.Y(n_6167)
);

AOI221xp5_ASAP7_75t_L g6168 ( 
.A1(n_6062),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.C(n_604),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_6047),
.Y(n_6169)
);

OAI21xp5_ASAP7_75t_L g6170 ( 
.A1(n_6096),
.A2(n_602),
.B(n_603),
.Y(n_6170)
);

AND2x2_ASAP7_75t_L g6171 ( 
.A(n_6078),
.B(n_6014),
.Y(n_6171)
);

INVx5_ASAP7_75t_L g6172 ( 
.A(n_6044),
.Y(n_6172)
);

OR2x2_ASAP7_75t_L g6173 ( 
.A(n_6121),
.B(n_602),
.Y(n_6173)
);

AOI22xp33_ASAP7_75t_L g6174 ( 
.A1(n_6118),
.A2(n_6110),
.B1(n_6112),
.B2(n_6108),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_6050),
.Y(n_6175)
);

INVxp67_ASAP7_75t_SL g6176 ( 
.A(n_6020),
.Y(n_6176)
);

NAND5xp2_ASAP7_75t_L g6177 ( 
.A(n_6121),
.B(n_606),
.C(n_603),
.D(n_605),
.E(n_607),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_6023),
.Y(n_6178)
);

AND2x2_ASAP7_75t_L g6179 ( 
.A(n_6095),
.B(n_605),
.Y(n_6179)
);

NAND2xp5_ASAP7_75t_L g6180 ( 
.A(n_6113),
.B(n_605),
.Y(n_6180)
);

INVx1_ASAP7_75t_L g6181 ( 
.A(n_6029),
.Y(n_6181)
);

NOR2xp33_ASAP7_75t_L g6182 ( 
.A(n_6032),
.B(n_606),
.Y(n_6182)
);

AND2x2_ASAP7_75t_L g6183 ( 
.A(n_6063),
.B(n_606),
.Y(n_6183)
);

OR2x2_ASAP7_75t_L g6184 ( 
.A(n_6039),
.B(n_607),
.Y(n_6184)
);

BUFx2_ASAP7_75t_L g6185 ( 
.A(n_6043),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_6046),
.Y(n_6186)
);

AND2x2_ASAP7_75t_L g6187 ( 
.A(n_6089),
.B(n_607),
.Y(n_6187)
);

NAND2xp5_ASAP7_75t_L g6188 ( 
.A(n_6104),
.B(n_608),
.Y(n_6188)
);

OAI31xp33_ASAP7_75t_L g6189 ( 
.A1(n_6093),
.A2(n_610),
.A3(n_608),
.B(n_609),
.Y(n_6189)
);

NAND2xp5_ASAP7_75t_SL g6190 ( 
.A(n_6074),
.B(n_608),
.Y(n_6190)
);

NAND2xp5_ASAP7_75t_L g6191 ( 
.A(n_6104),
.B(n_6119),
.Y(n_6191)
);

AOI221xp5_ASAP7_75t_L g6192 ( 
.A1(n_6056),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.C(n_612),
.Y(n_6192)
);

AND2x2_ASAP7_75t_L g6193 ( 
.A(n_6048),
.B(n_6051),
.Y(n_6193)
);

AOI22xp33_ASAP7_75t_L g6194 ( 
.A1(n_6071),
.A2(n_612),
.B1(n_609),
.B2(n_610),
.Y(n_6194)
);

AND2x2_ASAP7_75t_L g6195 ( 
.A(n_6059),
.B(n_6060),
.Y(n_6195)
);

AND2x2_ASAP7_75t_L g6196 ( 
.A(n_6067),
.B(n_613),
.Y(n_6196)
);

OR2x2_ASAP7_75t_L g6197 ( 
.A(n_6042),
.B(n_613),
.Y(n_6197)
);

AND2x2_ASAP7_75t_L g6198 ( 
.A(n_6068),
.B(n_613),
.Y(n_6198)
);

OAI321xp33_ASAP7_75t_L g6199 ( 
.A1(n_6033),
.A2(n_616),
.A3(n_618),
.B1(n_614),
.B2(n_615),
.C(n_617),
.Y(n_6199)
);

AND2x2_ASAP7_75t_L g6200 ( 
.A(n_6091),
.B(n_614),
.Y(n_6200)
);

AND2x2_ASAP7_75t_L g6201 ( 
.A(n_6035),
.B(n_614),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_6070),
.Y(n_6202)
);

NAND2xp5_ASAP7_75t_L g6203 ( 
.A(n_6107),
.B(n_615),
.Y(n_6203)
);

AND2x2_ASAP7_75t_L g6204 ( 
.A(n_6037),
.B(n_615),
.Y(n_6204)
);

AND2x2_ASAP7_75t_L g6205 ( 
.A(n_6040),
.B(n_616),
.Y(n_6205)
);

INVxp67_ASAP7_75t_SL g6206 ( 
.A(n_6073),
.Y(n_6206)
);

INVx1_ASAP7_75t_L g6207 ( 
.A(n_6120),
.Y(n_6207)
);

INVx3_ASAP7_75t_L g6208 ( 
.A(n_6045),
.Y(n_6208)
);

INVx3_ASAP7_75t_L g6209 ( 
.A(n_6111),
.Y(n_6209)
);

INVx2_ASAP7_75t_SL g6210 ( 
.A(n_6024),
.Y(n_6210)
);

AOI221xp5_ASAP7_75t_L g6211 ( 
.A1(n_6076),
.A2(n_619),
.B1(n_617),
.B2(n_618),
.C(n_620),
.Y(n_6211)
);

AND2x2_ASAP7_75t_L g6212 ( 
.A(n_6111),
.B(n_618),
.Y(n_6212)
);

AND2x2_ASAP7_75t_L g6213 ( 
.A(n_6116),
.B(n_619),
.Y(n_6213)
);

OAI21xp5_ASAP7_75t_SL g6214 ( 
.A1(n_6099),
.A2(n_619),
.B(n_620),
.Y(n_6214)
);

NAND2xp5_ASAP7_75t_L g6215 ( 
.A(n_6072),
.B(n_622),
.Y(n_6215)
);

INVx2_ASAP7_75t_L g6216 ( 
.A(n_6101),
.Y(n_6216)
);

INVx5_ASAP7_75t_L g6217 ( 
.A(n_6084),
.Y(n_6217)
);

INVx1_ASAP7_75t_L g6218 ( 
.A(n_6088),
.Y(n_6218)
);

HB1xp67_ASAP7_75t_L g6219 ( 
.A(n_6076),
.Y(n_6219)
);

AND2x2_ASAP7_75t_L g6220 ( 
.A(n_6109),
.B(n_622),
.Y(n_6220)
);

AOI211xp5_ASAP7_75t_SL g6221 ( 
.A1(n_6082),
.A2(n_6083),
.B(n_6026),
.C(n_6106),
.Y(n_6221)
);

OAI33xp33_ASAP7_75t_L g6222 ( 
.A1(n_6079),
.A2(n_6081),
.A3(n_6087),
.B1(n_6085),
.B2(n_6094),
.B3(n_6077),
.Y(n_6222)
);

AND2x2_ASAP7_75t_L g6223 ( 
.A(n_6075),
.B(n_622),
.Y(n_6223)
);

INVx1_ASAP7_75t_L g6224 ( 
.A(n_6079),
.Y(n_6224)
);

NAND2xp5_ASAP7_75t_L g6225 ( 
.A(n_6080),
.B(n_623),
.Y(n_6225)
);

INVx4_ASAP7_75t_L g6226 ( 
.A(n_6086),
.Y(n_6226)
);

INVx2_ASAP7_75t_L g6227 ( 
.A(n_6081),
.Y(n_6227)
);

INVx2_ASAP7_75t_SL g6228 ( 
.A(n_6115),
.Y(n_6228)
);

INVx1_ASAP7_75t_SL g6229 ( 
.A(n_6085),
.Y(n_6229)
);

AOI21xp5_ASAP7_75t_L g6230 ( 
.A1(n_6087),
.A2(n_623),
.B(n_624),
.Y(n_6230)
);

AOI221xp5_ASAP7_75t_L g6231 ( 
.A1(n_6049),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.C(n_627),
.Y(n_6231)
);

AND2x2_ASAP7_75t_L g6232 ( 
.A(n_6027),
.B(n_624),
.Y(n_6232)
);

INVxp67_ASAP7_75t_SL g6233 ( 
.A(n_6030),
.Y(n_6233)
);

NAND3xp33_ASAP7_75t_SL g6234 ( 
.A(n_6049),
.B(n_625),
.C(n_626),
.Y(n_6234)
);

INVx2_ASAP7_75t_SL g6235 ( 
.A(n_6025),
.Y(n_6235)
);

AND2x2_ASAP7_75t_L g6236 ( 
.A(n_6027),
.B(n_627),
.Y(n_6236)
);

HB1xp67_ASAP7_75t_L g6237 ( 
.A(n_6019),
.Y(n_6237)
);

OAI221xp5_ASAP7_75t_L g6238 ( 
.A1(n_6049),
.A2(n_629),
.B1(n_627),
.B2(n_628),
.C(n_630),
.Y(n_6238)
);

AOI221xp5_ASAP7_75t_L g6239 ( 
.A1(n_6049),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.C(n_631),
.Y(n_6239)
);

NAND3xp33_ASAP7_75t_L g6240 ( 
.A(n_6103),
.B(n_628),
.C(n_631),
.Y(n_6240)
);

INVxp67_ASAP7_75t_SL g6241 ( 
.A(n_6030),
.Y(n_6241)
);

OAI31xp33_ASAP7_75t_L g6242 ( 
.A1(n_6049),
.A2(n_633),
.A3(n_631),
.B(n_632),
.Y(n_6242)
);

INVx2_ASAP7_75t_L g6243 ( 
.A(n_6066),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_6030),
.Y(n_6244)
);

AND2x2_ASAP7_75t_L g6245 ( 
.A(n_6027),
.B(n_632),
.Y(n_6245)
);

NAND2xp5_ASAP7_75t_L g6246 ( 
.A(n_6049),
.B(n_632),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_6030),
.Y(n_6247)
);

INVx1_ASAP7_75t_L g6248 ( 
.A(n_6030),
.Y(n_6248)
);

NAND2xp5_ASAP7_75t_L g6249 ( 
.A(n_6231),
.B(n_633),
.Y(n_6249)
);

INVx2_ASAP7_75t_SL g6250 ( 
.A(n_6243),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_6237),
.Y(n_6251)
);

AND2x2_ASAP7_75t_L g6252 ( 
.A(n_6141),
.B(n_634),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_6140),
.Y(n_6253)
);

HB1xp67_ASAP7_75t_L g6254 ( 
.A(n_6134),
.Y(n_6254)
);

BUFx2_ASAP7_75t_L g6255 ( 
.A(n_6123),
.Y(n_6255)
);

AND2x2_ASAP7_75t_L g6256 ( 
.A(n_6232),
.B(n_634),
.Y(n_6256)
);

NAND2x1_ASAP7_75t_L g6257 ( 
.A(n_6143),
.B(n_634),
.Y(n_6257)
);

AND2x2_ASAP7_75t_L g6258 ( 
.A(n_6236),
.B(n_635),
.Y(n_6258)
);

INVxp67_ASAP7_75t_SL g6259 ( 
.A(n_6139),
.Y(n_6259)
);

AND2x2_ASAP7_75t_L g6260 ( 
.A(n_6245),
.B(n_635),
.Y(n_6260)
);

AND2x2_ASAP7_75t_L g6261 ( 
.A(n_6135),
.B(n_636),
.Y(n_6261)
);

INVx3_ASAP7_75t_L g6262 ( 
.A(n_6167),
.Y(n_6262)
);

AND2x2_ASAP7_75t_L g6263 ( 
.A(n_6235),
.B(n_636),
.Y(n_6263)
);

INVxp67_ASAP7_75t_SL g6264 ( 
.A(n_6188),
.Y(n_6264)
);

NAND2xp5_ASAP7_75t_L g6265 ( 
.A(n_6239),
.B(n_637),
.Y(n_6265)
);

NAND2xp5_ASAP7_75t_L g6266 ( 
.A(n_6242),
.B(n_637),
.Y(n_6266)
);

NAND2xp5_ASAP7_75t_L g6267 ( 
.A(n_6148),
.B(n_638),
.Y(n_6267)
);

INVx2_ASAP7_75t_SL g6268 ( 
.A(n_6172),
.Y(n_6268)
);

INVx1_ASAP7_75t_L g6269 ( 
.A(n_6212),
.Y(n_6269)
);

OR2x2_ASAP7_75t_L g6270 ( 
.A(n_6173),
.B(n_638),
.Y(n_6270)
);

INVx2_ASAP7_75t_L g6271 ( 
.A(n_6193),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_6185),
.Y(n_6272)
);

NAND2xp5_ASAP7_75t_L g6273 ( 
.A(n_6145),
.B(n_639),
.Y(n_6273)
);

NAND2xp5_ASAP7_75t_L g6274 ( 
.A(n_6122),
.B(n_639),
.Y(n_6274)
);

AND2x2_ASAP7_75t_L g6275 ( 
.A(n_6131),
.B(n_640),
.Y(n_6275)
);

INVx2_ASAP7_75t_L g6276 ( 
.A(n_6162),
.Y(n_6276)
);

OR2x2_ASAP7_75t_L g6277 ( 
.A(n_6191),
.B(n_640),
.Y(n_6277)
);

AND2x2_ASAP7_75t_L g6278 ( 
.A(n_6163),
.B(n_640),
.Y(n_6278)
);

NAND2xp5_ASAP7_75t_SL g6279 ( 
.A(n_6172),
.B(n_641),
.Y(n_6279)
);

INVx1_ASAP7_75t_L g6280 ( 
.A(n_6220),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_6200),
.Y(n_6281)
);

INVx2_ASAP7_75t_L g6282 ( 
.A(n_6162),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_6178),
.Y(n_6283)
);

AND2x2_ASAP7_75t_L g6284 ( 
.A(n_6195),
.B(n_641),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_6181),
.Y(n_6285)
);

INVx2_ASAP7_75t_L g6286 ( 
.A(n_6186),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_6213),
.Y(n_6287)
);

AND2x2_ASAP7_75t_L g6288 ( 
.A(n_6207),
.B(n_641),
.Y(n_6288)
);

AND2x2_ASAP7_75t_L g6289 ( 
.A(n_6154),
.B(n_642),
.Y(n_6289)
);

NAND2xp5_ASAP7_75t_L g6290 ( 
.A(n_6132),
.B(n_642),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_6157),
.Y(n_6291)
);

INVx2_ASAP7_75t_L g6292 ( 
.A(n_6172),
.Y(n_6292)
);

INVx1_ASAP7_75t_L g6293 ( 
.A(n_6153),
.Y(n_6293)
);

INVx2_ASAP7_75t_L g6294 ( 
.A(n_6209),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_6183),
.B(n_642),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_6156),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_6146),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_6197),
.Y(n_6298)
);

OR2x2_ASAP7_75t_L g6299 ( 
.A(n_6246),
.B(n_643),
.Y(n_6299)
);

NAND2x1_ASAP7_75t_L g6300 ( 
.A(n_6208),
.B(n_644),
.Y(n_6300)
);

INVx2_ASAP7_75t_L g6301 ( 
.A(n_6184),
.Y(n_6301)
);

AND2x2_ASAP7_75t_L g6302 ( 
.A(n_6179),
.B(n_644),
.Y(n_6302)
);

INVx1_ASAP7_75t_L g6303 ( 
.A(n_6223),
.Y(n_6303)
);

INVxp33_ASAP7_75t_L g6304 ( 
.A(n_6182),
.Y(n_6304)
);

AND2x2_ASAP7_75t_L g6305 ( 
.A(n_6149),
.B(n_6150),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_6165),
.Y(n_6306)
);

NAND2xp5_ASAP7_75t_SL g6307 ( 
.A(n_6217),
.B(n_645),
.Y(n_6307)
);

OR2x2_ASAP7_75t_L g6308 ( 
.A(n_6180),
.B(n_645),
.Y(n_6308)
);

INVx2_ASAP7_75t_L g6309 ( 
.A(n_6171),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_6196),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_6198),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_6187),
.Y(n_6312)
);

NAND2xp5_ASAP7_75t_L g6313 ( 
.A(n_6136),
.B(n_645),
.Y(n_6313)
);

AND2x4_ASAP7_75t_L g6314 ( 
.A(n_6130),
.B(n_646),
.Y(n_6314)
);

NAND2xp5_ASAP7_75t_L g6315 ( 
.A(n_6174),
.B(n_646),
.Y(n_6315)
);

INVx2_ASAP7_75t_L g6316 ( 
.A(n_6210),
.Y(n_6316)
);

AND2x2_ASAP7_75t_L g6317 ( 
.A(n_6233),
.B(n_647),
.Y(n_6317)
);

NAND2xp5_ASAP7_75t_L g6318 ( 
.A(n_6128),
.B(n_647),
.Y(n_6318)
);

INVx1_ASAP7_75t_L g6319 ( 
.A(n_6219),
.Y(n_6319)
);

INVx2_ASAP7_75t_L g6320 ( 
.A(n_6125),
.Y(n_6320)
);

NAND2xp5_ASAP7_75t_L g6321 ( 
.A(n_6241),
.B(n_648),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_6201),
.Y(n_6322)
);

INVx2_ASAP7_75t_L g6323 ( 
.A(n_6202),
.Y(n_6323)
);

INVx2_ASAP7_75t_L g6324 ( 
.A(n_6152),
.Y(n_6324)
);

OR2x2_ASAP7_75t_L g6325 ( 
.A(n_6142),
.B(n_648),
.Y(n_6325)
);

OR2x2_ASAP7_75t_L g6326 ( 
.A(n_6164),
.B(n_648),
.Y(n_6326)
);

INVx2_ASAP7_75t_L g6327 ( 
.A(n_6216),
.Y(n_6327)
);

NAND2xp5_ASAP7_75t_L g6328 ( 
.A(n_6221),
.B(n_649),
.Y(n_6328)
);

NAND2xp5_ASAP7_75t_L g6329 ( 
.A(n_6127),
.B(n_649),
.Y(n_6329)
);

INVx2_ASAP7_75t_L g6330 ( 
.A(n_6227),
.Y(n_6330)
);

INVx1_ASAP7_75t_L g6331 ( 
.A(n_6204),
.Y(n_6331)
);

INVx1_ASAP7_75t_L g6332 ( 
.A(n_6205),
.Y(n_6332)
);

INVx1_ASAP7_75t_SL g6333 ( 
.A(n_6151),
.Y(n_6333)
);

OR2x2_ASAP7_75t_L g6334 ( 
.A(n_6126),
.B(n_649),
.Y(n_6334)
);

INVx1_ASAP7_75t_L g6335 ( 
.A(n_6166),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_6169),
.Y(n_6336)
);

AND2x2_ASAP7_75t_L g6337 ( 
.A(n_6217),
.B(n_6137),
.Y(n_6337)
);

NAND2xp5_ASAP7_75t_L g6338 ( 
.A(n_6228),
.B(n_650),
.Y(n_6338)
);

NAND2xp5_ASAP7_75t_L g6339 ( 
.A(n_6226),
.B(n_650),
.Y(n_6339)
);

INVxp67_ASAP7_75t_SL g6340 ( 
.A(n_6215),
.Y(n_6340)
);

OR2x2_ASAP7_75t_L g6341 ( 
.A(n_6144),
.B(n_6161),
.Y(n_6341)
);

AND2x2_ASAP7_75t_L g6342 ( 
.A(n_6217),
.B(n_651),
.Y(n_6342)
);

NOR2x1_ASAP7_75t_L g6343 ( 
.A(n_6234),
.B(n_6238),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_6175),
.Y(n_6344)
);

OR2x2_ASAP7_75t_L g6345 ( 
.A(n_6158),
.B(n_651),
.Y(n_6345)
);

AND2x2_ASAP7_75t_L g6346 ( 
.A(n_6176),
.B(n_651),
.Y(n_6346)
);

INVxp67_ASAP7_75t_L g6347 ( 
.A(n_6177),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_6225),
.Y(n_6348)
);

OR2x2_ASAP7_75t_L g6349 ( 
.A(n_6124),
.B(n_652),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_6138),
.Y(n_6350)
);

INVx1_ASAP7_75t_L g6351 ( 
.A(n_6147),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_6206),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_6244),
.Y(n_6353)
);

AND2x2_ASAP7_75t_L g6354 ( 
.A(n_6247),
.B(n_652),
.Y(n_6354)
);

NOR3xp33_ASAP7_75t_L g6355 ( 
.A(n_6199),
.B(n_653),
.C(n_654),
.Y(n_6355)
);

AND2x4_ASAP7_75t_L g6356 ( 
.A(n_6170),
.B(n_653),
.Y(n_6356)
);

NAND2xp5_ASAP7_75t_L g6357 ( 
.A(n_6129),
.B(n_653),
.Y(n_6357)
);

AND2x2_ASAP7_75t_L g6358 ( 
.A(n_6248),
.B(n_6218),
.Y(n_6358)
);

NAND2xp5_ASAP7_75t_L g6359 ( 
.A(n_6214),
.B(n_6155),
.Y(n_6359)
);

AND2x2_ASAP7_75t_L g6360 ( 
.A(n_6250),
.B(n_6160),
.Y(n_6360)
);

INVx2_ASAP7_75t_L g6361 ( 
.A(n_6255),
.Y(n_6361)
);

NOR2xp33_ASAP7_75t_R g6362 ( 
.A(n_6268),
.B(n_6159),
.Y(n_6362)
);

OR2x2_ASAP7_75t_L g6363 ( 
.A(n_6313),
.B(n_6190),
.Y(n_6363)
);

AND2x2_ASAP7_75t_L g6364 ( 
.A(n_6289),
.B(n_6203),
.Y(n_6364)
);

BUFx2_ASAP7_75t_L g6365 ( 
.A(n_6314),
.Y(n_6365)
);

INVxp67_ASAP7_75t_L g6366 ( 
.A(n_6342),
.Y(n_6366)
);

HB1xp67_ASAP7_75t_L g6367 ( 
.A(n_6263),
.Y(n_6367)
);

INVx2_ASAP7_75t_L g6368 ( 
.A(n_6262),
.Y(n_6368)
);

AND2x2_ASAP7_75t_L g6369 ( 
.A(n_6284),
.B(n_6189),
.Y(n_6369)
);

NAND2xp5_ASAP7_75t_L g6370 ( 
.A(n_6347),
.B(n_6262),
.Y(n_6370)
);

OR2x2_ASAP7_75t_L g6371 ( 
.A(n_6273),
.B(n_6133),
.Y(n_6371)
);

INVx1_ASAP7_75t_SL g6372 ( 
.A(n_6314),
.Y(n_6372)
);

OR2x2_ASAP7_75t_L g6373 ( 
.A(n_6274),
.B(n_6229),
.Y(n_6373)
);

OR2x2_ASAP7_75t_L g6374 ( 
.A(n_6294),
.B(n_6240),
.Y(n_6374)
);

INVx2_ASAP7_75t_SL g6375 ( 
.A(n_6276),
.Y(n_6375)
);

INVxp67_ASAP7_75t_SL g6376 ( 
.A(n_6257),
.Y(n_6376)
);

AND2x2_ASAP7_75t_L g6377 ( 
.A(n_6271),
.B(n_6194),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_6257),
.Y(n_6378)
);

AND2x4_ASAP7_75t_L g6379 ( 
.A(n_6282),
.B(n_6224),
.Y(n_6379)
);

NAND3xp33_ASAP7_75t_SL g6380 ( 
.A(n_6355),
.B(n_6168),
.C(n_6192),
.Y(n_6380)
);

INVx2_ASAP7_75t_SL g6381 ( 
.A(n_6292),
.Y(n_6381)
);

OR2x2_ASAP7_75t_L g6382 ( 
.A(n_6270),
.B(n_6251),
.Y(n_6382)
);

INVx1_ASAP7_75t_SL g6383 ( 
.A(n_6337),
.Y(n_6383)
);

AND2x2_ASAP7_75t_L g6384 ( 
.A(n_6288),
.B(n_6230),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_6278),
.Y(n_6385)
);

OR2x2_ASAP7_75t_L g6386 ( 
.A(n_6328),
.B(n_6315),
.Y(n_6386)
);

AND2x4_ASAP7_75t_SL g6387 ( 
.A(n_6316),
.B(n_6222),
.Y(n_6387)
);

NOR3xp33_ASAP7_75t_SL g6388 ( 
.A(n_6352),
.B(n_6211),
.C(n_655),
.Y(n_6388)
);

AND2x4_ASAP7_75t_L g6389 ( 
.A(n_6272),
.B(n_655),
.Y(n_6389)
);

AND2x2_ASAP7_75t_L g6390 ( 
.A(n_6305),
.B(n_655),
.Y(n_6390)
);

BUFx3_ASAP7_75t_L g6391 ( 
.A(n_6286),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6254),
.Y(n_6392)
);

AND2x2_ASAP7_75t_L g6393 ( 
.A(n_6317),
.B(n_656),
.Y(n_6393)
);

NAND2xp5_ASAP7_75t_L g6394 ( 
.A(n_6261),
.B(n_656),
.Y(n_6394)
);

NAND2xp5_ASAP7_75t_L g6395 ( 
.A(n_6346),
.B(n_656),
.Y(n_6395)
);

NOR2xp33_ASAP7_75t_L g6396 ( 
.A(n_6279),
.B(n_6307),
.Y(n_6396)
);

NAND2x1_ASAP7_75t_SL g6397 ( 
.A(n_6354),
.B(n_657),
.Y(n_6397)
);

NOR2xp33_ASAP7_75t_L g6398 ( 
.A(n_6300),
.B(n_657),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_6252),
.Y(n_6399)
);

NAND2xp5_ASAP7_75t_L g6400 ( 
.A(n_6275),
.B(n_657),
.Y(n_6400)
);

BUFx2_ASAP7_75t_L g6401 ( 
.A(n_6309),
.Y(n_6401)
);

INVx2_ASAP7_75t_L g6402 ( 
.A(n_6327),
.Y(n_6402)
);

OR2x2_ASAP7_75t_L g6403 ( 
.A(n_6321),
.B(n_658),
.Y(n_6403)
);

OR2x2_ASAP7_75t_L g6404 ( 
.A(n_6266),
.B(n_658),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_6339),
.Y(n_6405)
);

NAND2xp33_ASAP7_75t_SL g6406 ( 
.A(n_6300),
.B(n_659),
.Y(n_6406)
);

OR2x2_ASAP7_75t_L g6407 ( 
.A(n_6357),
.B(n_659),
.Y(n_6407)
);

OR2x2_ASAP7_75t_L g6408 ( 
.A(n_6318),
.B(n_659),
.Y(n_6408)
);

NAND2xp5_ASAP7_75t_L g6409 ( 
.A(n_6356),
.B(n_660),
.Y(n_6409)
);

OR2x2_ASAP7_75t_L g6410 ( 
.A(n_6277),
.B(n_660),
.Y(n_6410)
);

NOR3xp33_ASAP7_75t_SL g6411 ( 
.A(n_6329),
.B(n_660),
.C(n_661),
.Y(n_6411)
);

HB1xp67_ASAP7_75t_L g6412 ( 
.A(n_6320),
.Y(n_6412)
);

AND2x4_ASAP7_75t_L g6413 ( 
.A(n_6323),
.B(n_661),
.Y(n_6413)
);

AND2x2_ASAP7_75t_L g6414 ( 
.A(n_6253),
.B(n_661),
.Y(n_6414)
);

NOR2xp33_ASAP7_75t_SL g6415 ( 
.A(n_6256),
.B(n_662),
.Y(n_6415)
);

NAND2xp5_ASAP7_75t_L g6416 ( 
.A(n_6356),
.B(n_662),
.Y(n_6416)
);

AND2x2_ASAP7_75t_L g6417 ( 
.A(n_6343),
.B(n_663),
.Y(n_6417)
);

OR2x2_ASAP7_75t_L g6418 ( 
.A(n_6290),
.B(n_664),
.Y(n_6418)
);

AND2x2_ASAP7_75t_L g6419 ( 
.A(n_6258),
.B(n_664),
.Y(n_6419)
);

AOI221xp5_ASAP7_75t_L g6420 ( 
.A1(n_6291),
.A2(n_667),
.B1(n_665),
.B2(n_666),
.C(n_668),
.Y(n_6420)
);

INVx2_ASAP7_75t_SL g6421 ( 
.A(n_6301),
.Y(n_6421)
);

NAND2xp5_ASAP7_75t_L g6422 ( 
.A(n_6302),
.B(n_665),
.Y(n_6422)
);

AND2x2_ASAP7_75t_L g6423 ( 
.A(n_6260),
.B(n_6297),
.Y(n_6423)
);

INVx1_ASAP7_75t_SL g6424 ( 
.A(n_6295),
.Y(n_6424)
);

AND2x2_ASAP7_75t_L g6425 ( 
.A(n_6280),
.B(n_665),
.Y(n_6425)
);

AND2x2_ASAP7_75t_L g6426 ( 
.A(n_6281),
.B(n_6303),
.Y(n_6426)
);

AND2x2_ASAP7_75t_L g6427 ( 
.A(n_6310),
.B(n_666),
.Y(n_6427)
);

OR2x2_ASAP7_75t_L g6428 ( 
.A(n_6299),
.B(n_666),
.Y(n_6428)
);

NAND2xp5_ASAP7_75t_L g6429 ( 
.A(n_6259),
.B(n_667),
.Y(n_6429)
);

OR2x2_ASAP7_75t_L g6430 ( 
.A(n_6345),
.B(n_667),
.Y(n_6430)
);

INVx2_ASAP7_75t_L g6431 ( 
.A(n_6330),
.Y(n_6431)
);

INVx2_ASAP7_75t_L g6432 ( 
.A(n_6283),
.Y(n_6432)
);

INVx3_ASAP7_75t_L g6433 ( 
.A(n_6285),
.Y(n_6433)
);

AND2x2_ASAP7_75t_L g6434 ( 
.A(n_6311),
.B(n_668),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_6338),
.Y(n_6435)
);

NAND2xp5_ASAP7_75t_L g6436 ( 
.A(n_6333),
.B(n_668),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_6308),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_6312),
.B(n_669),
.Y(n_6438)
);

NOR3xp33_ASAP7_75t_L g6439 ( 
.A(n_6249),
.B(n_669),
.C(n_670),
.Y(n_6439)
);

NAND2xp5_ASAP7_75t_L g6440 ( 
.A(n_6287),
.B(n_670),
.Y(n_6440)
);

AND2x2_ASAP7_75t_L g6441 ( 
.A(n_6358),
.B(n_670),
.Y(n_6441)
);

AND2x2_ASAP7_75t_L g6442 ( 
.A(n_6322),
.B(n_671),
.Y(n_6442)
);

NAND3xp33_ASAP7_75t_SL g6443 ( 
.A(n_6304),
.B(n_671),
.C(n_672),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_6325),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_6326),
.Y(n_6445)
);

AND2x2_ASAP7_75t_L g6446 ( 
.A(n_6331),
.B(n_672),
.Y(n_6446)
);

HB1xp67_ASAP7_75t_L g6447 ( 
.A(n_6293),
.Y(n_6447)
);

NAND2xp5_ASAP7_75t_L g6448 ( 
.A(n_6332),
.B(n_673),
.Y(n_6448)
);

NAND4xp25_ASAP7_75t_L g6449 ( 
.A(n_6359),
.B(n_675),
.C(n_673),
.D(n_674),
.Y(n_6449)
);

AND2x2_ASAP7_75t_L g6450 ( 
.A(n_6269),
.B(n_674),
.Y(n_6450)
);

NAND2xp5_ASAP7_75t_L g6451 ( 
.A(n_6340),
.B(n_675),
.Y(n_6451)
);

OAI31xp33_ASAP7_75t_L g6452 ( 
.A1(n_6319),
.A2(n_677),
.A3(n_675),
.B(n_676),
.Y(n_6452)
);

AOI222xp33_ASAP7_75t_L g6453 ( 
.A1(n_6296),
.A2(n_678),
.B1(n_680),
.B2(n_676),
.C1(n_677),
.C2(n_679),
.Y(n_6453)
);

INVx3_ASAP7_75t_L g6454 ( 
.A(n_6324),
.Y(n_6454)
);

AND2x2_ASAP7_75t_L g6455 ( 
.A(n_6298),
.B(n_676),
.Y(n_6455)
);

NAND2xp5_ASAP7_75t_SL g6456 ( 
.A(n_6341),
.B(n_677),
.Y(n_6456)
);

AND2x4_ASAP7_75t_L g6457 ( 
.A(n_6351),
.B(n_6353),
.Y(n_6457)
);

OAI33xp33_ASAP7_75t_L g6458 ( 
.A1(n_6335),
.A2(n_680),
.A3(n_682),
.B1(n_678),
.B2(n_679),
.B3(n_681),
.Y(n_6458)
);

AND2x2_ASAP7_75t_L g6459 ( 
.A(n_6306),
.B(n_679),
.Y(n_6459)
);

INVx3_ASAP7_75t_L g6460 ( 
.A(n_6349),
.Y(n_6460)
);

INVx2_ASAP7_75t_L g6461 ( 
.A(n_6334),
.Y(n_6461)
);

HB1xp67_ASAP7_75t_L g6462 ( 
.A(n_6336),
.Y(n_6462)
);

NAND2xp5_ASAP7_75t_L g6463 ( 
.A(n_6264),
.B(n_680),
.Y(n_6463)
);

INVx2_ASAP7_75t_SL g6464 ( 
.A(n_6344),
.Y(n_6464)
);

OR2x2_ASAP7_75t_L g6465 ( 
.A(n_6267),
.B(n_6265),
.Y(n_6465)
);

OR2x2_ASAP7_75t_L g6466 ( 
.A(n_6348),
.B(n_681),
.Y(n_6466)
);

AND2x2_ASAP7_75t_L g6467 ( 
.A(n_6350),
.B(n_681),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_6263),
.Y(n_6468)
);

AOI211x1_ASAP7_75t_SL g6469 ( 
.A1(n_6320),
.A2(n_684),
.B(n_682),
.C(n_683),
.Y(n_6469)
);

AOI21xp5_ASAP7_75t_L g6470 ( 
.A1(n_6279),
.A2(n_683),
.B(n_684),
.Y(n_6470)
);

CKINVDCx16_ASAP7_75t_R g6471 ( 
.A(n_6250),
.Y(n_6471)
);

NAND2xp5_ASAP7_75t_L g6472 ( 
.A(n_6250),
.B(n_683),
.Y(n_6472)
);

INVx1_ASAP7_75t_L g6473 ( 
.A(n_6263),
.Y(n_6473)
);

AND2x2_ASAP7_75t_L g6474 ( 
.A(n_6471),
.B(n_684),
.Y(n_6474)
);

AND2x2_ASAP7_75t_L g6475 ( 
.A(n_6383),
.B(n_685),
.Y(n_6475)
);

HB1xp67_ASAP7_75t_L g6476 ( 
.A(n_6412),
.Y(n_6476)
);

INVx3_ASAP7_75t_L g6477 ( 
.A(n_6379),
.Y(n_6477)
);

AND2x4_ASAP7_75t_L g6478 ( 
.A(n_6381),
.B(n_685),
.Y(n_6478)
);

NAND2xp5_ASAP7_75t_L g6479 ( 
.A(n_6376),
.B(n_685),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_6361),
.Y(n_6480)
);

AND2x2_ASAP7_75t_L g6481 ( 
.A(n_6441),
.B(n_6390),
.Y(n_6481)
);

AND2x2_ASAP7_75t_L g6482 ( 
.A(n_6393),
.B(n_686),
.Y(n_6482)
);

NAND2xp5_ASAP7_75t_L g6483 ( 
.A(n_6375),
.B(n_686),
.Y(n_6483)
);

NAND2xp5_ASAP7_75t_L g6484 ( 
.A(n_6372),
.B(n_686),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_6365),
.Y(n_6485)
);

INVx1_ASAP7_75t_L g6486 ( 
.A(n_6472),
.Y(n_6486)
);

AND2x2_ASAP7_75t_L g6487 ( 
.A(n_6417),
.B(n_6369),
.Y(n_6487)
);

INVx1_ASAP7_75t_L g6488 ( 
.A(n_6409),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_6391),
.Y(n_6489)
);

INVx1_ASAP7_75t_SL g6490 ( 
.A(n_6362),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_6416),
.Y(n_6491)
);

AND2x2_ASAP7_75t_L g6492 ( 
.A(n_6360),
.B(n_687),
.Y(n_6492)
);

INVx2_ASAP7_75t_L g6493 ( 
.A(n_6402),
.Y(n_6493)
);

OR2x2_ASAP7_75t_L g6494 ( 
.A(n_6368),
.B(n_687),
.Y(n_6494)
);

AND2x2_ASAP7_75t_L g6495 ( 
.A(n_6455),
.B(n_687),
.Y(n_6495)
);

INVx1_ASAP7_75t_L g6496 ( 
.A(n_6413),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_6413),
.Y(n_6497)
);

NAND2xp5_ASAP7_75t_L g6498 ( 
.A(n_6387),
.B(n_688),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_6389),
.Y(n_6499)
);

OR2x6_ASAP7_75t_L g6500 ( 
.A(n_6370),
.B(n_6431),
.Y(n_6500)
);

NOR2xp33_ASAP7_75t_L g6501 ( 
.A(n_6378),
.B(n_689),
.Y(n_6501)
);

NAND2xp5_ASAP7_75t_L g6502 ( 
.A(n_6469),
.B(n_690),
.Y(n_6502)
);

AND2x2_ASAP7_75t_L g6503 ( 
.A(n_6414),
.B(n_690),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6389),
.Y(n_6504)
);

INVx1_ASAP7_75t_L g6505 ( 
.A(n_6401),
.Y(n_6505)
);

NAND2xp5_ASAP7_75t_L g6506 ( 
.A(n_6419),
.B(n_690),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_6379),
.Y(n_6507)
);

INVxp67_ASAP7_75t_L g6508 ( 
.A(n_6415),
.Y(n_6508)
);

O2A1O1Ixp33_ASAP7_75t_L g6509 ( 
.A1(n_6443),
.A2(n_693),
.B(n_691),
.C(n_692),
.Y(n_6509)
);

AND2x2_ASAP7_75t_L g6510 ( 
.A(n_6425),
.B(n_691),
.Y(n_6510)
);

AND2x4_ASAP7_75t_L g6511 ( 
.A(n_6421),
.B(n_6454),
.Y(n_6511)
);

NAND2xp5_ASAP7_75t_L g6512 ( 
.A(n_6398),
.B(n_691),
.Y(n_6512)
);

AND2x2_ASAP7_75t_L g6513 ( 
.A(n_6427),
.B(n_692),
.Y(n_6513)
);

AND2x2_ASAP7_75t_L g6514 ( 
.A(n_6434),
.B(n_692),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_6367),
.Y(n_6515)
);

AOI221xp5_ASAP7_75t_L g6516 ( 
.A1(n_6380),
.A2(n_695),
.B1(n_693),
.B2(n_694),
.C(n_696),
.Y(n_6516)
);

NAND2xp5_ASAP7_75t_L g6517 ( 
.A(n_6453),
.B(n_694),
.Y(n_6517)
);

NAND2xp5_ASAP7_75t_L g6518 ( 
.A(n_6384),
.B(n_695),
.Y(n_6518)
);

INVx1_ASAP7_75t_L g6519 ( 
.A(n_6374),
.Y(n_6519)
);

AND2x2_ASAP7_75t_L g6520 ( 
.A(n_6459),
.B(n_696),
.Y(n_6520)
);

INVx1_ASAP7_75t_L g6521 ( 
.A(n_6429),
.Y(n_6521)
);

NAND2xp5_ASAP7_75t_L g6522 ( 
.A(n_6364),
.B(n_697),
.Y(n_6522)
);

INVx1_ASAP7_75t_L g6523 ( 
.A(n_6404),
.Y(n_6523)
);

NAND3xp33_ASAP7_75t_L g6524 ( 
.A(n_6452),
.B(n_697),
.C(n_698),
.Y(n_6524)
);

INVx2_ASAP7_75t_L g6525 ( 
.A(n_6392),
.Y(n_6525)
);

AND2x2_ASAP7_75t_L g6526 ( 
.A(n_6450),
.B(n_698),
.Y(n_6526)
);

AND2x2_ASAP7_75t_L g6527 ( 
.A(n_6438),
.B(n_699),
.Y(n_6527)
);

INVx2_ASAP7_75t_L g6528 ( 
.A(n_6382),
.Y(n_6528)
);

NAND2xp5_ASAP7_75t_L g6529 ( 
.A(n_6470),
.B(n_699),
.Y(n_6529)
);

INVx1_ASAP7_75t_L g6530 ( 
.A(n_6422),
.Y(n_6530)
);

AOI211xp5_ASAP7_75t_L g6531 ( 
.A1(n_6396),
.A2(n_6456),
.B(n_6371),
.C(n_6366),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_6428),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_6410),
.Y(n_6533)
);

NAND2x1p5_ASAP7_75t_L g6534 ( 
.A(n_6407),
.B(n_700),
.Y(n_6534)
);

OR2x2_ASAP7_75t_L g6535 ( 
.A(n_6449),
.B(n_700),
.Y(n_6535)
);

OR2x2_ASAP7_75t_L g6536 ( 
.A(n_6430),
.B(n_700),
.Y(n_6536)
);

INVxp67_ASAP7_75t_L g6537 ( 
.A(n_6406),
.Y(n_6537)
);

AND2x4_ASAP7_75t_SL g6538 ( 
.A(n_6423),
.B(n_701),
.Y(n_6538)
);

AND2x2_ASAP7_75t_L g6539 ( 
.A(n_6442),
.B(n_701),
.Y(n_6539)
);

OAI22xp5_ASAP7_75t_L g6540 ( 
.A1(n_6408),
.A2(n_703),
.B1(n_701),
.B2(n_702),
.Y(n_6540)
);

OR2x2_ASAP7_75t_L g6541 ( 
.A(n_6424),
.B(n_702),
.Y(n_6541)
);

AND2x2_ASAP7_75t_L g6542 ( 
.A(n_6446),
.B(n_702),
.Y(n_6542)
);

INVx1_ASAP7_75t_L g6543 ( 
.A(n_6377),
.Y(n_6543)
);

HB1xp67_ASAP7_75t_L g6544 ( 
.A(n_6447),
.Y(n_6544)
);

BUFx2_ASAP7_75t_SL g6545 ( 
.A(n_6432),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6397),
.B(n_6420),
.Y(n_6546)
);

INVx1_ASAP7_75t_L g6547 ( 
.A(n_6436),
.Y(n_6547)
);

NAND2xp5_ASAP7_75t_L g6548 ( 
.A(n_6467),
.B(n_703),
.Y(n_6548)
);

HB1xp67_ASAP7_75t_L g6549 ( 
.A(n_6462),
.Y(n_6549)
);

INVx1_ASAP7_75t_SL g6550 ( 
.A(n_6490),
.Y(n_6550)
);

AND2x2_ASAP7_75t_L g6551 ( 
.A(n_6474),
.B(n_6411),
.Y(n_6551)
);

INVx1_ASAP7_75t_L g6552 ( 
.A(n_6478),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_6478),
.Y(n_6553)
);

NAND2xp33_ASAP7_75t_SL g6554 ( 
.A(n_6498),
.B(n_6388),
.Y(n_6554)
);

AND2x2_ASAP7_75t_L g6555 ( 
.A(n_6475),
.B(n_6385),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_6476),
.Y(n_6556)
);

AND2x4_ASAP7_75t_L g6557 ( 
.A(n_6507),
.B(n_6457),
.Y(n_6557)
);

AND2x2_ASAP7_75t_L g6558 ( 
.A(n_6503),
.B(n_6399),
.Y(n_6558)
);

OR2x2_ASAP7_75t_L g6559 ( 
.A(n_6489),
.B(n_6403),
.Y(n_6559)
);

OR2x2_ASAP7_75t_L g6560 ( 
.A(n_6477),
.B(n_6463),
.Y(n_6560)
);

AND2x2_ASAP7_75t_L g6561 ( 
.A(n_6510),
.B(n_6426),
.Y(n_6561)
);

AOI211xp5_ASAP7_75t_SL g6562 ( 
.A1(n_6537),
.A2(n_6451),
.B(n_6439),
.C(n_6405),
.Y(n_6562)
);

NAND2xp5_ASAP7_75t_L g6563 ( 
.A(n_6511),
.B(n_6468),
.Y(n_6563)
);

HB1xp67_ASAP7_75t_L g6564 ( 
.A(n_6511),
.Y(n_6564)
);

NOR2xp33_ASAP7_75t_L g6565 ( 
.A(n_6480),
.B(n_6395),
.Y(n_6565)
);

AND2x2_ASAP7_75t_L g6566 ( 
.A(n_6513),
.B(n_6473),
.Y(n_6566)
);

NAND2xp5_ASAP7_75t_L g6567 ( 
.A(n_6493),
.B(n_6464),
.Y(n_6567)
);

OR2x2_ASAP7_75t_L g6568 ( 
.A(n_6479),
.B(n_6394),
.Y(n_6568)
);

INVx1_ASAP7_75t_SL g6569 ( 
.A(n_6545),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_6492),
.Y(n_6570)
);

INVx2_ASAP7_75t_L g6571 ( 
.A(n_6500),
.Y(n_6571)
);

HB1xp67_ASAP7_75t_L g6572 ( 
.A(n_6500),
.Y(n_6572)
);

NAND2xp5_ASAP7_75t_SL g6573 ( 
.A(n_6516),
.B(n_6457),
.Y(n_6573)
);

AND2x2_ASAP7_75t_L g6574 ( 
.A(n_6514),
.B(n_6460),
.Y(n_6574)
);

INVx2_ASAP7_75t_SL g6575 ( 
.A(n_6505),
.Y(n_6575)
);

NOR2xp33_ASAP7_75t_L g6576 ( 
.A(n_6535),
.B(n_6400),
.Y(n_6576)
);

NAND2xp5_ASAP7_75t_L g6577 ( 
.A(n_6485),
.B(n_6444),
.Y(n_6577)
);

INVx2_ASAP7_75t_L g6578 ( 
.A(n_6525),
.Y(n_6578)
);

OAI21xp5_ASAP7_75t_L g6579 ( 
.A1(n_6524),
.A2(n_6373),
.B(n_6440),
.Y(n_6579)
);

NOR3xp33_ASAP7_75t_SL g6580 ( 
.A(n_6501),
.B(n_6458),
.C(n_6445),
.Y(n_6580)
);

INVx2_ASAP7_75t_L g6581 ( 
.A(n_6496),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6484),
.Y(n_6582)
);

NAND2xp5_ASAP7_75t_L g6583 ( 
.A(n_6526),
.B(n_6437),
.Y(n_6583)
);

AOI221xp5_ASAP7_75t_L g6584 ( 
.A1(n_6509),
.A2(n_6433),
.B1(n_6435),
.B2(n_6461),
.C(n_6448),
.Y(n_6584)
);

NAND2xp5_ASAP7_75t_L g6585 ( 
.A(n_6527),
.B(n_6465),
.Y(n_6585)
);

NAND2xp5_ASAP7_75t_L g6586 ( 
.A(n_6539),
.B(n_6418),
.Y(n_6586)
);

NAND2xp5_ASAP7_75t_SL g6587 ( 
.A(n_6502),
.B(n_6528),
.Y(n_6587)
);

INVx2_ASAP7_75t_SL g6588 ( 
.A(n_6538),
.Y(n_6588)
);

INVx2_ASAP7_75t_L g6589 ( 
.A(n_6497),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_6499),
.Y(n_6590)
);

AOI21xp5_ASAP7_75t_L g6591 ( 
.A1(n_6517),
.A2(n_6466),
.B(n_6386),
.Y(n_6591)
);

NAND2xp5_ASAP7_75t_L g6592 ( 
.A(n_6542),
.B(n_6363),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6483),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_6545),
.Y(n_6594)
);

AOI322xp5_ASAP7_75t_L g6595 ( 
.A1(n_6543),
.A2(n_709),
.A3(n_708),
.B1(n_706),
.B2(n_704),
.C1(n_705),
.C2(n_707),
.Y(n_6595)
);

INVx1_ASAP7_75t_L g6596 ( 
.A(n_6494),
.Y(n_6596)
);

NAND2x1_ASAP7_75t_L g6597 ( 
.A(n_6504),
.B(n_704),
.Y(n_6597)
);

NAND2x1_ASAP7_75t_L g6598 ( 
.A(n_6519),
.B(n_704),
.Y(n_6598)
);

OR2x2_ASAP7_75t_L g6599 ( 
.A(n_6522),
.B(n_705),
.Y(n_6599)
);

OAI21xp33_ASAP7_75t_SL g6600 ( 
.A1(n_6487),
.A2(n_705),
.B(n_706),
.Y(n_6600)
);

OR2x2_ASAP7_75t_L g6601 ( 
.A(n_6506),
.B(n_706),
.Y(n_6601)
);

INVx1_ASAP7_75t_L g6602 ( 
.A(n_6541),
.Y(n_6602)
);

INVx2_ASAP7_75t_L g6603 ( 
.A(n_6534),
.Y(n_6603)
);

INVxp33_ASAP7_75t_L g6604 ( 
.A(n_6529),
.Y(n_6604)
);

NAND2xp5_ASAP7_75t_L g6605 ( 
.A(n_6495),
.B(n_707),
.Y(n_6605)
);

OR2x2_ASAP7_75t_L g6606 ( 
.A(n_6518),
.B(n_708),
.Y(n_6606)
);

INVx1_ASAP7_75t_L g6607 ( 
.A(n_6544),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6549),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_6536),
.Y(n_6609)
);

OR2x2_ASAP7_75t_L g6610 ( 
.A(n_6548),
.B(n_708),
.Y(n_6610)
);

AND2x2_ASAP7_75t_L g6611 ( 
.A(n_6520),
.B(n_710),
.Y(n_6611)
);

AND2x2_ASAP7_75t_L g6612 ( 
.A(n_6481),
.B(n_710),
.Y(n_6612)
);

NAND2xp5_ASAP7_75t_L g6613 ( 
.A(n_6482),
.B(n_711),
.Y(n_6613)
);

OR2x2_ASAP7_75t_L g6614 ( 
.A(n_6512),
.B(n_712),
.Y(n_6614)
);

NAND2xp33_ASAP7_75t_L g6615 ( 
.A(n_6515),
.B(n_712),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_6508),
.B(n_712),
.Y(n_6616)
);

INVxp67_ASAP7_75t_L g6617 ( 
.A(n_6546),
.Y(n_6617)
);

AOI22xp33_ASAP7_75t_L g6618 ( 
.A1(n_6523),
.A2(n_715),
.B1(n_713),
.B2(n_714),
.Y(n_6618)
);

INVx2_ASAP7_75t_L g6619 ( 
.A(n_6532),
.Y(n_6619)
);

AND2x2_ASAP7_75t_L g6620 ( 
.A(n_6533),
.B(n_713),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_6540),
.Y(n_6621)
);

AND2x2_ASAP7_75t_L g6622 ( 
.A(n_6547),
.B(n_6530),
.Y(n_6622)
);

INVxp67_ASAP7_75t_SL g6623 ( 
.A(n_6531),
.Y(n_6623)
);

INVx6_ASAP7_75t_L g6624 ( 
.A(n_6488),
.Y(n_6624)
);

INVx1_ASAP7_75t_L g6625 ( 
.A(n_6491),
.Y(n_6625)
);

AND2x2_ASAP7_75t_L g6626 ( 
.A(n_6521),
.B(n_713),
.Y(n_6626)
);

AND2x2_ASAP7_75t_L g6627 ( 
.A(n_6486),
.B(n_714),
.Y(n_6627)
);

INVx1_ASAP7_75t_L g6628 ( 
.A(n_6564),
.Y(n_6628)
);

INVx2_ASAP7_75t_SL g6629 ( 
.A(n_6557),
.Y(n_6629)
);

NAND2xp5_ASAP7_75t_SL g6630 ( 
.A(n_6550),
.B(n_714),
.Y(n_6630)
);

OAI22xp5_ASAP7_75t_L g6631 ( 
.A1(n_6569),
.A2(n_718),
.B1(n_716),
.B2(n_717),
.Y(n_6631)
);

AOI22xp33_ASAP7_75t_L g6632 ( 
.A1(n_6572),
.A2(n_718),
.B1(n_716),
.B2(n_717),
.Y(n_6632)
);

OR2x2_ASAP7_75t_L g6633 ( 
.A(n_6594),
.B(n_716),
.Y(n_6633)
);

INVxp33_ASAP7_75t_L g6634 ( 
.A(n_6563),
.Y(n_6634)
);

INVx2_ASAP7_75t_SL g6635 ( 
.A(n_6557),
.Y(n_6635)
);

OR2x2_ASAP7_75t_L g6636 ( 
.A(n_6597),
.B(n_717),
.Y(n_6636)
);

A2O1A1Ixp33_ASAP7_75t_L g6637 ( 
.A1(n_6595),
.A2(n_721),
.B(n_719),
.C(n_720),
.Y(n_6637)
);

INVx2_ASAP7_75t_L g6638 ( 
.A(n_6571),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_6598),
.Y(n_6639)
);

A2O1A1Ixp33_ASAP7_75t_L g6640 ( 
.A1(n_6600),
.A2(n_722),
.B(n_719),
.C(n_721),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_6567),
.Y(n_6641)
);

INVx2_ASAP7_75t_L g6642 ( 
.A(n_6578),
.Y(n_6642)
);

NAND2xp5_ASAP7_75t_SL g6643 ( 
.A(n_6575),
.B(n_719),
.Y(n_6643)
);

OAI31xp33_ASAP7_75t_SL g6644 ( 
.A1(n_6623),
.A2(n_724),
.A3(n_722),
.B(n_723),
.Y(n_6644)
);

A2O1A1Ixp33_ASAP7_75t_L g6645 ( 
.A1(n_6565),
.A2(n_725),
.B(n_722),
.C(n_724),
.Y(n_6645)
);

HB1xp67_ASAP7_75t_L g6646 ( 
.A(n_6552),
.Y(n_6646)
);

OR2x2_ASAP7_75t_L g6647 ( 
.A(n_6556),
.B(n_724),
.Y(n_6647)
);

AND2x4_ASAP7_75t_SL g6648 ( 
.A(n_6603),
.B(n_725),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6620),
.Y(n_6649)
);

INVx1_ASAP7_75t_L g6650 ( 
.A(n_6553),
.Y(n_6650)
);

A2O1A1Ixp33_ASAP7_75t_L g6651 ( 
.A1(n_6576),
.A2(n_727),
.B(n_725),
.C(n_726),
.Y(n_6651)
);

AOI32xp33_ASAP7_75t_L g6652 ( 
.A1(n_6554),
.A2(n_728),
.A3(n_726),
.B1(n_727),
.B2(n_729),
.Y(n_6652)
);

NAND2xp5_ASAP7_75t_L g6653 ( 
.A(n_6612),
.B(n_727),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_6559),
.Y(n_6654)
);

AOI22xp5_ASAP7_75t_L g6655 ( 
.A1(n_6588),
.A2(n_730),
.B1(n_728),
.B2(n_729),
.Y(n_6655)
);

OAI22xp33_ASAP7_75t_L g6656 ( 
.A1(n_6562),
.A2(n_6590),
.B1(n_6608),
.B2(n_6607),
.Y(n_6656)
);

INVx1_ASAP7_75t_SL g6657 ( 
.A(n_6581),
.Y(n_6657)
);

AOI21xp33_ASAP7_75t_SL g6658 ( 
.A1(n_6573),
.A2(n_728),
.B(n_729),
.Y(n_6658)
);

INVx2_ASAP7_75t_L g6659 ( 
.A(n_6589),
.Y(n_6659)
);

AND2x2_ASAP7_75t_L g6660 ( 
.A(n_6561),
.B(n_730),
.Y(n_6660)
);

NOR2xp33_ASAP7_75t_L g6661 ( 
.A(n_6613),
.B(n_730),
.Y(n_6661)
);

OR2x2_ASAP7_75t_L g6662 ( 
.A(n_6605),
.B(n_731),
.Y(n_6662)
);

NOR3x1_ASAP7_75t_L g6663 ( 
.A(n_6579),
.B(n_731),
.C(n_732),
.Y(n_6663)
);

INVxp67_ASAP7_75t_SL g6664 ( 
.A(n_6616),
.Y(n_6664)
);

NOR2xp33_ASAP7_75t_L g6665 ( 
.A(n_6570),
.B(n_732),
.Y(n_6665)
);

INVx2_ASAP7_75t_L g6666 ( 
.A(n_6619),
.Y(n_6666)
);

NAND2xp5_ASAP7_75t_L g6667 ( 
.A(n_6611),
.B(n_732),
.Y(n_6667)
);

AOI21xp33_ASAP7_75t_SL g6668 ( 
.A1(n_6587),
.A2(n_733),
.B(n_734),
.Y(n_6668)
);

AOI32xp33_ASAP7_75t_L g6669 ( 
.A1(n_6551),
.A2(n_735),
.A3(n_733),
.B1(n_734),
.B2(n_736),
.Y(n_6669)
);

OAI221xp5_ASAP7_75t_L g6670 ( 
.A1(n_6618),
.A2(n_736),
.B1(n_734),
.B2(n_735),
.C(n_737),
.Y(n_6670)
);

NAND2xp5_ASAP7_75t_L g6671 ( 
.A(n_6555),
.B(n_735),
.Y(n_6671)
);

INVxp67_ASAP7_75t_SL g6672 ( 
.A(n_6577),
.Y(n_6672)
);

NAND2xp5_ASAP7_75t_L g6673 ( 
.A(n_6627),
.B(n_736),
.Y(n_6673)
);

INVxp67_ASAP7_75t_L g6674 ( 
.A(n_6626),
.Y(n_6674)
);

AOI21xp5_ASAP7_75t_L g6675 ( 
.A1(n_6615),
.A2(n_737),
.B(n_738),
.Y(n_6675)
);

AND2x2_ASAP7_75t_L g6676 ( 
.A(n_6558),
.B(n_739),
.Y(n_6676)
);

AOI322xp5_ASAP7_75t_L g6677 ( 
.A1(n_6621),
.A2(n_744),
.A3(n_743),
.B1(n_741),
.B2(n_739),
.C1(n_740),
.C2(n_742),
.Y(n_6677)
);

INVx1_ASAP7_75t_L g6678 ( 
.A(n_6574),
.Y(n_6678)
);

INVxp67_ASAP7_75t_SL g6679 ( 
.A(n_6629),
.Y(n_6679)
);

INVx4_ASAP7_75t_L g6680 ( 
.A(n_6638),
.Y(n_6680)
);

INVx2_ASAP7_75t_L g6681 ( 
.A(n_6635),
.Y(n_6681)
);

INVx1_ASAP7_75t_L g6682 ( 
.A(n_6628),
.Y(n_6682)
);

NAND2xp5_ASAP7_75t_L g6683 ( 
.A(n_6657),
.B(n_6566),
.Y(n_6683)
);

NAND2xp5_ASAP7_75t_L g6684 ( 
.A(n_6642),
.B(n_6580),
.Y(n_6684)
);

NAND2xp5_ASAP7_75t_L g6685 ( 
.A(n_6677),
.B(n_6659),
.Y(n_6685)
);

XOR2x2_ASAP7_75t_L g6686 ( 
.A(n_6653),
.B(n_6586),
.Y(n_6686)
);

INVx2_ASAP7_75t_L g6687 ( 
.A(n_6666),
.Y(n_6687)
);

NAND4xp25_ASAP7_75t_L g6688 ( 
.A(n_6678),
.B(n_6584),
.C(n_6641),
.D(n_6654),
.Y(n_6688)
);

INVx1_ASAP7_75t_L g6689 ( 
.A(n_6636),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_6633),
.Y(n_6690)
);

INVx1_ASAP7_75t_SL g6691 ( 
.A(n_6648),
.Y(n_6691)
);

XOR2x2_ASAP7_75t_L g6692 ( 
.A(n_6667),
.B(n_6585),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_6646),
.Y(n_6693)
);

INVxp67_ASAP7_75t_SL g6694 ( 
.A(n_6656),
.Y(n_6694)
);

AND2x2_ASAP7_75t_L g6695 ( 
.A(n_6660),
.B(n_6602),
.Y(n_6695)
);

INVx1_ASAP7_75t_L g6696 ( 
.A(n_6647),
.Y(n_6696)
);

AND2x2_ASAP7_75t_L g6697 ( 
.A(n_6676),
.B(n_6609),
.Y(n_6697)
);

NOR2xp33_ASAP7_75t_L g6698 ( 
.A(n_6634),
.B(n_6617),
.Y(n_6698)
);

AOI32xp33_ASAP7_75t_L g6699 ( 
.A1(n_6650),
.A2(n_6604),
.A3(n_6596),
.B1(n_6622),
.B2(n_6625),
.Y(n_6699)
);

OA21x2_ASAP7_75t_L g6700 ( 
.A1(n_6671),
.A2(n_6591),
.B(n_6582),
.Y(n_6700)
);

OAI21x1_ASAP7_75t_SL g6701 ( 
.A1(n_6658),
.A2(n_6592),
.B(n_6583),
.Y(n_6701)
);

AND2x2_ASAP7_75t_L g6702 ( 
.A(n_6672),
.B(n_6560),
.Y(n_6702)
);

NAND2x1p5_ASAP7_75t_L g6703 ( 
.A(n_6663),
.B(n_6610),
.Y(n_6703)
);

NAND2xp5_ASAP7_75t_L g6704 ( 
.A(n_6644),
.B(n_6593),
.Y(n_6704)
);

INVx1_ASAP7_75t_L g6705 ( 
.A(n_6631),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6673),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6655),
.Y(n_6707)
);

NAND2xp5_ASAP7_75t_L g6708 ( 
.A(n_6632),
.B(n_6599),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_6662),
.Y(n_6709)
);

OAI21x1_ASAP7_75t_SL g6710 ( 
.A1(n_6639),
.A2(n_6601),
.B(n_6614),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_6649),
.B(n_6606),
.Y(n_6711)
);

AND2x2_ASAP7_75t_L g6712 ( 
.A(n_6674),
.B(n_6661),
.Y(n_6712)
);

NAND2xp5_ASAP7_75t_SL g6713 ( 
.A(n_6668),
.B(n_6568),
.Y(n_6713)
);

NAND2xp5_ASAP7_75t_L g6714 ( 
.A(n_6640),
.B(n_6669),
.Y(n_6714)
);

AND2x2_ASAP7_75t_L g6715 ( 
.A(n_6665),
.B(n_6624),
.Y(n_6715)
);

INVxp33_ASAP7_75t_L g6716 ( 
.A(n_6630),
.Y(n_6716)
);

OR2x2_ASAP7_75t_L g6717 ( 
.A(n_6643),
.B(n_740),
.Y(n_6717)
);

AND4x1_ASAP7_75t_L g6718 ( 
.A(n_6651),
.B(n_6624),
.C(n_742),
.D(n_740),
.Y(n_6718)
);

INVxp67_ASAP7_75t_L g6719 ( 
.A(n_6670),
.Y(n_6719)
);

NAND2xp5_ASAP7_75t_L g6720 ( 
.A(n_6652),
.B(n_741),
.Y(n_6720)
);

INVxp67_ASAP7_75t_L g6721 ( 
.A(n_6675),
.Y(n_6721)
);

NAND2xp5_ASAP7_75t_L g6722 ( 
.A(n_6637),
.B(n_741),
.Y(n_6722)
);

AND2x2_ASAP7_75t_L g6723 ( 
.A(n_6664),
.B(n_6668),
.Y(n_6723)
);

NAND2xp5_ASAP7_75t_L g6724 ( 
.A(n_6645),
.B(n_742),
.Y(n_6724)
);

INVx1_ASAP7_75t_L g6725 ( 
.A(n_6629),
.Y(n_6725)
);

NAND2x1_ASAP7_75t_SL g6726 ( 
.A(n_6628),
.B(n_743),
.Y(n_6726)
);

CKINVDCx20_ASAP7_75t_R g6727 ( 
.A(n_6629),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_L g6728 ( 
.A(n_6629),
.B(n_744),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6629),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6629),
.Y(n_6730)
);

AND2x2_ASAP7_75t_L g6731 ( 
.A(n_6629),
.B(n_744),
.Y(n_6731)
);

HB1xp67_ASAP7_75t_L g6732 ( 
.A(n_6629),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6629),
.Y(n_6733)
);

NAND2xp5_ASAP7_75t_L g6734 ( 
.A(n_6629),
.B(n_745),
.Y(n_6734)
);

XNOR2xp5_ASAP7_75t_L g6735 ( 
.A(n_6629),
.B(n_745),
.Y(n_6735)
);

XNOR2x2_ASAP7_75t_L g6736 ( 
.A(n_6657),
.B(n_745),
.Y(n_6736)
);

XOR2x2_ASAP7_75t_L g6737 ( 
.A(n_6735),
.B(n_746),
.Y(n_6737)
);

AND2x2_ASAP7_75t_SL g6738 ( 
.A(n_6680),
.B(n_746),
.Y(n_6738)
);

NAND2xp5_ASAP7_75t_L g6739 ( 
.A(n_6694),
.B(n_6679),
.Y(n_6739)
);

INVx2_ASAP7_75t_L g6740 ( 
.A(n_6680),
.Y(n_6740)
);

O2A1O1Ixp5_ASAP7_75t_L g6741 ( 
.A1(n_6681),
.A2(n_6687),
.B(n_6729),
.C(n_6725),
.Y(n_6741)
);

NAND2xp5_ASAP7_75t_L g6742 ( 
.A(n_6732),
.B(n_747),
.Y(n_6742)
);

BUFx2_ASAP7_75t_L g6743 ( 
.A(n_6727),
.Y(n_6743)
);

NOR2xp33_ASAP7_75t_L g6744 ( 
.A(n_6730),
.B(n_747),
.Y(n_6744)
);

OAI21xp33_ASAP7_75t_SL g6745 ( 
.A1(n_6688),
.A2(n_747),
.B(n_748),
.Y(n_6745)
);

NAND2x1_ASAP7_75t_L g6746 ( 
.A(n_6733),
.B(n_748),
.Y(n_6746)
);

NAND2xp5_ASAP7_75t_L g6747 ( 
.A(n_6731),
.B(n_749),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_6683),
.Y(n_6748)
);

AND3x2_ASAP7_75t_L g6749 ( 
.A(n_6721),
.B(n_749),
.C(n_750),
.Y(n_6749)
);

AOI22xp5_ASAP7_75t_L g6750 ( 
.A1(n_6698),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.Y(n_6750)
);

INVx1_ASAP7_75t_L g6751 ( 
.A(n_6702),
.Y(n_6751)
);

AND2x2_ASAP7_75t_L g6752 ( 
.A(n_6697),
.B(n_750),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_6728),
.Y(n_6753)
);

XOR2xp5_ASAP7_75t_L g6754 ( 
.A(n_6692),
.B(n_751),
.Y(n_6754)
);

INVx1_ASAP7_75t_L g6755 ( 
.A(n_6734),
.Y(n_6755)
);

INVxp67_ASAP7_75t_L g6756 ( 
.A(n_6684),
.Y(n_6756)
);

OAI21xp5_ASAP7_75t_SL g6757 ( 
.A1(n_6699),
.A2(n_752),
.B(n_753),
.Y(n_6757)
);

NAND2xp5_ASAP7_75t_L g6758 ( 
.A(n_6691),
.B(n_752),
.Y(n_6758)
);

AND2x2_ASAP7_75t_L g6759 ( 
.A(n_6695),
.B(n_753),
.Y(n_6759)
);

A2O1A1Ixp33_ASAP7_75t_L g6760 ( 
.A1(n_6693),
.A2(n_755),
.B(n_753),
.C(n_754),
.Y(n_6760)
);

XNOR2x1_ASAP7_75t_L g6761 ( 
.A(n_6736),
.B(n_754),
.Y(n_6761)
);

NAND2xp5_ASAP7_75t_L g6762 ( 
.A(n_6682),
.B(n_754),
.Y(n_6762)
);

NAND2xp5_ASAP7_75t_L g6763 ( 
.A(n_6689),
.B(n_755),
.Y(n_6763)
);

AND2x2_ASAP7_75t_L g6764 ( 
.A(n_6715),
.B(n_755),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6685),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_6720),
.Y(n_6766)
);

NAND2xp5_ASAP7_75t_L g6767 ( 
.A(n_6719),
.B(n_756),
.Y(n_6767)
);

HB1xp67_ASAP7_75t_L g6768 ( 
.A(n_6739),
.Y(n_6768)
);

NOR2x1_ASAP7_75t_L g6769 ( 
.A(n_6757),
.B(n_6705),
.Y(n_6769)
);

NAND2xp5_ASAP7_75t_L g6770 ( 
.A(n_6751),
.B(n_6726),
.Y(n_6770)
);

OAI211xp5_ASAP7_75t_L g6771 ( 
.A1(n_6745),
.A2(n_6722),
.B(n_6704),
.C(n_6714),
.Y(n_6771)
);

NAND2xp5_ASAP7_75t_SL g6772 ( 
.A(n_6740),
.B(n_6724),
.Y(n_6772)
);

INVxp67_ASAP7_75t_L g6773 ( 
.A(n_6743),
.Y(n_6773)
);

INVx1_ASAP7_75t_SL g6774 ( 
.A(n_6748),
.Y(n_6774)
);

AND2x2_ASAP7_75t_L g6775 ( 
.A(n_6764),
.B(n_6700),
.Y(n_6775)
);

INVx1_ASAP7_75t_L g6776 ( 
.A(n_6741),
.Y(n_6776)
);

INVx1_ASAP7_75t_SL g6777 ( 
.A(n_6746),
.Y(n_6777)
);

NAND2xp5_ASAP7_75t_L g6778 ( 
.A(n_6749),
.B(n_6690),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6758),
.Y(n_6779)
);

INVx2_ASAP7_75t_L g6780 ( 
.A(n_6756),
.Y(n_6780)
);

AOI22xp33_ASAP7_75t_L g6781 ( 
.A1(n_6765),
.A2(n_6707),
.B1(n_6696),
.B2(n_6723),
.Y(n_6781)
);

XNOR2xp5_ASAP7_75t_L g6782 ( 
.A(n_6754),
.B(n_6686),
.Y(n_6782)
);

OR2x2_ASAP7_75t_L g6783 ( 
.A(n_6747),
.B(n_6703),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_6752),
.Y(n_6784)
);

INVx1_ASAP7_75t_L g6785 ( 
.A(n_6759),
.Y(n_6785)
);

NAND3xp33_ASAP7_75t_L g6786 ( 
.A(n_6744),
.B(n_6718),
.C(n_6713),
.Y(n_6786)
);

OAI21xp5_ASAP7_75t_SL g6787 ( 
.A1(n_6750),
.A2(n_6716),
.B(n_6711),
.Y(n_6787)
);

A2O1A1Ixp33_ASAP7_75t_L g6788 ( 
.A1(n_6742),
.A2(n_6717),
.B(n_6709),
.C(n_6708),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6763),
.Y(n_6789)
);

INVx1_ASAP7_75t_L g6790 ( 
.A(n_6762),
.Y(n_6790)
);

INVx1_ASAP7_75t_SL g6791 ( 
.A(n_6738),
.Y(n_6791)
);

OAI22xp5_ASAP7_75t_SL g6792 ( 
.A1(n_6767),
.A2(n_6700),
.B1(n_6706),
.B2(n_6701),
.Y(n_6792)
);

INVx1_ASAP7_75t_L g6793 ( 
.A(n_6761),
.Y(n_6793)
);

NOR2xp67_ASAP7_75t_SL g6794 ( 
.A(n_6776),
.B(n_6766),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_6775),
.Y(n_6795)
);

NAND2x1p5_ASAP7_75t_L g6796 ( 
.A(n_6774),
.B(n_6753),
.Y(n_6796)
);

NOR3xp33_ASAP7_75t_L g6797 ( 
.A(n_6771),
.B(n_6760),
.C(n_6755),
.Y(n_6797)
);

NAND2xp5_ASAP7_75t_L g6798 ( 
.A(n_6768),
.B(n_6712),
.Y(n_6798)
);

AND2x2_ASAP7_75t_L g6799 ( 
.A(n_6773),
.B(n_6737),
.Y(n_6799)
);

NAND3xp33_ASAP7_75t_L g6800 ( 
.A(n_6781),
.B(n_6710),
.C(n_756),
.Y(n_6800)
);

INVx1_ASAP7_75t_L g6801 ( 
.A(n_6792),
.Y(n_6801)
);

NAND2xp5_ASAP7_75t_L g6802 ( 
.A(n_6780),
.B(n_6777),
.Y(n_6802)
);

NAND2xp5_ASAP7_75t_L g6803 ( 
.A(n_6784),
.B(n_757),
.Y(n_6803)
);

NOR2xp33_ASAP7_75t_L g6804 ( 
.A(n_6785),
.B(n_6787),
.Y(n_6804)
);

INVx1_ASAP7_75t_L g6805 ( 
.A(n_6782),
.Y(n_6805)
);

INVx1_ASAP7_75t_L g6806 ( 
.A(n_6769),
.Y(n_6806)
);

NAND4xp75_ASAP7_75t_L g6807 ( 
.A(n_6772),
.B(n_759),
.C(n_757),
.D(n_758),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_6783),
.Y(n_6808)
);

OAI322xp33_ASAP7_75t_L g6809 ( 
.A1(n_6778),
.A2(n_757),
.A3(n_758),
.B1(n_759),
.B2(n_760),
.C1(n_761),
.C2(n_762),
.Y(n_6809)
);

NAND3xp33_ASAP7_75t_L g6810 ( 
.A(n_6786),
.B(n_758),
.C(n_760),
.Y(n_6810)
);

NOR2xp33_ASAP7_75t_L g6811 ( 
.A(n_6793),
.B(n_760),
.Y(n_6811)
);

NAND2xp5_ASAP7_75t_L g6812 ( 
.A(n_6788),
.B(n_761),
.Y(n_6812)
);

NOR2x1_ASAP7_75t_L g6813 ( 
.A(n_6770),
.B(n_761),
.Y(n_6813)
);

AOI21xp5_ASAP7_75t_L g6814 ( 
.A1(n_6779),
.A2(n_762),
.B(n_763),
.Y(n_6814)
);

OAI22xp33_ASAP7_75t_L g6815 ( 
.A1(n_6791),
.A2(n_765),
.B1(n_763),
.B2(n_764),
.Y(n_6815)
);

OAI22xp5_ASAP7_75t_L g6816 ( 
.A1(n_6795),
.A2(n_6789),
.B1(n_6790),
.B2(n_765),
.Y(n_6816)
);

AOI221xp5_ASAP7_75t_L g6817 ( 
.A1(n_6809),
.A2(n_766),
.B1(n_763),
.B2(n_764),
.C(n_767),
.Y(n_6817)
);

AOI31xp33_ASAP7_75t_L g6818 ( 
.A1(n_6801),
.A2(n_767),
.A3(n_764),
.B(n_766),
.Y(n_6818)
);

NAND2x1p5_ASAP7_75t_L g6819 ( 
.A(n_6794),
.B(n_766),
.Y(n_6819)
);

AOI22xp33_ASAP7_75t_L g6820 ( 
.A1(n_6808),
.A2(n_770),
.B1(n_768),
.B2(n_769),
.Y(n_6820)
);

O2A1O1Ixp5_ASAP7_75t_L g6821 ( 
.A1(n_6798),
.A2(n_770),
.B(n_768),
.C(n_769),
.Y(n_6821)
);

O2A1O1Ixp33_ASAP7_75t_L g6822 ( 
.A1(n_6815),
.A2(n_772),
.B(n_770),
.C(n_771),
.Y(n_6822)
);

AOI21xp33_ASAP7_75t_L g6823 ( 
.A1(n_6802),
.A2(n_772),
.B(n_773),
.Y(n_6823)
);

INVxp67_ASAP7_75t_L g6824 ( 
.A(n_6812),
.Y(n_6824)
);

AOI21xp33_ASAP7_75t_L g6825 ( 
.A1(n_6810),
.A2(n_773),
.B(n_774),
.Y(n_6825)
);

OAI22xp5_ASAP7_75t_L g6826 ( 
.A1(n_6800),
.A2(n_775),
.B1(n_773),
.B2(n_774),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_6796),
.Y(n_6827)
);

A2O1A1Ixp33_ASAP7_75t_L g6828 ( 
.A1(n_6811),
.A2(n_776),
.B(n_774),
.C(n_775),
.Y(n_6828)
);

NAND2xp5_ASAP7_75t_L g6829 ( 
.A(n_6814),
.B(n_6805),
.Y(n_6829)
);

BUFx6f_ASAP7_75t_L g6830 ( 
.A(n_6806),
.Y(n_6830)
);

AOI221xp5_ASAP7_75t_L g6831 ( 
.A1(n_6804),
.A2(n_777),
.B1(n_775),
.B2(n_776),
.C(n_778),
.Y(n_6831)
);

OAI22xp5_ASAP7_75t_L g6832 ( 
.A1(n_6803),
.A2(n_778),
.B1(n_776),
.B2(n_777),
.Y(n_6832)
);

OAI21xp33_ASAP7_75t_L g6833 ( 
.A1(n_6799),
.A2(n_777),
.B(n_778),
.Y(n_6833)
);

AO22x2_ASAP7_75t_L g6834 ( 
.A1(n_6807),
.A2(n_781),
.B1(n_779),
.B2(n_780),
.Y(n_6834)
);

AOI22xp33_ASAP7_75t_L g6835 ( 
.A1(n_6797),
.A2(n_6813),
.B1(n_781),
.B2(n_779),
.Y(n_6835)
);

NAND2xp5_ASAP7_75t_SL g6836 ( 
.A(n_6795),
.B(n_779),
.Y(n_6836)
);

OAI22xp33_ASAP7_75t_SL g6837 ( 
.A1(n_6795),
.A2(n_782),
.B1(n_780),
.B2(n_781),
.Y(n_6837)
);

INVx1_ASAP7_75t_L g6838 ( 
.A(n_6795),
.Y(n_6838)
);

INVx1_ASAP7_75t_L g6839 ( 
.A(n_6795),
.Y(n_6839)
);

NOR4xp25_ASAP7_75t_L g6840 ( 
.A(n_6833),
.B(n_783),
.C(n_780),
.D(n_782),
.Y(n_6840)
);

AND5x1_ASAP7_75t_L g6841 ( 
.A(n_6817),
.B(n_785),
.C(n_782),
.D(n_784),
.E(n_786),
.Y(n_6841)
);

NOR3xp33_ASAP7_75t_L g6842 ( 
.A(n_6838),
.B(n_784),
.C(n_785),
.Y(n_6842)
);

NOR2xp33_ASAP7_75t_L g6843 ( 
.A(n_6839),
.B(n_784),
.Y(n_6843)
);

NAND3xp33_ASAP7_75t_L g6844 ( 
.A(n_6823),
.B(n_786),
.C(n_787),
.Y(n_6844)
);

AND2x2_ASAP7_75t_SL g6845 ( 
.A(n_6827),
.B(n_786),
.Y(n_6845)
);

OA22x2_ASAP7_75t_L g6846 ( 
.A1(n_6826),
.A2(n_789),
.B1(n_787),
.B2(n_788),
.Y(n_6846)
);

NAND3xp33_ASAP7_75t_L g6847 ( 
.A(n_6835),
.B(n_787),
.C(n_788),
.Y(n_6847)
);

OAI211xp5_ASAP7_75t_SL g6848 ( 
.A1(n_6831),
.A2(n_790),
.B(n_788),
.C(n_789),
.Y(n_6848)
);

NOR2xp33_ASAP7_75t_L g6849 ( 
.A(n_6830),
.B(n_790),
.Y(n_6849)
);

A2O1A1Ixp33_ASAP7_75t_L g6850 ( 
.A1(n_6822),
.A2(n_792),
.B(n_790),
.C(n_791),
.Y(n_6850)
);

NAND2x1_ASAP7_75t_L g6851 ( 
.A(n_6830),
.B(n_791),
.Y(n_6851)
);

AND2x4_ASAP7_75t_L g6852 ( 
.A(n_6829),
.B(n_791),
.Y(n_6852)
);

NAND4xp25_ASAP7_75t_L g6853 ( 
.A(n_6820),
.B(n_794),
.C(n_792),
.D(n_793),
.Y(n_6853)
);

NOR2xp33_ASAP7_75t_L g6854 ( 
.A(n_6836),
.B(n_792),
.Y(n_6854)
);

NOR3x1_ASAP7_75t_L g6855 ( 
.A(n_6832),
.B(n_793),
.C(n_794),
.Y(n_6855)
);

NAND4xp75_ASAP7_75t_L g6856 ( 
.A(n_6821),
.B(n_795),
.C(n_793),
.D(n_794),
.Y(n_6856)
);

NOR3xp33_ASAP7_75t_L g6857 ( 
.A(n_6816),
.B(n_795),
.C(n_796),
.Y(n_6857)
);

INVx1_ASAP7_75t_SL g6858 ( 
.A(n_6819),
.Y(n_6858)
);

AND2x2_ASAP7_75t_L g6859 ( 
.A(n_6834),
.B(n_796),
.Y(n_6859)
);

AND4x1_ASAP7_75t_L g6860 ( 
.A(n_6828),
.B(n_799),
.C(n_797),
.D(n_798),
.Y(n_6860)
);

NAND2xp5_ASAP7_75t_L g6861 ( 
.A(n_6818),
.B(n_6837),
.Y(n_6861)
);

OR5x1_ASAP7_75t_L g6862 ( 
.A(n_6825),
.B(n_799),
.C(n_797),
.D(n_798),
.E(n_800),
.Y(n_6862)
);

NAND3xp33_ASAP7_75t_L g6863 ( 
.A(n_6824),
.B(n_797),
.C(n_798),
.Y(n_6863)
);

AND2x2_ASAP7_75t_L g6864 ( 
.A(n_6838),
.B(n_800),
.Y(n_6864)
);

AOI22xp5_ASAP7_75t_L g6865 ( 
.A1(n_6838),
.A2(n_802),
.B1(n_800),
.B2(n_801),
.Y(n_6865)
);

NOR2x2_ASAP7_75t_L g6866 ( 
.A(n_6856),
.B(n_801),
.Y(n_6866)
);

AOI211xp5_ASAP7_75t_L g6867 ( 
.A1(n_6843),
.A2(n_804),
.B(n_802),
.C(n_803),
.Y(n_6867)
);

AOI22xp5_ASAP7_75t_L g6868 ( 
.A1(n_6864),
.A2(n_804),
.B1(n_802),
.B2(n_803),
.Y(n_6868)
);

OAI211xp5_ASAP7_75t_SL g6869 ( 
.A1(n_6861),
.A2(n_807),
.B(n_805),
.C(n_806),
.Y(n_6869)
);

AOI211xp5_ASAP7_75t_L g6870 ( 
.A1(n_6848),
.A2(n_6853),
.B(n_6844),
.C(n_6854),
.Y(n_6870)
);

AND2x2_ASAP7_75t_L g6871 ( 
.A(n_6859),
.B(n_805),
.Y(n_6871)
);

OAI32xp33_ASAP7_75t_L g6872 ( 
.A1(n_6857),
.A2(n_807),
.A3(n_805),
.B1(n_806),
.B2(n_808),
.Y(n_6872)
);

OA22x2_ASAP7_75t_L g6873 ( 
.A1(n_6852),
.A2(n_6858),
.B1(n_6865),
.B2(n_6851),
.Y(n_6873)
);

AOI211xp5_ASAP7_75t_L g6874 ( 
.A1(n_6842),
.A2(n_6863),
.B(n_6847),
.C(n_6849),
.Y(n_6874)
);

AOI322xp5_ASAP7_75t_L g6875 ( 
.A1(n_6852),
.A2(n_808),
.A3(n_809),
.B1(n_810),
.B2(n_811),
.C1(n_812),
.C2(n_813),
.Y(n_6875)
);

OAI21xp5_ASAP7_75t_SL g6876 ( 
.A1(n_6850),
.A2(n_809),
.B(n_810),
.Y(n_6876)
);

OAI21xp33_ASAP7_75t_L g6877 ( 
.A1(n_6840),
.A2(n_810),
.B(n_811),
.Y(n_6877)
);

INVxp33_ASAP7_75t_L g6878 ( 
.A(n_6846),
.Y(n_6878)
);

AOI21xp5_ASAP7_75t_L g6879 ( 
.A1(n_6845),
.A2(n_811),
.B(n_812),
.Y(n_6879)
);

AOI221x1_ASAP7_75t_L g6880 ( 
.A1(n_6841),
.A2(n_814),
.B1(n_812),
.B2(n_813),
.C(n_815),
.Y(n_6880)
);

XNOR2xp5_ASAP7_75t_L g6881 ( 
.A(n_6860),
.B(n_6862),
.Y(n_6881)
);

INVx1_ASAP7_75t_L g6882 ( 
.A(n_6855),
.Y(n_6882)
);

HB1xp67_ASAP7_75t_L g6883 ( 
.A(n_6871),
.Y(n_6883)
);

OAI211xp5_ASAP7_75t_SL g6884 ( 
.A1(n_6870),
.A2(n_815),
.B(n_813),
.C(n_814),
.Y(n_6884)
);

OAI21xp5_ASAP7_75t_SL g6885 ( 
.A1(n_6878),
.A2(n_814),
.B(n_816),
.Y(n_6885)
);

NOR2x1_ASAP7_75t_L g6886 ( 
.A(n_6882),
.B(n_6876),
.Y(n_6886)
);

NOR4xp25_ASAP7_75t_L g6887 ( 
.A(n_6869),
.B(n_818),
.C(n_816),
.D(n_817),
.Y(n_6887)
);

OR2x2_ASAP7_75t_L g6888 ( 
.A(n_6868),
.B(n_816),
.Y(n_6888)
);

NAND2xp5_ASAP7_75t_L g6889 ( 
.A(n_6875),
.B(n_817),
.Y(n_6889)
);

NOR3xp33_ASAP7_75t_L g6890 ( 
.A(n_6867),
.B(n_818),
.C(n_819),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_6872),
.Y(n_6891)
);

AO22x2_ASAP7_75t_L g6892 ( 
.A1(n_6880),
.A2(n_821),
.B1(n_819),
.B2(n_820),
.Y(n_6892)
);

HB1xp67_ASAP7_75t_L g6893 ( 
.A(n_6881),
.Y(n_6893)
);

XNOR2xp5_ASAP7_75t_L g6894 ( 
.A(n_6873),
.B(n_819),
.Y(n_6894)
);

AOI221xp5_ASAP7_75t_L g6895 ( 
.A1(n_6885),
.A2(n_6879),
.B1(n_6877),
.B2(n_6874),
.C(n_6866),
.Y(n_6895)
);

AOI22xp33_ASAP7_75t_L g6896 ( 
.A1(n_6893),
.A2(n_6883),
.B1(n_6886),
.B2(n_6894),
.Y(n_6896)
);

INVx1_ASAP7_75t_L g6897 ( 
.A(n_6892),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6892),
.Y(n_6898)
);

NOR3xp33_ASAP7_75t_SL g6899 ( 
.A(n_6884),
.B(n_820),
.C(n_821),
.Y(n_6899)
);

AOI21xp5_ASAP7_75t_L g6900 ( 
.A1(n_6897),
.A2(n_6898),
.B(n_6887),
.Y(n_6900)
);

A2O1A1Ixp33_ASAP7_75t_L g6901 ( 
.A1(n_6895),
.A2(n_6888),
.B(n_6889),
.C(n_6890),
.Y(n_6901)
);

NOR2x1_ASAP7_75t_SL g6902 ( 
.A(n_6896),
.B(n_6891),
.Y(n_6902)
);

INVx1_ASAP7_75t_SL g6903 ( 
.A(n_6899),
.Y(n_6903)
);

NOR4xp25_ASAP7_75t_L g6904 ( 
.A(n_6903),
.B(n_822),
.C(n_820),
.D(n_821),
.Y(n_6904)
);

OAI22xp5_ASAP7_75t_L g6905 ( 
.A1(n_6901),
.A2(n_825),
.B1(n_823),
.B2(n_824),
.Y(n_6905)
);

AND2x4_ASAP7_75t_L g6906 ( 
.A(n_6904),
.B(n_6902),
.Y(n_6906)
);

AOI22xp5_ASAP7_75t_L g6907 ( 
.A1(n_6906),
.A2(n_6900),
.B1(n_6905),
.B2(n_825),
.Y(n_6907)
);

OAI22xp5_ASAP7_75t_L g6908 ( 
.A1(n_6907),
.A2(n_825),
.B1(n_823),
.B2(n_824),
.Y(n_6908)
);

AOI21xp5_ASAP7_75t_L g6909 ( 
.A1(n_6908),
.A2(n_865),
.B(n_864),
.Y(n_6909)
);

AOI221xp5_ASAP7_75t_L g6910 ( 
.A1(n_6909),
.A2(n_826),
.B1(n_823),
.B2(n_824),
.C(n_827),
.Y(n_6910)
);

OAI22xp5_ASAP7_75t_L g6911 ( 
.A1(n_6910),
.A2(n_866),
.B1(n_867),
.B2(n_865),
.Y(n_6911)
);

OAI21xp5_ASAP7_75t_L g6912 ( 
.A1(n_6911),
.A2(n_869),
.B(n_866),
.Y(n_6912)
);

BUFx2_ASAP7_75t_L g6913 ( 
.A(n_6912),
.Y(n_6913)
);

OR2x6_ASAP7_75t_L g6914 ( 
.A(n_6913),
.B(n_871),
.Y(n_6914)
);

AOI22xp5_ASAP7_75t_L g6915 ( 
.A1(n_6914),
.A2(n_872),
.B1(n_873),
.B2(n_871),
.Y(n_6915)
);

AOI211xp5_ASAP7_75t_L g6916 ( 
.A1(n_6915),
.A2(n_873),
.B(n_876),
.C(n_872),
.Y(n_6916)
);


endmodule