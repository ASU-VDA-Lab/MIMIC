module fake_jpeg_16623_n_396 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_46),
.Y(n_84)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_79),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_17),
.A2(n_14),
.B(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_51),
.B(n_54),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_53),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_14),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_21),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_57),
.Y(n_137)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_60),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_75),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_30),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_22),
.B(n_13),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_42),
.B1(n_37),
.B2(n_22),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_85),
.A2(n_102),
.B1(n_108),
.B2(n_1),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_89),
.B(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_29),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_44),
.A2(n_42),
.B1(n_37),
.B2(n_24),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_61),
.C(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_114),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_58),
.A2(n_39),
.B1(n_32),
.B2(n_29),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_SL g167 ( 
.A(n_104),
.B(n_125),
.C(n_35),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_42),
.B1(n_70),
.B2(n_67),
.Y(n_108)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_49),
.B(n_32),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_110),
.B(n_112),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_24),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_55),
.B(n_24),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_113),
.B(n_123),
.Y(n_171)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_39),
.B1(n_25),
.B2(n_27),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_117),
.A2(n_126),
.B1(n_129),
.B2(n_133),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_38),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_38),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_48),
.A2(n_39),
.B1(n_37),
.B2(n_25),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_50),
.A2(n_27),
.B1(n_40),
.B2(n_34),
.Y(n_129)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_63),
.A2(n_27),
.B1(n_40),
.B2(n_3),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_64),
.B(n_34),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_134),
.B(n_41),
.Y(n_185)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_28),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_66),
.B(n_31),
.Y(n_139)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

OR2x2_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_31),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_140),
.A2(n_147),
.B(n_117),
.C(n_126),
.Y(n_190)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_20),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_145),
.B(n_185),
.Y(n_216)
);

OR2x2_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_20),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_81),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_155),
.Y(n_195)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_88),
.A2(n_100),
.B1(n_135),
.B2(n_106),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_173),
.B1(n_15),
.B2(n_11),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_87),
.B(n_73),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_84),
.B(n_28),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_168),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_104),
.A2(n_41),
.B(n_9),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_157),
.A2(n_11),
.B(n_4),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_92),
.Y(n_158)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_101),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_166),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_97),
.Y(n_166)
);

OAI211xp5_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_96),
.B(n_15),
.C(n_86),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_1),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_92),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_35),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_177),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_90),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_178),
.Y(n_220)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_35),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_115),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_183),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_2),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_188),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g181 ( 
.A1(n_106),
.A2(n_15),
.B1(n_35),
.B2(n_30),
.Y(n_181)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_119),
.A2(n_30),
.B1(n_41),
.B2(n_35),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_107),
.B1(n_95),
.B2(n_5),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_88),
.A2(n_15),
.B1(n_11),
.B2(n_9),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_168),
.B1(n_180),
.B2(n_173),
.Y(n_210)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_99),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_103),
.B(n_2),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_190),
.B(n_219),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_146),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_203),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_100),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_196),
.B(n_201),
.C(n_206),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_185),
.A2(n_95),
.B1(n_107),
.B2(n_114),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_231),
.B(n_183),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_198),
.B(n_213),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_96),
.Y(n_201)
);

OA22x2_ASAP7_75t_L g270 ( 
.A1(n_202),
.A2(n_210),
.B1(n_205),
.B2(n_231),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_150),
.B1(n_170),
.B2(n_6),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_155),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_146),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_218),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_159),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_131),
.B1(n_121),
.B2(n_93),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_225),
.B1(n_227),
.B2(n_158),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_148),
.Y(n_218)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_157),
.A2(n_131),
.B1(n_121),
.B2(n_93),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_156),
.A2(n_96),
.B1(n_118),
.B2(n_91),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_91),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_229),
.B(n_2),
.Y(n_262)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_142),
.Y(n_232)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g275 ( 
.A1(n_234),
.A2(n_242),
.B(n_243),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_147),
.B(n_153),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_237),
.A2(n_252),
.B(n_198),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_145),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_240),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_145),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_171),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_257),
.C(n_268),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_163),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_244),
.B(n_245),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_162),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_141),
.B1(n_172),
.B2(n_182),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_247),
.A2(n_250),
.B1(n_256),
.B2(n_263),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_182),
.B1(n_181),
.B2(n_169),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_140),
.B(n_165),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_201),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_255),
.B(n_264),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_182),
.B1(n_181),
.B2(n_151),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_197),
.B(n_86),
.C(n_151),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_187),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_262),
.B(n_207),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_216),
.A2(n_215),
.B1(n_210),
.B2(n_190),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_223),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_216),
.B(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_225),
.A2(n_6),
.B1(n_7),
.B2(n_202),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_266),
.A2(n_243),
.B1(n_240),
.B2(n_247),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_208),
.A2(n_6),
.B(n_7),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_SL g300 ( 
.A1(n_267),
.A2(n_269),
.B(n_259),
.C(n_265),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_227),
.C(n_209),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_205),
.A2(n_209),
.B1(n_218),
.B2(n_193),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_193),
.B1(n_230),
.B2(n_199),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_221),
.B(n_191),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_285),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_290),
.B(n_298),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_213),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_282),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_294),
.B1(n_296),
.B2(n_297),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_212),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_291),
.C(n_241),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_246),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_287),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_199),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_288),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_222),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_223),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_270),
.A2(n_226),
.B1(n_233),
.B2(n_232),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_194),
.B1(n_226),
.B2(n_257),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_194),
.B1(n_242),
.B2(n_245),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_239),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_255),
.B1(n_238),
.B2(n_266),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_283),
.B(n_294),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_235),
.B(n_268),
.Y(n_301)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_303),
.A2(n_306),
.B(n_324),
.Y(n_342)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_300),
.A2(n_234),
.B(n_252),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_275),
.A2(n_248),
.B1(n_244),
.B2(n_256),
.Y(n_308)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_297),
.A2(n_248),
.B1(n_250),
.B2(n_258),
.Y(n_310)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_320),
.C(n_322),
.Y(n_327)
);

AOI22x1_ASAP7_75t_L g312 ( 
.A1(n_293),
.A2(n_267),
.B1(n_235),
.B2(n_239),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_312),
.A2(n_319),
.B1(n_314),
.B2(n_318),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_237),
.Y(n_313)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_314),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_253),
.Y(n_315)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_290),
.A2(n_253),
.B1(n_293),
.B2(n_296),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_319),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_284),
.C(n_274),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_276),
.C(n_281),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_278),
.A2(n_300),
.B(n_276),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_299),
.C(n_289),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.C(n_286),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_277),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_332),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_324),
.B(n_288),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_280),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_336),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_308),
.B(n_280),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_316),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_337),
.B(n_321),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_320),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_343),
.C(n_323),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_302),
.A2(n_303),
.B(n_312),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_317),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_305),
.C(n_326),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_344),
.A2(n_304),
.B1(n_310),
.B2(n_309),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_348),
.A2(n_351),
.B1(n_353),
.B2(n_358),
.Y(n_368)
);

AO21x1_ASAP7_75t_L g349 ( 
.A1(n_342),
.A2(n_302),
.B(n_312),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_354),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_306),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_356),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_334),
.B(n_305),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_331),
.B(n_325),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_315),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_355),
.A2(n_359),
.B1(n_362),
.B2(n_346),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_343),
.C(n_327),
.Y(n_370)
);

INVx11_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_309),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_335),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_361),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_336),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

BUFx12_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_363),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_346),
.B1(n_345),
.B2(n_339),
.Y(n_364)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_372),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_371),
.C(n_373),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_327),
.C(n_332),
.Y(n_371)
);

FAx1_ASAP7_75t_SL g372 ( 
.A(n_354),
.B(n_342),
.CI(n_329),
.CON(n_372),
.SN(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_349),
.A2(n_356),
.B1(n_360),
.B2(n_347),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_369),
.A2(n_350),
.B(n_361),
.Y(n_376)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_376),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_371),
.A2(n_352),
.B(n_347),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_380),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_352),
.C(n_370),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_374),
.A2(n_364),
.B1(n_369),
.B2(n_373),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_383),
.B(n_384),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_378),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_366),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_378),
.C(n_365),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_386),
.A2(n_387),
.B(n_382),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_368),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_384),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_389),
.A2(n_390),
.B1(n_386),
.B2(n_375),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_391),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_392),
.B(n_377),
.Y(n_393)
);

AO21x1_ASAP7_75t_L g394 ( 
.A1(n_393),
.A2(n_372),
.B(n_363),
.Y(n_394)
);

A2O1A1Ixp33_ASAP7_75t_L g395 ( 
.A1(n_394),
.A2(n_372),
.B(n_365),
.C(n_363),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_385),
.Y(n_396)
);


endmodule