module real_aes_7676_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_693;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_224;
wire n_639;
wire n_587;
wire n_546;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_0), .A2(n_205), .B1(n_510), .B2(n_513), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_1), .A2(n_196), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_2), .A2(n_89), .B1(n_517), .B2(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_3), .B(n_291), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_4), .A2(n_134), .B1(n_281), .B2(n_297), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_5), .A2(n_23), .B1(n_310), .B2(n_584), .Y(n_612) );
INVx1_ASAP7_75t_L g727 ( .A(n_6), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_7), .A2(n_220), .B1(n_356), .B2(n_358), .C(n_360), .Y(n_355) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_8), .A2(n_182), .B1(n_480), .B2(n_544), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_9), .B(n_638), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_10), .A2(n_21), .B1(n_475), .B2(n_476), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_11), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_12), .Y(n_532) );
AOI222xp33_ASAP7_75t_L g370 ( .A1(n_13), .A2(n_105), .B1(n_131), .B2(n_294), .C1(n_371), .C2(n_373), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g239 ( .A1(n_14), .A2(n_114), .B1(n_240), .B2(n_255), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_15), .A2(n_119), .B1(n_429), .B2(n_498), .Y(n_497) );
OA22x2_ASAP7_75t_L g451 ( .A1(n_16), .A2(n_452), .B1(n_453), .B2(n_484), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_16), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_17), .A2(n_157), .B1(n_240), .B2(n_447), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_18), .A2(n_99), .B1(n_305), .B2(n_405), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_19), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_20), .A2(n_193), .B1(n_479), .B2(n_480), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_22), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_24), .A2(n_213), .B1(n_275), .B2(n_280), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_25), .Y(n_397) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_26), .A2(n_70), .B1(n_244), .B2(n_249), .Y(n_252) );
INVx1_ASAP7_75t_L g694 ( .A(n_26), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_27), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_28), .A2(n_33), .B1(n_374), .B2(n_434), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_29), .A2(n_52), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_30), .A2(n_195), .B1(n_345), .B2(n_630), .C(n_631), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_31), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g642 ( .A1(n_32), .A2(n_86), .B1(n_132), .B2(n_373), .C1(n_643), .C2(n_644), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_34), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_35), .A2(n_48), .B1(n_570), .B2(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_36), .A2(n_214), .B1(n_294), .B2(n_297), .Y(n_293) );
AOI222xp33_ASAP7_75t_L g613 ( .A1(n_37), .A2(n_106), .B1(n_163), .B2(n_495), .C1(n_570), .C2(n_571), .Y(n_613) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_38), .A2(n_72), .B1(n_244), .B2(n_245), .Y(n_254) );
INVx1_ASAP7_75t_L g695 ( .A(n_38), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_39), .Y(n_351) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_40), .A2(n_194), .B1(n_304), .B2(n_522), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_41), .A2(n_103), .B1(n_260), .B2(n_604), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_42), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_43), .A2(n_221), .B1(n_260), .B2(n_264), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_44), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_45), .A2(n_67), .B1(n_504), .B2(n_506), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_46), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_47), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_49), .A2(n_198), .B1(n_403), .B2(n_611), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_50), .A2(n_490), .B1(n_491), .B2(n_525), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_50), .Y(n_490) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_51), .A2(n_113), .B1(n_280), .B2(n_297), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_53), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_54), .A2(n_107), .B1(n_401), .B2(n_403), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_55), .A2(n_158), .B1(n_308), .B2(n_447), .Y(n_714) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_56), .A2(n_96), .B1(n_405), .B2(n_406), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_57), .A2(n_118), .B1(n_619), .B2(n_621), .C(n_623), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_58), .B(n_357), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_59), .A2(n_120), .B1(n_637), .B2(n_638), .C(n_639), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_60), .A2(n_184), .B1(n_350), .B2(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_61), .A2(n_212), .B1(n_294), .B2(n_374), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_62), .B(n_285), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_63), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_64), .A2(n_129), .B1(n_255), .B2(n_512), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_65), .A2(n_318), .B1(n_375), .B2(n_376), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_65), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_66), .A2(n_617), .B1(n_645), .B2(n_646), .Y(n_616) );
INVx1_ASAP7_75t_L g645 ( .A(n_66), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_68), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_69), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_71), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_73), .Y(n_325) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_74), .A2(n_174), .B1(n_446), .B2(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g229 ( .A(n_75), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_76), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_77), .A2(n_116), .B1(n_374), .B2(n_393), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_78), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_79), .A2(n_178), .B1(n_426), .B2(n_464), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_80), .A2(n_95), .B1(n_580), .B2(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g226 ( .A(n_81), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_82), .A2(n_156), .B1(n_255), .B2(n_512), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_83), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_84), .A2(n_117), .B1(n_479), .B2(n_611), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_85), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_87), .A2(n_137), .B1(n_357), .B2(n_436), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_88), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g432 ( .A1(n_90), .A2(n_110), .B1(n_433), .B2(n_434), .Y(n_432) );
OA22x2_ASAP7_75t_L g378 ( .A1(n_91), .A2(n_379), .B1(n_380), .B2(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_91), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_92), .A2(n_93), .B1(n_515), .B2(n_517), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_94), .A2(n_109), .B1(n_297), .B2(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_97), .A2(n_177), .B1(n_401), .B2(n_580), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_98), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_100), .A2(n_133), .B1(n_240), .B2(n_604), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_101), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_102), .A2(n_180), .B1(n_306), .B2(n_583), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_104), .A2(n_148), .B1(n_323), .B2(n_401), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g438 ( .A1(n_108), .A2(n_183), .B1(n_412), .B2(n_439), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_111), .A2(n_179), .B1(n_677), .B2(n_679), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_112), .Y(n_664) );
INVx2_ASAP7_75t_L g230 ( .A(n_115), .Y(n_230) );
INVx1_ASAP7_75t_L g548 ( .A(n_121), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_122), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_123), .B(n_291), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_124), .B(n_285), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_125), .A2(n_216), .B1(n_582), .B2(n_584), .Y(n_581) );
AND2x6_ASAP7_75t_L g225 ( .A(n_126), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_126), .Y(n_688) );
AO22x2_ASAP7_75t_L g243 ( .A1(n_127), .A2(n_187), .B1(n_244), .B2(n_245), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_128), .A2(n_172), .B1(n_240), .B2(n_345), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_130), .A2(n_208), .B1(n_275), .B2(n_280), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_135), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_136), .A2(n_197), .B1(n_264), .B2(n_409), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_138), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_139), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_140), .A2(n_176), .B1(n_295), .B2(n_297), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_141), .B(n_356), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_142), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_143), .B(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_144), .Y(n_624) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_145), .A2(n_153), .B1(n_411), .B2(n_412), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_146), .A2(n_698), .B1(n_699), .B2(n_715), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_146), .Y(n_715) );
AO22x2_ASAP7_75t_L g248 ( .A1(n_147), .A2(n_200), .B1(n_244), .B2(n_249), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_149), .A2(n_219), .B1(n_308), .B2(n_310), .Y(n_307) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_150), .A2(n_201), .B1(n_409), .B2(n_513), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_151), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_152), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_154), .B(n_436), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_155), .A2(n_185), .B1(n_308), .B2(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_159), .A2(n_162), .B1(n_255), .B2(n_737), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_160), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_161), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_164), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g301 ( .A1(n_165), .A2(n_217), .B1(n_302), .B2(n_305), .Y(n_301) );
AOI22xp33_ASAP7_75t_SL g441 ( .A1(n_166), .A2(n_169), .B1(n_334), .B2(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_167), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_168), .A2(n_170), .B1(n_411), .B2(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_171), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_173), .B(n_291), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_175), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_181), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_186), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_187), .B(n_693), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_188), .Y(n_650) );
OA22x2_ASAP7_75t_L g419 ( .A1(n_189), .A2(n_420), .B1(n_421), .B2(n_449), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_189), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_190), .A2(n_223), .B(n_231), .C(n_696), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_191), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_192), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_199), .Y(n_706) );
INVx1_ASAP7_75t_L g691 ( .A(n_200), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_202), .Y(n_496) );
OA22x2_ASAP7_75t_L g555 ( .A1(n_203), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_555) );
CKINVDCx16_ASAP7_75t_R g556 ( .A(n_203), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_204), .B(n_356), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_206), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_207), .Y(n_654) );
INVx1_ASAP7_75t_L g244 ( .A(n_209), .Y(n_244) );
INVx1_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_210), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_211), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_215), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_218), .Y(n_424) );
INVx2_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_226), .Y(n_687) );
OA21x2_ASAP7_75t_L g720 ( .A1(n_227), .A2(n_686), .B(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_594), .B1(n_681), .B2(n_682), .C(n_683), .Y(n_231) );
INVx1_ASAP7_75t_L g681 ( .A(n_232), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_553), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_414), .B1(n_415), .B2(n_552), .Y(n_233) );
INVx1_ASAP7_75t_L g552 ( .A(n_234), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_314), .B1(n_315), .B2(n_413), .Y(n_234) );
INVx1_ASAP7_75t_L g413 ( .A(n_235), .Y(n_413) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
XOR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_313), .Y(n_236) );
NAND3x1_ASAP7_75t_L g237 ( .A(n_238), .B(n_266), .C(n_300), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_259), .Y(n_238) );
BUFx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx3_ASAP7_75t_L g409 ( .A(n_241), .Y(n_409) );
BUFx3_ASAP7_75t_L g440 ( .A(n_241), .Y(n_440) );
BUFx3_ASAP7_75t_L g522 ( .A(n_241), .Y(n_522) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_250), .Y(n_241) );
AND2x2_ASAP7_75t_L g312 ( .A(n_242), .B(n_292), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_242), .B(n_292), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_242), .B(n_250), .Y(n_354) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_243), .B(n_248), .Y(n_258) );
INVx2_ASAP7_75t_L g263 ( .A(n_243), .Y(n_263) );
AND2x2_ASAP7_75t_L g279 ( .A(n_243), .B(n_252), .Y(n_279) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g249 ( .A(n_246), .Y(n_249) );
INVx1_ASAP7_75t_L g282 ( .A(n_247), .Y(n_282) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g262 ( .A(n_248), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g273 ( .A(n_248), .Y(n_273) );
INVx1_ASAP7_75t_L g278 ( .A(n_248), .Y(n_278) );
AND2x4_ASAP7_75t_L g261 ( .A(n_250), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g265 ( .A(n_250), .B(n_257), .Y(n_265) );
AND2x2_ASAP7_75t_L g309 ( .A(n_250), .B(n_272), .Y(n_309) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
OR2x2_ASAP7_75t_L g289 ( .A(n_251), .B(n_254), .Y(n_289) );
AND2x2_ASAP7_75t_L g292 ( .A(n_251), .B(n_254), .Y(n_292) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g271 ( .A(n_252), .B(n_254), .Y(n_271) );
INVx1_ASAP7_75t_L g256 ( .A(n_253), .Y(n_256) );
AND2x2_ASAP7_75t_L g296 ( .A(n_253), .B(n_278), .Y(n_296) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_256), .B(n_279), .Y(n_364) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x6_ASAP7_75t_L g336 ( .A(n_258), .B(n_299), .Y(n_336) );
BUFx2_ASAP7_75t_L g679 ( .A(n_260), .Y(n_679) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx3_ASAP7_75t_L g324 ( .A(n_261), .Y(n_324) );
BUFx3_ASAP7_75t_L g403 ( .A(n_261), .Y(n_403) );
INVx2_ASAP7_75t_L g483 ( .A(n_261), .Y(n_483) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_261), .Y(n_512) );
AND2x4_ASAP7_75t_L g287 ( .A(n_262), .B(n_288), .Y(n_287) );
AND2x6_ASAP7_75t_L g291 ( .A(n_262), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g387 ( .A(n_262), .Y(n_387) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_262), .B(n_292), .Y(n_390) );
AND2x2_ASAP7_75t_L g272 ( .A(n_263), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g628 ( .A(n_264), .Y(n_628) );
BUFx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
BUFx3_ASAP7_75t_L g327 ( .A(n_265), .Y(n_327) );
BUFx3_ASAP7_75t_L g447 ( .A(n_265), .Y(n_447) );
BUFx2_ASAP7_75t_SL g480 ( .A(n_265), .Y(n_480) );
BUFx2_ASAP7_75t_L g513 ( .A(n_265), .Y(n_513) );
INVx1_ASAP7_75t_L g593 ( .A(n_265), .Y(n_593) );
BUFx3_ASAP7_75t_L g602 ( .A(n_265), .Y(n_602) );
NOR2x1_ASAP7_75t_L g266 ( .A(n_267), .B(n_283), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_274), .Y(n_267) );
BUFx2_ASAP7_75t_L g372 ( .A(n_269), .Y(n_372) );
INVx4_ASAP7_75t_L g643 ( .A(n_269), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_269), .A2(n_706), .B(n_707), .Y(n_705) );
INVx4_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx3_ASAP7_75t_L g395 ( .A(n_270), .Y(n_395) );
INVx2_ASAP7_75t_L g462 ( .A(n_270), .Y(n_462) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_270), .Y(n_495) );
INVx2_ASAP7_75t_SL g659 ( .A(n_270), .Y(n_659) );
AND2x6_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x4_ASAP7_75t_L g281 ( .A(n_271), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g368 ( .A(n_271), .Y(n_368) );
AND2x6_ASAP7_75t_L g304 ( .A(n_272), .B(n_288), .Y(n_304) );
AND2x4_ASAP7_75t_L g306 ( .A(n_272), .B(n_292), .Y(n_306) );
BUFx4f_ASAP7_75t_L g429 ( .A(n_275), .Y(n_429) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx12f_ASAP7_75t_L g374 ( .A(n_276), .Y(n_374) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_276), .Y(n_466) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g295 ( .A(n_279), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g297 ( .A(n_279), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g507 ( .A(n_280), .Y(n_507) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx3_ASAP7_75t_L g434 ( .A(n_281), .Y(n_434) );
INVx1_ASAP7_75t_L g369 ( .A(n_282), .Y(n_369) );
NAND3xp33_ASAP7_75t_L g283 ( .A(n_284), .B(n_290), .C(n_293), .Y(n_283) );
BUFx2_ASAP7_75t_L g637 ( .A(n_285), .Y(n_637) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx5_ASAP7_75t_L g357 ( .A(n_286), .Y(n_357) );
INVx2_ASAP7_75t_L g536 ( .A(n_286), .Y(n_536) );
INVx4_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g386 ( .A(n_289), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g359 ( .A(n_291), .Y(n_359) );
BUFx2_ASAP7_75t_L g436 ( .A(n_291), .Y(n_436) );
BUFx4f_ASAP7_75t_L g638 ( .A(n_291), .Y(n_638) );
BUFx4f_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_295), .Y(n_393) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_295), .Y(n_426) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_295), .Y(n_539) );
BUFx2_ASAP7_75t_L g433 ( .A(n_297), .Y(n_433) );
INVx1_ASAP7_75t_L g505 ( .A(n_297), .Y(n_505) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_307), .Y(n_300) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g446 ( .A(n_303), .Y(n_446) );
INVx5_ASAP7_75t_SL g544 ( .A(n_303), .Y(n_544) );
INVx2_ASAP7_75t_L g580 ( .A(n_303), .Y(n_580) );
INVx4_ASAP7_75t_L g626 ( .A(n_303), .Y(n_626) );
INVx11_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx11_ASAP7_75t_L g342 ( .A(n_304), .Y(n_342) );
BUFx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx6_ASAP7_75t_L g346 ( .A(n_306), .Y(n_346) );
BUFx3_ASAP7_75t_L g412 ( .A(n_306), .Y(n_412) );
BUFx3_ASAP7_75t_L g670 ( .A(n_306), .Y(n_670) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_308), .Y(n_520) );
INVx3_ASAP7_75t_L g620 ( .A(n_308), .Y(n_620) );
BUFx3_ASAP7_75t_L g669 ( .A(n_308), .Y(n_669) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_SL g350 ( .A(n_309), .Y(n_350) );
INVx2_ASAP7_75t_L g402 ( .A(n_309), .Y(n_402) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx5_ASAP7_75t_L g405 ( .A(n_311), .Y(n_405) );
INVx1_ASAP7_75t_L g443 ( .A(n_311), .Y(n_443) );
BUFx3_ASAP7_75t_L g516 ( .A(n_311), .Y(n_516) );
INVx4_ASAP7_75t_L g583 ( .A(n_311), .Y(n_583) );
INVx2_ASAP7_75t_L g737 ( .A(n_311), .Y(n_737) );
INVx8_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_377), .B2(n_378), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g376 ( .A(n_318), .Y(n_376) );
AND4x1_ASAP7_75t_L g318 ( .A(n_319), .B(n_337), .C(n_355), .D(n_370), .Y(n_318) );
NOR2xp33_ASAP7_75t_SL g319 ( .A(n_320), .B(n_328), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_325), .B2(n_326), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVxp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B1(n_332), .B2(n_333), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_330), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
BUFx2_ASAP7_75t_R g330 ( .A(n_331), .Y(n_330) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g406 ( .A(n_335), .Y(n_406) );
BUFx2_ASAP7_75t_L g584 ( .A(n_335), .Y(n_584) );
BUFx2_ASAP7_75t_L g635 ( .A(n_335), .Y(n_635) );
INVx6_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g476 ( .A(n_336), .Y(n_476) );
INVx1_ASAP7_75t_SL g517 ( .A(n_336), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_347), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_343), .B2(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx4_ASAP7_75t_L g411 ( .A(n_342), .Y(n_411) );
INVx4_ASAP7_75t_L g479 ( .A(n_342), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_344), .A2(n_586), .B1(n_587), .B2(n_588), .Y(n_585) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g524 ( .A(n_346), .Y(n_524) );
INVx3_ASAP7_75t_L g611 ( .A(n_346), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_351), .B2(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g588 ( .A(n_353), .Y(n_588) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_365), .B2(n_366), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_362), .A2(n_366), .B1(n_640), .B2(n_641), .Y(n_639) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx4_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_367), .B1(n_397), .B2(n_398), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_364), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_455) );
OAI22xp33_ASAP7_75t_SL g573 ( .A1(n_364), .A2(n_574), .B1(n_575), .B2(n_576), .Y(n_573) );
BUFx3_ASAP7_75t_L g663 ( .A(n_364), .Y(n_663) );
BUFx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_367), .Y(n_459) );
OR2x6_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI222xp33_ASAP7_75t_L g423 ( .A1(n_372), .A2(n_424), .B1(n_425), .B2(n_427), .C1(n_428), .C2(n_430), .Y(n_423) );
BUFx4f_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g572 ( .A(n_374), .Y(n_572) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND3x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_399), .C(n_407), .Y(n_381) );
NOR3xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_391), .C(n_396), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_388), .B2(n_389), .Y(n_383) );
BUFx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_386), .Y(n_469) );
BUFx3_ASAP7_75t_L g564 ( .A(n_389), .Y(n_564) );
OAI22xp5_ASAP7_75t_SL g653 ( .A1(n_389), .A2(n_469), .B1(n_654), .B2(n_655), .Y(n_653) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g472 ( .A(n_390), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx4_ASAP7_75t_L g499 ( .A(n_393), .Y(n_499) );
BUFx2_ASAP7_75t_L g570 ( .A(n_393), .Y(n_570) );
INVx3_ASAP7_75t_L g567 ( .A(n_395), .Y(n_567) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_404), .Y(n_399) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g604 ( .A(n_402), .Y(n_604) );
INVx1_ASAP7_75t_L g591 ( .A(n_403), .Y(n_591) );
BUFx2_ASAP7_75t_L g475 ( .A(n_405), .Y(n_475) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g622 ( .A(n_409), .Y(n_622) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_485), .B1(n_550), .B2(n_551), .Y(n_415) );
INVx1_ASAP7_75t_L g550 ( .A(n_416), .Y(n_550) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_450), .B2(n_451), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g449 ( .A(n_421), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_437), .C(n_444), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_431), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
OAI222xp33_ASAP7_75t_L g656 ( .A1(n_428), .A2(n_657), .B1(n_658), .B2(n_659), .C1(n_660), .C2(n_661), .Y(n_656) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
BUFx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g484 ( .A(n_453), .Y(n_484) );
NAND2x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_473), .Y(n_453) );
NOR3xp33_ASAP7_75t_SL g454 ( .A(n_455), .B(n_460), .C(n_467), .Y(n_454) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g575 ( .A(n_459), .Y(n_575) );
OAI21xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_463), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_462), .A2(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_470), .B2(n_471), .Y(n_467) );
INVx1_ASAP7_75t_L g562 ( .A(n_469), .Y(n_562) );
OA211x2_ASAP7_75t_L g605 ( .A1(n_471), .A2(n_606), .B(n_607), .C(n_608), .Y(n_605) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND4x1_ASAP7_75t_L g473 ( .A(n_474), .B(n_477), .C(n_478), .D(n_481), .Y(n_473) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g551 ( .A(n_485), .Y(n_551) );
OAI22xp5_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_487), .B1(n_526), .B2(n_549), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g525 ( .A(n_491), .Y(n_525) );
NAND3x1_ASAP7_75t_L g491 ( .A(n_492), .B(n_508), .C(n_518), .Y(n_491) );
NOR2x1_ASAP7_75t_L g492 ( .A(n_493), .B(n_500), .Y(n_492) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_496), .B(n_497), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .C(n_503), .Y(n_500) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .Y(n_508) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx4_ASAP7_75t_L g630 ( .A(n_511), .Y(n_630) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
BUFx4f_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g678 ( .A(n_522), .Y(n_678) );
INVx1_ASAP7_75t_L g549 ( .A(n_526), .Y(n_549) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
XOR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_548), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_530), .B(n_540), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .C(n_538), .Y(n_534) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_539), .Y(n_644) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_577), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_566), .C(n_573), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI21xp33_ASAP7_75t_SL g566 ( .A1(n_567), .A2(n_568), .B(n_569), .Y(n_566) );
OAI21xp5_ASAP7_75t_SL g726 ( .A1(n_567), .A2(n_727), .B(n_728), .Y(n_726) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI22xp5_ASAP7_75t_SL g662 ( .A1(n_575), .A2(n_663), .B1(n_664), .B2(n_665), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_585), .C(n_589), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g673 ( .A(n_583), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_592), .B2(n_593), .Y(n_589) );
INVx1_ASAP7_75t_L g682 ( .A(n_594), .Y(n_682) );
AOI22xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_648), .B1(n_649), .B2(n_680), .Y(n_594) );
INVx1_ASAP7_75t_L g680 ( .A(n_595), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_615), .B1(n_616), .B2(n_647), .Y(n_595) );
INVx1_ASAP7_75t_L g647 ( .A(n_596), .Y(n_647) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
XOR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_614), .Y(n_598) );
NAND4xp75_ASAP7_75t_L g599 ( .A(n_600), .B(n_605), .C(n_609), .D(n_613), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g646 ( .A(n_617), .Y(n_646) );
AND4x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_629), .C(n_636), .D(n_642), .Y(n_617) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_627), .B2(n_628), .Y(n_623) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_SL g657 ( .A(n_644), .Y(n_657) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
XNOR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_666), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_656), .C(n_662), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_674), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .Y(n_667) );
INVx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_685), .B(n_689), .Y(n_684) );
OR2x2_ASAP7_75t_SL g743 ( .A(n_685), .B(n_690), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_686), .Y(n_717) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_687), .B(n_719), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g719 ( .A(n_688), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
OAI322xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_716), .A3(n_718), .B1(n_720), .B2(n_722), .C1(n_723), .C2(n_741), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND3x1_ASAP7_75t_SL g700 ( .A(n_701), .B(n_704), .C(n_712), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_705), .B(n_708), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .C(n_711), .Y(n_708) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
BUFx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
XOR2x2_ASAP7_75t_L g723 ( .A(n_722), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_725), .B(n_733), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_729), .Y(n_725) );
NAND3xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .C(n_732), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_738), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
endmodule