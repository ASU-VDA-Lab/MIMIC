module fake_jpeg_12711_n_582 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_582);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_582;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx3_ASAP7_75t_SL g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_2),
.B(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_66),
.B(n_68),
.Y(n_144)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g143 ( 
.A(n_69),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_13),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_70),
.B(n_71),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_74),
.B(n_84),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_76),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_83),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_12),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_50),
.Y(n_89)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_12),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_90),
.B(n_93),
.Y(n_157)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_95),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_34),
.B(n_11),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_97),
.B(n_111),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_34),
.B(n_11),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_123),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_17),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_103),
.Y(n_127)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

BUFx12f_ASAP7_75t_SL g111 ( 
.A(n_23),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_17),
.Y(n_113)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_40),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_31),
.Y(n_124)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_90),
.B(n_55),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_149),
.B(n_155),
.Y(n_270)
);

BUFx4f_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_66),
.B(n_55),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_156),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_81),
.A2(n_28),
.B1(n_59),
.B2(n_40),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_166),
.A2(n_45),
.B1(n_21),
.B2(n_47),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_SL g168 ( 
.A1(n_114),
.A2(n_38),
.B(n_26),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_201),
.Y(n_209)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_95),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_84),
.B(n_59),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_92),
.B(n_51),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_62),
.Y(n_199)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_63),
.Y(n_200)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_95),
.B(n_38),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_38),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_202),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_204),
.B(n_208),
.Y(n_278)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_178),
.B(n_105),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g211 ( 
.A(n_145),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_211),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_212),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_202),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_214),
.B(n_228),
.Y(n_314)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_216),
.Y(n_305)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_191),
.A2(n_106),
.B1(n_38),
.B2(n_99),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_219),
.A2(n_229),
.B1(n_230),
.B2(n_271),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_221),
.B(n_243),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_222),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_41),
.B1(n_51),
.B2(n_94),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_224),
.A2(n_258),
.B(n_29),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_183),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_225),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_89),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_260),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_139),
.B(n_41),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_140),
.A2(n_100),
.B1(n_98),
.B2(n_83),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_127),
.A2(n_77),
.B1(n_54),
.B2(n_49),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_232),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_129),
.B(n_75),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_235),
.B(n_172),
.C(n_173),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_157),
.B(n_32),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_236),
.B(n_237),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_144),
.B(n_32),
.Y(n_237)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_155),
.B(n_33),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_239),
.B(n_244),
.Y(n_329)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_241),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_152),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_144),
.B(n_44),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_44),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_245),
.B(n_262),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_181),
.A2(n_73),
.B1(n_64),
.B2(n_54),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_252),
.B1(n_229),
.B2(n_224),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_190),
.Y(n_249)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_142),
.Y(n_254)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_151),
.Y(n_255)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

INVx11_ASAP7_75t_L g257 ( 
.A(n_143),
.Y(n_257)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

OR2x4_ASAP7_75t_L g258 ( 
.A(n_149),
.B(n_22),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_192),
.Y(n_259)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_166),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_143),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_264),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_198),
.B(n_22),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_171),
.A2(n_21),
.B1(n_47),
.B2(n_45),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_29),
.B1(n_227),
.B2(n_265),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_175),
.Y(n_264)
);

CKINVDCx9p33_ASAP7_75t_R g265 ( 
.A(n_175),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_265),
.Y(n_318)
);

CKINVDCx12_ASAP7_75t_R g266 ( 
.A(n_136),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_266),
.Y(n_322)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_269),
.Y(n_296)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_147),
.Y(n_268)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_128),
.B(n_69),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_154),
.A2(n_185),
.B1(n_174),
.B2(n_164),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_167),
.Y(n_272)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_131),
.Y(n_273)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_206),
.B(n_49),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_277),
.B(n_323),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_279),
.A2(n_280),
.B1(n_300),
.B2(n_208),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_246),
.A2(n_148),
.B1(n_173),
.B2(n_187),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_209),
.B(n_142),
.CI(n_33),
.CON(n_281),
.SN(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_324),
.B(n_258),
.C(n_269),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_219),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_289),
.B(n_320),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_311),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_241),
.A2(n_163),
.B1(n_126),
.B2(n_43),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_252),
.A2(n_195),
.B1(n_187),
.B2(n_146),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_209),
.A2(n_43),
.B(n_130),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_306),
.A2(n_230),
.B(n_240),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_220),
.B(n_195),
.C(n_153),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_271),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_242),
.A2(n_161),
.B1(n_165),
.B2(n_137),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_235),
.A2(n_165),
.B1(n_162),
.B2(n_141),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_235),
.A2(n_162),
.B1(n_141),
.B2(n_138),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_328),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_138),
.Y(n_323)
);

AOI32xp33_ASAP7_75t_L g324 ( 
.A1(n_225),
.A2(n_137),
.A3(n_133),
.B1(n_5),
.B2(n_6),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_247),
.Y(n_327)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_208),
.A2(n_133),
.B1(n_3),
.B2(n_6),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_330),
.B(n_346),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_285),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_339),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_333),
.A2(n_338),
.B1(n_356),
.B2(n_299),
.Y(n_380)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_282),
.Y(n_335)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_257),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_340),
.Y(n_389)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_291),
.Y(n_342)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_342),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_343),
.B(n_316),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_213),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_348),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_276),
.A2(n_204),
.B(n_218),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_345),
.A2(n_288),
.B(n_312),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_207),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_283),
.B(n_249),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_215),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_352),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_259),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_359),
.Y(n_398)
);

INVx13_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_250),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_275),
.Y(n_353)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_317),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_357),
.Y(n_395)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_355),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_279),
.A2(n_231),
.B1(n_248),
.B2(n_223),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_318),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_292),
.B(n_254),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_366),
.Y(n_405)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_364),
.Y(n_376)
);

INVx13_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g363 ( 
.A(n_284),
.B(n_210),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_363),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_278),
.B(n_234),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_277),
.B(n_217),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_368),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_226),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_296),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_369),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_302),
.B(n_281),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_370),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_278),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_371),
.A2(n_299),
.B1(n_328),
.B2(n_281),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_347),
.C(n_341),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_381),
.C(n_390),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_333),
.A2(n_290),
.B1(n_321),
.B2(n_320),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_374),
.A2(n_380),
.B1(n_407),
.B2(n_376),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_341),
.B(n_278),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_379),
.B(n_388),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_308),
.C(n_289),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_361),
.A2(n_300),
.B1(n_280),
.B2(n_306),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_383),
.A2(n_396),
.B1(n_404),
.B2(n_367),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

FAx1_ASAP7_75t_SL g387 ( 
.A(n_365),
.B(n_319),
.CI(n_310),
.CON(n_387),
.SN(n_387)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_392),
.Y(n_416)
);

AND2x2_ASAP7_75t_SL g388 ( 
.A(n_343),
.B(n_309),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_361),
.A2(n_316),
.B1(n_313),
.B2(n_304),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_350),
.C(n_345),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_368),
.Y(n_438)
);

FAx1_ASAP7_75t_L g403 ( 
.A(n_330),
.B(n_307),
.CI(n_293),
.CON(n_403),
.SN(n_403)
);

AO22x2_ASAP7_75t_L g420 ( 
.A1(n_403),
.A2(n_363),
.B1(n_339),
.B2(n_360),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_274),
.B1(n_293),
.B2(n_305),
.Y(n_404)
);

BUFx12_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_408),
.Y(n_442)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_398),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_424),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_398),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_426),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_414),
.A2(n_407),
.B1(n_392),
.B2(n_403),
.Y(n_444)
);

OAI21xp33_ASAP7_75t_L g415 ( 
.A1(n_394),
.A2(n_369),
.B(n_364),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_415),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_332),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_417),
.B(n_418),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_357),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_402),
.Y(n_419)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_419),
.Y(n_447)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_420),
.Y(n_460)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_402),
.Y(n_421)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_421),
.Y(n_461)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_346),
.Y(n_423)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_354),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_389),
.Y(n_425)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_425),
.Y(n_469)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_401),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_431),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_405),
.B(n_334),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_429),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_387),
.B(n_355),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_331),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_430),
.A2(n_377),
.B(n_376),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_383),
.A2(n_331),
.B1(n_338),
.B2(n_356),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_406),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_433),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_377),
.A2(n_331),
.B1(n_367),
.B2(n_363),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_435),
.Y(n_459)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_382),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_387),
.B(n_334),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_436),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_374),
.A2(n_364),
.B1(n_336),
.B2(n_353),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_437),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_390),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_340),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_373),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_444),
.A2(n_446),
.B1(n_455),
.B2(n_458),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_445),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_414),
.A2(n_372),
.B1(n_381),
.B2(n_404),
.Y(n_446)
);

NOR2x1_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_376),
.Y(n_451)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

NAND2x1_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_382),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_408),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_410),
.A2(n_432),
.B1(n_416),
.B2(n_413),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_410),
.A2(n_375),
.B1(n_397),
.B2(n_379),
.Y(n_458)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_463),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_440),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_409),
.B(n_393),
.Y(n_465)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_465),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_420),
.A2(n_430),
.B1(n_431),
.B2(n_411),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_466),
.A2(n_400),
.B1(n_408),
.B2(n_336),
.Y(n_492)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_470),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_454),
.B(n_438),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_471),
.B(n_481),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_468),
.A2(n_411),
.B(n_420),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_472),
.A2(n_483),
.B(n_469),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_473),
.B(n_461),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_L g474 ( 
.A1(n_445),
.A2(n_420),
.B(n_434),
.C(n_419),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_479),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_388),
.C(n_440),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_480),
.C(n_482),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_312),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_388),
.C(n_435),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_335),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_427),
.C(n_426),
.Y(n_482)
);

XOR2x2_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_425),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_443),
.A2(n_421),
.B1(n_422),
.B2(n_375),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_484),
.A2(n_489),
.B1(n_495),
.B2(n_485),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_441),
.Y(n_485)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_399),
.C(n_400),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_442),
.C(n_452),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_449),
.B(n_351),
.Y(n_488)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_465),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_399),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_493),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_492),
.A2(n_456),
.B1(n_442),
.B2(n_459),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_453),
.B(n_351),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_448),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_457),
.A2(n_305),
.B1(n_274),
.B2(n_342),
.Y(n_495)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_496),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_483),
.A2(n_444),
.B1(n_457),
.B2(n_456),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_505),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_511),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_477),
.A2(n_459),
.B1(n_460),
.B2(n_467),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_491),
.A2(n_467),
.B1(n_463),
.B2(n_460),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_516),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_507),
.B(n_508),
.C(n_490),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_452),
.C(n_448),
.Y(n_508)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_509),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_486),
.A2(n_469),
.B1(n_462),
.B2(n_461),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_451),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_515),
.Y(n_530)
);

FAx1_ASAP7_75t_SL g513 ( 
.A(n_475),
.B(n_451),
.CI(n_462),
.CON(n_513),
.SN(n_513)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_513),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_514),
.A2(n_470),
.B(n_447),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_482),
.A2(n_447),
.B1(n_359),
.B2(n_337),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_510),
.B(n_478),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_518),
.B(n_526),
.Y(n_534)
);

BUFx12_ASAP7_75t_L g522 ( 
.A(n_513),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_523),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_511),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_504),
.Y(n_525)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_525),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_503),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_527),
.A2(n_531),
.B(n_532),
.Y(n_541)
);

AOI221xp5_ASAP7_75t_L g529 ( 
.A1(n_508),
.A2(n_476),
.B1(n_495),
.B2(n_491),
.C(n_474),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_529),
.B(n_498),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_501),
.A2(n_493),
.B(n_492),
.Y(n_531)
);

INVx13_ASAP7_75t_L g532 ( 
.A(n_502),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_509),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_519),
.A2(n_500),
.B1(n_507),
.B2(n_515),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_535),
.B(n_537),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_517),
.B(n_501),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_547),
.Y(n_553)
);

XNOR2x1_ASAP7_75t_L g557 ( 
.A(n_539),
.B(n_545),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_512),
.C(n_516),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_542),
.C(n_544),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_528),
.A2(n_505),
.B1(n_473),
.B2(n_497),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_528),
.A2(n_497),
.B1(n_286),
.B2(n_315),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_530),
.B(n_362),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_521),
.C(n_524),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_546),
.B(n_534),
.C(n_304),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_533),
.B(n_286),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_540),
.B(n_521),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_548),
.B(n_551),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_520),
.C(n_522),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_550),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_522),
.C(n_532),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_543),
.B(n_362),
.Y(n_551)
);

INVx11_ASAP7_75t_L g552 ( 
.A(n_539),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_552),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_315),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_551),
.Y(n_565)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_556),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_554),
.C(n_550),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_561),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_549),
.A2(n_232),
.B1(n_303),
.B2(n_216),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_565),
.B(n_566),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_303),
.C(n_256),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_562),
.B(n_558),
.Y(n_567)
);

AO21x1_ASAP7_75t_L g574 ( 
.A1(n_567),
.A2(n_572),
.B(n_566),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_563),
.C(n_560),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_568),
.B(n_570),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_564),
.B(n_553),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_561),
.B(n_536),
.Y(n_572)
);

AOI322xp5_ASAP7_75t_L g576 ( 
.A1(n_574),
.A2(n_569),
.A3(n_571),
.B1(n_557),
.B2(n_267),
.C1(n_212),
.C2(n_205),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_567),
.A2(n_557),
.B(n_267),
.Y(n_575)
);

A2O1A1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_575),
.A2(n_1),
.B(n_3),
.C(n_7),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_576),
.B(n_577),
.C(n_573),
.Y(n_578)
);

FAx1_ASAP7_75t_SL g579 ( 
.A(n_578),
.B(n_238),
.CI(n_233),
.CON(n_579),
.SN(n_579)
);

MAJx2_ASAP7_75t_L g580 ( 
.A(n_579),
.B(n_233),
.C(n_8),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_580),
.A2(n_579),
.B(n_9),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_581),
.B(n_9),
.Y(n_582)
);


endmodule