module fake_jpeg_25802_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_16),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_32),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_16),
.B1(n_32),
.B2(n_20),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_56),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_32),
.B1(n_20),
.B2(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_34),
.B1(n_33),
.B2(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_20),
.B1(n_29),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_25),
.B1(n_29),
.B2(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_41),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_77),
.B(n_92),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_65),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_67),
.B(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_19),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_78),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_51),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_75),
.C(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_80),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_30),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_28),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_39),
.CI(n_41),
.CON(n_83),
.SN(n_83)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_97),
.A3(n_34),
.B1(n_33),
.B2(n_24),
.Y(n_130)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_57),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_90),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_113)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_96),
.B(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_48),
.A2(n_26),
.B(n_35),
.C(n_22),
.D(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_28),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_54),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_53),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_56),
.B(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_104),
.B1(n_50),
.B2(n_27),
.Y(n_119)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_26),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_75),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_50),
.B1(n_58),
.B2(n_54),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_115),
.B1(n_121),
.B2(n_126),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_63),
.A2(n_50),
.B1(n_47),
.B2(n_61),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_31),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_50),
.B1(n_27),
.B2(n_31),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_50),
.B1(n_27),
.B2(n_31),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_26),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_132),
.B1(n_94),
.B2(n_91),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_35),
.B1(n_24),
.B2(n_23),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_35),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_141),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_73),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_64),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_64),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_152),
.B1(n_121),
.B2(n_131),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_84),
.B1(n_83),
.B2(n_90),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_73),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_163),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_83),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_129),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_84),
.B(n_90),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_162),
.B(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_77),
.Y(n_161)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_66),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_122),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_114),
.B(n_122),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_170),
.B(n_189),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_124),
.B(n_126),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_172),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_130),
.B1(n_124),
.B2(n_78),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_181),
.B1(n_185),
.B2(n_192),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_128),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_179),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_146),
.B1(n_152),
.B2(n_155),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_184),
.B1(n_187),
.B2(n_193),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_0),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_85),
.B1(n_87),
.B2(n_79),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_89),
.B1(n_95),
.B2(n_66),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_99),
.B1(n_88),
.B2(n_104),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_129),
.B1(n_88),
.B2(n_106),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_106),
.B(n_127),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_127),
.B(n_118),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_24),
.B(n_1),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_144),
.A2(n_110),
.B1(n_134),
.B2(n_100),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_156),
.B1(n_164),
.B2(n_142),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_166),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_201),
.B1(n_218),
.B2(n_221),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_163),
.B1(n_110),
.B2(n_143),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_203),
.B1(n_204),
.B2(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_166),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_149),
.C(n_148),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_211),
.C(n_222),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_118),
.B1(n_134),
.B2(n_149),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_91),
.B1(n_153),
.B2(n_70),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_9),
.C(n_14),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_177),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_213),
.B1(n_220),
.B2(n_223),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_172),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_170),
.A2(n_3),
.B(n_4),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_189),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_192),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_194),
.B1(n_180),
.B2(n_196),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_187),
.B1(n_191),
.B2(n_182),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_7),
.C(n_13),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_15),
.B1(n_7),
.B2(n_11),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_173),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_227),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_173),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_168),
.C(n_171),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_233),
.C(n_244),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_171),
.C(n_178),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_208),
.A2(n_196),
.B1(n_183),
.B2(n_169),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_236),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_193),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_190),
.B1(n_195),
.B2(n_174),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_199),
.Y(n_248)
);

XOR2x2_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_201),
.Y(n_241)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_242),
.CI(n_213),
.CON(n_253),
.SN(n_253)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_203),
.B(n_195),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_11),
.C(n_15),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_197),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_248),
.A2(n_261),
.B1(n_263),
.B2(n_250),
.Y(n_277)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_199),
.C(n_216),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_251),
.C(n_258),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_209),
.C(n_211),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_260),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_222),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_257),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_204),
.C(n_206),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_214),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_241),
.B(n_242),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_270),
.B(n_254),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_237),
.B1(n_238),
.B2(n_226),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_272),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_212),
.B1(n_225),
.B2(n_5),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_278),
.B1(n_253),
.B2(n_251),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_225),
.B(n_212),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_246),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_3),
.B1(n_6),
.B2(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_262),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_246),
.C(n_258),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_276),
.C(n_271),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_257),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_286),
.A2(n_288),
.B(n_270),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_278),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_290),
.B(n_294),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_287),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_275),
.B(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_267),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_284),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_284),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_291),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_SL g306 ( 
.A(n_304),
.B(n_298),
.C(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_293),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_306),
.Y(n_307)
);

AOI221xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_302),
.B1(n_292),
.B2(n_266),
.C(n_272),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_6),
.B1(n_254),
.B2(n_304),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_6),
.Y(n_311)
);


endmodule