module fake_jpeg_18656_n_410 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_49),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_53),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_69),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_63),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_68),
.Y(n_75)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_70),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_29),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_13),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_35),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_36),
.B1(n_32),
.B2(n_34),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_77),
.B1(n_93),
.B2(n_97),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_32),
.B1(n_19),
.B2(n_33),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_43),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_71),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_98),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_32),
.B1(n_19),
.B2(n_33),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_24),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_24),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_101),
.A2(n_60),
.B1(n_56),
.B2(n_16),
.Y(n_152)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_30),
.C(n_24),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_31),
.B1(n_28),
.B2(n_37),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_109),
.B1(n_111),
.B2(n_66),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_46),
.A2(n_37),
.B1(n_17),
.B2(n_27),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_61),
.A2(n_26),
.B1(n_19),
.B2(n_33),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_37),
.B1(n_27),
.B2(n_17),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_17),
.B1(n_27),
.B2(n_26),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_51),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_131),
.Y(n_160)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_118),
.B(n_134),
.Y(n_166)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_121),
.Y(n_171)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_26),
.B1(n_15),
.B2(n_24),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_35),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_140),
.CI(n_101),
.CON(n_156),
.SN(n_156)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_16),
.B1(n_53),
.B2(n_60),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_124),
.A2(n_80),
.B1(n_92),
.B2(n_72),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_58),
.B1(n_55),
.B2(n_44),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_125),
.A2(n_148),
.B1(n_85),
.B2(n_80),
.Y(n_175)
);

OR2x2_ASAP7_75t_SL g128 ( 
.A(n_84),
.B(n_108),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_152),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_42),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_15),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_146),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_96),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_137),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_30),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_30),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_143),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_75),
.B(n_15),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_53),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_110),
.B1(n_91),
.B2(n_78),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_100),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_30),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_77),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_95),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_102),
.B(n_101),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_92),
.C(n_30),
.Y(n_173)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_161),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_56),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_164),
.B(n_165),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_75),
.C(n_91),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_75),
.B(n_88),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_173),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_95),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_189),
.B(n_152),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_175),
.A2(n_178),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_136),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_147),
.B1(n_132),
.B2(n_149),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_110),
.B(n_72),
.C(n_88),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_191),
.B(n_2),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_181),
.B1(n_193),
.B2(n_125),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_135),
.A2(n_112),
.B1(n_83),
.B2(n_35),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_131),
.B(n_116),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_124),
.C(n_146),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_112),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_115),
.A2(n_16),
.B(n_1),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_115),
.B1(n_113),
.B2(n_142),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_113),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_203),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_142),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_197),
.B(n_201),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_142),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_199),
.B(n_225),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_118),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_200),
.B(n_211),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_166),
.B(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_153),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_232),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_205),
.A2(n_213),
.B1(n_214),
.B2(n_224),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_117),
.B(n_119),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_206),
.A2(n_216),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_120),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_221),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_130),
.B1(n_145),
.B2(n_154),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_124),
.B1(n_133),
.B2(n_121),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_127),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_222),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_155),
.B(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_156),
.B(n_124),
.C(n_139),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_231),
.C(n_157),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_163),
.B(n_0),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_181),
.B1(n_180),
.B2(n_222),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_185),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_156),
.B(n_5),
.C(n_6),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_160),
.B(n_5),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_158),
.B(n_172),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_240),
.B(n_256),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_170),
.B(n_158),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_218),
.B1(n_213),
.B2(n_203),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_247),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_157),
.B1(n_189),
.B2(n_184),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_244),
.A2(n_258),
.B1(n_220),
.B2(n_204),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_196),
.B(n_161),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_173),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_251),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_157),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_195),
.B(n_159),
.C(n_184),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_261),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_159),
.B(n_174),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_202),
.B1(n_205),
.B2(n_189),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_199),
.A2(n_178),
.B(n_174),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_201),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_264),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_197),
.B(n_179),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_206),
.A2(n_175),
.B(n_187),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_199),
.B(n_210),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_209),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_280),
.Y(n_300)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_316)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_277),
.B1(n_279),
.B2(n_282),
.Y(n_304)
);

BUFx12f_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_278),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_258),
.A2(n_214),
.B1(n_229),
.B2(n_232),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_254),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_233),
.A2(n_230),
.B1(n_194),
.B2(n_210),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_281),
.A2(n_256),
.B1(n_233),
.B2(n_252),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_241),
.A2(n_259),
.B1(n_240),
.B2(n_267),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_231),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_286),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_228),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_221),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_290),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_234),
.B(n_169),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_288),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_169),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_239),
.B(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_244),
.A2(n_224),
.B1(n_187),
.B2(n_217),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_208),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_235),
.B(n_162),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_236),
.A2(n_207),
.B1(n_226),
.B2(n_162),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_273),
.B(n_247),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_309),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_250),
.C(n_237),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_306),
.C(n_314),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_237),
.C(n_242),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_308),
.A2(n_310),
.B1(n_279),
.B2(n_295),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_251),
.C(n_248),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_293),
.A2(n_266),
.B1(n_248),
.B2(n_249),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_249),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_312),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_266),
.Y(n_312)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_168),
.C(n_238),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_168),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_322),
.C(n_278),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_319),
.A2(n_290),
.B1(n_291),
.B2(n_271),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_6),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_329),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_286),
.Y(n_327)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_314),
.A2(n_296),
.B1(n_282),
.B2(n_270),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_328),
.A2(n_334),
.B1(n_341),
.B2(n_318),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_284),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_305),
.A2(n_281),
.B1(n_295),
.B2(n_287),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_330),
.A2(n_331),
.B1(n_337),
.B2(n_340),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_269),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_335),
.Y(n_354)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_305),
.A2(n_296),
.B1(n_283),
.B2(n_278),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_278),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_343),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_299),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_304),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_340)
);

NOR2x1_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_7),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_342),
.A2(n_303),
.B(n_319),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_304),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

BUFx12_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_347),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_349),
.A2(n_351),
.B(n_10),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_302),
.C(n_306),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_350),
.B(n_325),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_SL g351 ( 
.A1(n_334),
.A2(n_310),
.B(n_317),
.C(n_309),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_356),
.Y(n_364)
);

BUFx12_ASAP7_75t_L g355 ( 
.A(n_341),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_355),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_339),
.Y(n_356)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_308),
.B(n_322),
.Y(n_358)
);

AOI31xp33_ASAP7_75t_L g363 ( 
.A1(n_358),
.A2(n_323),
.A3(n_312),
.B(n_325),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_311),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_360),
.B(n_336),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_353),
.A2(n_342),
.B1(n_323),
.B2(n_337),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_365),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_371),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_373),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_336),
.Y(n_370)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_370),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_9),
.C(n_10),
.Y(n_371)
);

XOR2x2_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_9),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_372),
.A2(n_374),
.B(n_373),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_9),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_374),
.A2(n_355),
.B(n_359),
.Y(n_380)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_377),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_355),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_381),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_380),
.A2(n_351),
.B(n_347),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_370),
.B(n_348),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_345),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_385),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_350),
.C(n_356),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_364),
.C(n_369),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_347),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_383),
.A2(n_362),
.B(n_368),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_388),
.B(n_390),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_379),
.A2(n_368),
.B(n_372),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_365),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_391),
.B(n_394),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_384),
.C(n_376),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_379),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_351),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g404 ( 
.A(n_395),
.B(n_397),
.CI(n_11),
.CON(n_404),
.SN(n_404)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_396),
.B(n_400),
.C(n_389),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_392),
.A2(n_371),
.B(n_11),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_11),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_401),
.B(n_403),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_402),
.B(n_404),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_386),
.C(n_393),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_398),
.C(n_404),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_405),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_408),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_11),
.Y(n_410)
);


endmodule