module real_jpeg_29269_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_314, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_314;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_0),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_0),
.A2(n_30),
.B1(n_55),
.B2(n_56),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_0),
.A2(n_30),
.B1(n_62),
.B2(n_63),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_1),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_1),
.A2(n_46),
.B1(n_62),
.B2(n_63),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_62),
.Y(n_93)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_2),
.Y(n_96)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_3),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_153),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_153),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_153),
.Y(n_246)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_5),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_160),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_160),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_160),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_6),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_8),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_102),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_102),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_102),
.Y(n_241)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_10),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_136),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_136),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_136),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_11),
.A2(n_40),
.B1(n_55),
.B2(n_56),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_61)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_15),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_SL g165 ( 
.A1(n_15),
.A2(n_33),
.B(n_37),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_15),
.B(n_35),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_15),
.A2(n_55),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_15),
.B(n_55),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_15),
.B(n_59),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_15),
.A2(n_92),
.B1(n_96),
.B2(n_252),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_15),
.A2(n_36),
.B(n_268),
.Y(n_267)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_16),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_17),
.A2(n_55),
.B1(n_56),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_17),
.A2(n_62),
.B1(n_63),
.B2(n_71),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_17),
.A2(n_36),
.B1(n_37),
.B2(n_71),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_103),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_75),
.C(n_81),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_23),
.B(n_75),
.CI(n_81),
.CON(n_137),
.SN(n_137)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_74),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_24),
.A2(n_25),
.B1(n_105),
.B2(n_113),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_25),
.B(n_43),
.C(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_39),
.B2(n_41),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_26),
.A2(n_31),
.B1(n_41),
.B2(n_100),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_33),
.Y(n_34)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_28),
.A2(n_38),
.B(n_164),
.C(n_165),
.Y(n_163)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_31),
.A2(n_41),
.B1(n_158),
.B2(n_161),
.Y(n_157)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_32),
.A2(n_35),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_32),
.A2(n_35),
.B1(n_101),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_32),
.A2(n_35),
.B1(n_135),
.B2(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_32),
.A2(n_35),
.B1(n_159),
.B2(n_196),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_49),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_36),
.A2(n_53),
.A3(n_56),
.B1(n_269),
.B2(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_37),
.B(n_164),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_60),
.B1(n_72),
.B2(n_73),
.Y(n_42)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_57),
.B2(n_59),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_48),
.B1(n_52),
.B2(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_47),
.A2(n_57),
.B1(n_59),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_47),
.A2(n_59),
.B1(n_78),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_47),
.A2(n_59),
.B1(n_127),
.B2(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_47),
.A2(n_59),
.B1(n_190),
.B2(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_48),
.A2(n_52),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_48),
.A2(n_52),
.B1(n_169),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_48),
.A2(n_52),
.B1(n_202),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_53),
.Y(n_278)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_56),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g229 ( 
.A1(n_55),
.A2(n_63),
.A3(n_69),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_55),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_60),
.A2(n_73),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_67),
.B(n_70),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_67),
.B1(n_70),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_61),
.A2(n_67),
.B1(n_87),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_61),
.A2(n_67),
.B1(n_133),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_61),
.A2(n_67),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_61),
.A2(n_67),
.B1(n_227),
.B2(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_61),
.B(n_164),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_61),
.A2(n_67),
.B1(n_194),
.B2(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_62),
.B(n_66),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_62),
.B(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_76),
.B(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_98),
.B(n_99),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_83),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_84),
.A2(n_85),
.B1(n_91),
.B2(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_88),
.A2(n_90),
.B1(n_149),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_88),
.A2(n_90),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_98),
.B1(n_99),
.B2(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B(n_97),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_97),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_92),
.A2(n_130),
.B1(n_131),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_92),
.A2(n_94),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_92),
.A2(n_96),
.B1(n_246),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_92),
.A2(n_94),
.B1(n_241),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_93),
.A2(n_95),
.B1(n_146),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_93),
.A2(n_95),
.B1(n_167),
.B2(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_93),
.A2(n_95),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

INVx5_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_99),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_110),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_138),
.B(n_310),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_137),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_118),
.B(n_137),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_124),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_123),
.Y(n_181)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_124),
.A2(n_125),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.C(n_134),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_126),
.B(n_128),
.CI(n_134),
.CON(n_175),
.SN(n_175)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_132),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_137),
.Y(n_312)
);

AOI321xp33_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_177),
.A3(n_182),
.B1(n_304),
.B2(n_309),
.C(n_314),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_140),
.A2(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_172),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_141),
.B(n_172),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_156),
.C(n_171),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_142),
.B(n_171),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_151),
.C(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_147),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_162),
.C(n_168),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_168),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_162),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_166),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_164),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_175),
.C(n_176),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_175),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_178),
.B(n_179),
.Y(n_309)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_212),
.C(n_217),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_206),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_184),
.B(n_206),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_197),
.C(n_198),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_185),
.B(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_195),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_192),
.C(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_197),
.Y(n_302)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_200),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_203),
.B(n_205),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_204),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_209),
.C(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_213),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_214),
.B(n_215),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_298),
.B(n_303),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_284),
.B(n_297),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_262),
.B(n_283),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_242),
.B(n_261),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_232),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_222),
.B(n_232),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_237),
.C(n_239),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_240),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_249),
.B(n_260),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_248),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_254),
.B(n_259),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_264),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_275),
.B1(n_281),
.B2(n_282),
.Y(n_264)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_265)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_274),
.C(n_282),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_272),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_275),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_279),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_293),
.C(n_295),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);


endmodule