module fake_jpeg_11735_n_109 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_35),
.B1(n_41),
.B2(n_3),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_45),
.B1(n_44),
.B2(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_60),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_7),
.B(n_8),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_3),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_5),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_68),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_18),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_6),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_20),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_12),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_86),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_88),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_90),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_15),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_21),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_68),
.B(n_78),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_82),
.C(n_89),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_78),
.B1(n_23),
.B2(n_25),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_89),
.B1(n_83),
.B2(n_34),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_81),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_93),
.B1(n_97),
.B2(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_104),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_26),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_108),
.Y(n_109)
);


endmodule