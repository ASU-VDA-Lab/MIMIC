module fake_jpeg_30734_n_500 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_500);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_500;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_19),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_93),
.Y(n_105)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_90),
.Y(n_113)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_1),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_75),
.B(n_96),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_94),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_30),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_43),
.B1(n_39),
.B2(n_47),
.Y(n_115)
);

CKINVDCx6p67_ASAP7_75t_R g96 ( 
.A(n_39),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_98),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_33),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_26),
.B1(n_46),
.B2(n_42),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_101),
.B(n_145),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_52),
.A2(n_67),
.B1(n_58),
.B2(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_102),
.A2(n_111),
.B1(n_120),
.B2(n_151),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_87),
.B1(n_54),
.B2(n_64),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_107),
.A2(n_132),
.B1(n_136),
.B2(n_144),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_47),
.B1(n_43),
.B2(n_41),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_115),
.A2(n_14),
.B1(n_5),
.B2(n_7),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_43),
.B1(n_49),
.B2(n_17),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_82),
.A2(n_46),
.B1(n_42),
.B2(n_37),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_90),
.B1(n_96),
.B2(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_75),
.B(n_37),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_1),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_93),
.B1(n_95),
.B2(n_39),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_35),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_35),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_80),
.A2(n_49),
.B1(n_16),
.B2(n_17),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_80),
.A2(n_39),
.B1(n_44),
.B2(n_16),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_155),
.B1(n_34),
.B2(n_32),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_80),
.A2(n_44),
.B1(n_38),
.B2(n_28),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_164),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_38),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_160),
.B(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_161),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_28),
.C(n_34),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_162),
.B(n_168),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_48),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_166),
.A2(n_170),
.B1(n_180),
.B2(n_194),
.Y(n_223)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_109),
.B(n_48),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_32),
.A3(n_30),
.B1(n_48),
.B2(n_18),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_173),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_18),
.B1(n_30),
.B2(n_48),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_171),
.A2(n_188),
.B1(n_199),
.B2(n_141),
.Y(n_233)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_117),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g240 ( 
.A(n_174),
.B(n_114),
.Y(n_240)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_176),
.B(n_181),
.Y(n_242)
);

BUFx4f_ASAP7_75t_SL g177 ( 
.A(n_116),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_100),
.A2(n_30),
.B1(n_3),
.B2(n_4),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_138),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_184),
.B(n_186),
.Y(n_243)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_2),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_108),
.Y(n_187)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_110),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_193),
.Y(n_244)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_5),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_120),
.B1(n_111),
.B2(n_102),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_112),
.B(n_8),
.C(n_9),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_200),
.Y(n_208)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_135),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_100),
.B(n_9),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_154),
.B(n_10),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_SL g248 ( 
.A(n_202),
.B(n_10),
.C(n_11),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_104),
.B1(n_128),
.B2(n_134),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_210),
.A2(n_237),
.B1(n_247),
.B2(n_126),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_246),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_160),
.A2(n_104),
.B1(n_128),
.B2(n_134),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_230),
.A2(n_201),
.B1(n_175),
.B2(n_178),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_165),
.B(n_174),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_157),
.A2(n_166),
.B1(n_196),
.B2(n_169),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_140),
.B1(n_118),
.B2(n_122),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

AO21x2_ASAP7_75t_L g245 ( 
.A1(n_188),
.A2(n_157),
.B(n_177),
.Y(n_245)
);

AOI22x1_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_188),
.B1(n_205),
.B2(n_165),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_173),
.A2(n_103),
.B1(n_123),
.B2(n_122),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_158),
.A2(n_118),
.B1(n_123),
.B2(n_126),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_202),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_250),
.B(n_263),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_158),
.B(n_164),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_251),
.A2(n_255),
.B(n_279),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_162),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_252),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_158),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_259),
.Y(n_291)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_202),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_187),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_163),
.C(n_168),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_231),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_211),
.B(n_163),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_280),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_262),
.A2(n_272),
.B1(n_276),
.B2(n_277),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_224),
.B(n_168),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_227),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_265),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_170),
.B1(n_185),
.B2(n_191),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_281),
.B1(n_245),
.B2(n_240),
.Y(n_288)
);

NOR3xp33_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_197),
.C(n_188),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_183),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_182),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_223),
.A2(n_195),
.B1(n_192),
.B2(n_172),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_223),
.A2(n_177),
.B1(n_167),
.B2(n_14),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_11),
.B(n_13),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_213),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_245),
.A2(n_234),
.B1(n_239),
.B2(n_247),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_228),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_287),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_239),
.B1(n_219),
.B2(n_230),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_286),
.Y(n_304)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_214),
.Y(n_285)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_288),
.A2(n_254),
.B1(n_284),
.B2(n_264),
.Y(n_335)
);

OAI32xp33_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_245),
.A3(n_231),
.B1(n_228),
.B2(n_222),
.Y(n_289)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_279),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_305),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_249),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_298),
.C(n_260),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_236),
.Y(n_351)
);

BUFx24_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_226),
.B1(n_218),
.B2(n_209),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_287),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_SL g303 ( 
.A1(n_269),
.A2(n_209),
.B(n_218),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_303),
.A2(n_321),
.B1(n_272),
.B2(n_276),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_285),
.Y(n_305)
);

AO21x2_ASAP7_75t_L g307 ( 
.A1(n_250),
.A2(n_226),
.B(n_214),
.Y(n_307)
);

AOI22x1_ASAP7_75t_L g331 ( 
.A1(n_307),
.A2(n_250),
.B1(n_281),
.B2(n_277),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_273),
.A2(n_229),
.B(n_221),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_258),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_278),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_274),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_316),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_270),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_319),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_254),
.A2(n_216),
.B1(n_221),
.B2(n_235),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_273),
.A2(n_229),
.B(n_216),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_312),
.Y(n_326)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_296),
.B(n_263),
.CI(n_251),
.CON(n_327),
.SN(n_327)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_328),
.Y(n_366)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_329),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_330),
.B(n_351),
.Y(n_376)
);

AOI22x1_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_307),
.B1(n_304),
.B2(n_315),
.Y(n_362)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_339),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_334),
.A2(n_338),
.B1(n_310),
.B2(n_304),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_335),
.A2(n_294),
.B1(n_307),
.B2(n_293),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_255),
.C(n_256),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_292),
.C(n_322),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_310),
.A2(n_262),
.B1(n_271),
.B2(n_275),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_341),
.A2(n_300),
.B(n_323),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_345),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_311),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_348),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_286),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_299),
.Y(n_348)
);

OAI32xp33_ASAP7_75t_SL g349 ( 
.A1(n_315),
.A2(n_235),
.A3(n_236),
.B1(n_302),
.B2(n_289),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_302),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_299),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_352),
.B(n_290),
.Y(n_370)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_354),
.Y(n_377)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_309),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_309),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_318),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_359),
.A2(n_363),
.B1(n_364),
.B2(n_381),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_347),
.A2(n_315),
.B(n_294),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_361),
.A2(n_375),
.B(n_350),
.Y(n_391)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_324),
.A2(n_307),
.B1(n_292),
.B2(n_296),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_351),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_369),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_368),
.A2(n_328),
.B1(n_329),
.B2(n_332),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_291),
.Y(n_369)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_313),
.C(n_301),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_371),
.B(n_349),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_335),
.Y(n_402)
);

INVx3_ASAP7_75t_SL g373 ( 
.A(n_336),
.Y(n_373)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_308),
.C(n_306),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_380),
.C(n_350),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_324),
.A2(n_334),
.B1(n_346),
.B2(n_336),
.Y(n_378)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_342),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_384),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_290),
.C(n_323),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_343),
.A2(n_307),
.B1(n_316),
.B2(n_305),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_345),
.Y(n_384)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_SL g389 ( 
.A(n_376),
.B(n_299),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_389),
.B(n_397),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_391),
.A2(n_406),
.B(n_361),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_357),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_395),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_357),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_396),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_365),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_399),
.B(n_402),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_400),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_405),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_376),
.B(n_349),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_SL g406 ( 
.A(n_372),
.B(n_341),
.C(n_331),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_374),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_409),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_331),
.C(n_355),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_408),
.B(n_363),
.C(n_368),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_364),
.A2(n_341),
.B1(n_325),
.B2(n_326),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_377),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_411),
.A2(n_381),
.B1(n_393),
.B2(n_387),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_416),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_425),
.Y(n_435)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_392),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_401),
.A2(n_356),
.B1(n_362),
.B2(n_375),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_428),
.Y(n_445)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_424),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_371),
.C(n_377),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_360),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_431),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_387),
.A2(n_406),
.B1(n_393),
.B2(n_402),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_396),
.Y(n_429)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_429),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_388),
.B(n_399),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_400),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_420),
.A2(n_403),
.B1(n_405),
.B2(n_404),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_419),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_449),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_414),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_436),
.B(n_440),
.Y(n_455)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_432),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_383),
.Y(n_443)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_443),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_413),
.A2(n_391),
.B1(n_392),
.B2(n_408),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_444),
.A2(n_415),
.B1(n_423),
.B2(n_425),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_416),
.A2(n_409),
.B(n_362),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_446),
.A2(n_427),
.B(n_382),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_366),
.Y(n_448)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_448),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_385),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_464),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_448),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_439),
.B(n_426),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_461),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_457),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_419),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_460),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_430),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_445),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_446),
.A2(n_412),
.B(n_431),
.Y(n_462)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_462),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_430),
.C(n_388),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_433),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_444),
.B(n_412),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_442),
.Y(n_466)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_445),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_472),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_447),
.C(n_448),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_474),
.B(n_476),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_358),
.Y(n_475)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_475),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_458),
.C(n_463),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_437),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_477),
.B(n_457),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_480),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_467),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_459),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_481),
.B(n_474),
.Y(n_487)
);

INVx11_ASAP7_75t_L g484 ( 
.A(n_475),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_484),
.B(n_465),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_471),
.A2(n_462),
.B(n_464),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_486),
.B(n_469),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_487),
.B(n_488),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_479),
.Y(n_488)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_490),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_491),
.A2(n_485),
.B(n_482),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_494),
.A2(n_489),
.B(n_478),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_495),
.A2(n_496),
.B(n_492),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_493),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_497),
.A2(n_481),
.B(n_483),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_498),
.B(n_339),
.C(n_468),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_318),
.Y(n_500)
);


endmodule