module fake_jpeg_6143_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_8),
.B(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_19),
.B1(n_13),
.B2(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_47),
.B1(n_19),
.B2(n_25),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_13),
.B1(n_19),
.B2(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_55),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_28),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_32),
.Y(n_58)
);

OA22x2_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_22),
.B1(n_34),
.B2(n_32),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_45),
.B1(n_24),
.B2(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_65),
.B(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_21),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_18),
.B(n_34),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_16),
.B1(n_25),
.B2(n_26),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_45),
.C(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_23),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_80),
.B1(n_23),
.B2(n_64),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_78),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_55),
.B1(n_59),
.B2(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_90),
.Y(n_101)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_83),
.B(n_76),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_69),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_94),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_68),
.C(n_24),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_56),
.B1(n_58),
.B2(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_65),
.B1(n_60),
.B2(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_71),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_17),
.B1(n_24),
.B2(n_18),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_68),
.A3(n_80),
.B1(n_24),
.B2(n_50),
.C1(n_18),
.C2(n_81),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_71),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_104),
.B(n_18),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_73),
.B(n_75),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_107),
.B(n_108),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_94),
.C(n_96),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

OAI322xp33_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_88),
.A3(n_97),
.B1(n_93),
.B2(n_90),
.C1(n_92),
.C2(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_116),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_99),
.B(n_100),
.C(n_102),
.D(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_115),
.B(n_116),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_12),
.A3(n_10),
.B1(n_7),
.B2(n_5),
.C1(n_2),
.C2(n_4),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_123),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_107),
.B1(n_104),
.B2(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_120),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_118),
.A2(n_121),
.B(n_114),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_128),
.B(n_125),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_113),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_120),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_134)
);

OAI31xp33_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_117),
.A3(n_12),
.B(n_7),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_133),
.B(n_5),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_3),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_136),
.B(n_5),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_6),
.Y(n_139)
);


endmodule