module fake_jpeg_18821_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_42),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_33),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_34),
.B1(n_25),
.B2(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_59),
.B1(n_23),
.B2(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_34),
.B1(n_25),
.B2(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_64),
.B(n_79),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_43),
.B1(n_41),
.B2(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_76),
.B1(n_86),
.B2(n_50),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_45),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_43),
.B1(n_41),
.B2(n_34),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_77),
.B1(n_78),
.B2(n_84),
.Y(n_111)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx4f_ASAP7_75t_SL g98 ( 
.A(n_73),
.Y(n_98)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_16),
.B1(n_54),
.B2(n_60),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_19),
.B1(n_44),
.B2(n_37),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_44),
.B1(n_27),
.B2(n_20),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_22),
.B1(n_30),
.B2(n_27),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_24),
.B1(n_30),
.B2(n_22),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_80),
.A2(n_82),
.B1(n_95),
.B2(n_50),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_24),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_24),
.B1(n_30),
.B2(n_22),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_83),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_40),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_17),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_38),
.B1(n_17),
.B2(n_31),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_93),
.Y(n_109)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_31),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_16),
.B(n_18),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_101),
.B(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_112),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_115),
.B1(n_119),
.B2(n_121),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_116),
.B1(n_124),
.B2(n_70),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_77),
.A2(n_69),
.B1(n_66),
.B2(n_50),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_13),
.B(n_10),
.Y(n_117)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_39),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_123),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_60),
.B1(n_38),
.B2(n_39),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_81),
.A2(n_32),
.B1(n_18),
.B2(n_40),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_21),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_32),
.B1(n_16),
.B2(n_36),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_29),
.B1(n_40),
.B2(n_36),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_21),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_36),
.C(n_73),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_127),
.B(n_128),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_74),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_153),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_100),
.B1(n_121),
.B2(n_119),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_137),
.B(n_145),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_110),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_113),
.B1(n_106),
.B2(n_126),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_74),
.C(n_26),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_141),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_72),
.Y(n_143)
);

OR2x6_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_105),
.B(n_87),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_146),
.B(n_148),
.Y(n_185)
);

OR2x4_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_26),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_106),
.B1(n_148),
.B2(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_73),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_65),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_155),
.B(n_154),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_96),
.C(n_101),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_163),
.C(n_29),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_157),
.A2(n_158),
.B1(n_177),
.B2(n_186),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_118),
.B1(n_116),
.B2(n_123),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_151),
.B1(n_89),
.B2(n_68),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_103),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_125),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_122),
.C(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_122),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_178),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_110),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_143),
.B(n_147),
.Y(n_176)
);

AO21x2_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_98),
.B(n_138),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_91),
.B1(n_95),
.B2(n_92),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_68),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_94),
.B1(n_106),
.B2(n_97),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_140),
.B1(n_89),
.B2(n_68),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_72),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_182),
.B(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_72),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_126),
.B1(n_102),
.B2(n_99),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_193),
.B1(n_204),
.B2(n_206),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_131),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_197),
.B(n_202),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_98),
.B(n_110),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g233 ( 
.A(n_190),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_192),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_131),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_14),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_198),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_130),
.B(n_138),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_180),
.B(n_13),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_203),
.B1(n_210),
.B2(n_212),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_201),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_99),
.B1(n_102),
.B2(n_132),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_26),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_8),
.B(n_15),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_219),
.B1(n_184),
.B2(n_163),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_29),
.B1(n_14),
.B2(n_12),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_158),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_29),
.B1(n_14),
.B2(n_12),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_178),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_11),
.C(n_10),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_162),
.C(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_11),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_235),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_221),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_230),
.C(n_241),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_174),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_237),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_161),
.C(n_170),
.Y(n_230)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_196),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_193),
.A2(n_168),
.B1(n_177),
.B2(n_164),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_187),
.B1(n_194),
.B2(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_179),
.C(n_164),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_168),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_207),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_195),
.Y(n_245)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_239),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_252),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_219),
.C(n_205),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_233),
.C(n_229),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_214),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_244),
.A2(n_209),
.B1(n_217),
.B2(n_218),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_198),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_189),
.B(n_207),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_214),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_194),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_264),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_191),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_263),
.A2(n_265),
.B1(n_232),
.B2(n_204),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_220),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_235),
.A2(n_202),
.B1(n_210),
.B2(n_190),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_247),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_267),
.A2(n_226),
.B1(n_232),
.B2(n_265),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_242),
.C(n_223),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_274),
.C(n_279),
.Y(n_298)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_223),
.C(n_221),
.Y(n_274)
);

AOI21x1_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_190),
.B(n_233),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_277),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_240),
.C(n_222),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_236),
.C(n_226),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_0),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_283),
.A2(n_258),
.B1(n_234),
.B2(n_211),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_254),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_287),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_253),
.B(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_296),
.C(n_280),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_254),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_250),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_289),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_257),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_294),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_293),
.B1(n_297),
.B2(n_269),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_9),
.C(n_2),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_266),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_299),
.B(n_4),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_300),
.A2(n_306),
.B(n_309),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_279),
.C(n_282),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_307),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_276),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_288),
.C(n_9),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_272),
.C(n_276),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_285),
.B(n_283),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_289),
.B(n_291),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_306),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_1),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_1),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_1),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_311),
.Y(n_326)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_322),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_302),
.C(n_5),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_328),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_312),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_327),
.B(n_324),
.C(n_323),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_324),
.C2(n_330),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_6),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_6),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_7),
.B(n_324),
.Y(n_335)
);


endmodule