module fake_netlist_6_285_n_130 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_3, n_14, n_0, n_4, n_22, n_13, n_11, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_130);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_13;
input n_11;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_130;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_127;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_129;
wire n_121;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_122;
wire n_45;
wire n_34;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_1),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_2),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_39),
.B1(n_33),
.B2(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_29),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_33),
.B1(n_6),
.B2(n_3),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_11),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR3xp33_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_3),
.C(n_6),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_8),
.Y(n_64)
);

OAI21x1_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_45),
.B(n_49),
.Y(n_65)
);

OAI21x1_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_45),
.B(n_49),
.Y(n_66)
);

AO31x2_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_54),
.A3(n_51),
.B(n_50),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_54),
.B(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_47),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_54),
.B(n_44),
.Y(n_71)
);

OAI21x1_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_44),
.B(n_49),
.Y(n_72)
);

OAI22x1_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_60),
.B1(n_55),
.B2(n_63),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

AOI21x1_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_49),
.B(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_58),
.B1(n_51),
.B2(n_50),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_69),
.B(n_62),
.C(n_48),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_43),
.B(n_57),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_43),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_67),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_66),
.B(n_13),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_86),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

OA21x2_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_80),
.B(n_75),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_88),
.B(n_81),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_86),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_91),
.B1(n_85),
.B2(n_87),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_98),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_102),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_95),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_93),
.B(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_102),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_100),
.B(n_89),
.C(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_114),
.B(n_108),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_89),
.B(n_94),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_107),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_118),
.C(n_112),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_111),
.C(n_116),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_111),
.C(n_113),
.Y(n_123)
);

NOR4xp25_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_117),
.C(n_18),
.D(n_24),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_15),
.Y(n_125)
);

OAI221xp5_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_79),
.B1(n_93),
.B2(n_94),
.C(n_121),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_126),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_79),
.B(n_93),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_94),
.B1(n_79),
.B2(n_93),
.Y(n_130)
);


endmodule