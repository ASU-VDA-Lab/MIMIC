module fake_jpeg_11791_n_304 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_165;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_294;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_46),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_50),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_8),
.C(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_16),
.B1(n_24),
.B2(n_41),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_52),
.B(n_58),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g116 ( 
.A(n_53),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_17),
.B(n_7),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx9p33_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_26),
.B(n_9),
.Y(n_60)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_5),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_67),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_0),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_19),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_70),
.Y(n_89)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_31),
.B(n_10),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_15),
.B(n_10),
.C(n_11),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_74),
.B(n_14),
.Y(n_126)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_44),
.A2(n_28),
.B1(n_25),
.B2(n_33),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_79),
.A2(n_91),
.B1(n_96),
.B2(n_101),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_85),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_37),
.B1(n_22),
.B2(n_28),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_120),
.B1(n_125),
.B2(n_100),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_43),
.B1(n_63),
.B2(n_48),
.Y(n_96)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx24_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_37),
.B1(n_22),
.B2(n_41),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_122),
.Y(n_128)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_54),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_118),
.B1(n_71),
.B2(n_42),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_119),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_113),
.A2(n_101),
.B1(n_109),
.B2(n_95),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_71),
.A2(n_36),
.B1(n_34),
.B2(n_16),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_61),
.A2(n_18),
.B1(n_35),
.B2(n_32),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_53),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_111),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_77),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_14),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_79),
.A2(n_74),
.B1(n_59),
.B2(n_35),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_127),
.A2(n_135),
.B1(n_133),
.B2(n_166),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_46),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_134),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_82),
.B(n_55),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_90),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_66),
.B1(n_73),
.B2(n_76),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_141),
.B1(n_161),
.B2(n_135),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_0),
.B(n_1),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_142),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_102),
.B1(n_96),
.B2(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_93),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_165),
.Y(n_171)
);

OR2x2_ASAP7_75t_SL g146 ( 
.A(n_93),
.B(n_88),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_168),
.B(n_117),
.C(n_97),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_84),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_152),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_92),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_154),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_87),
.Y(n_154)
);

INVx2_ASAP7_75t_R g156 ( 
.A(n_92),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_160),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_92),
.Y(n_157)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_114),
.B(n_83),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_86),
.B1(n_80),
.B2(n_98),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_105),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_156),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_105),
.A2(n_78),
.B1(n_97),
.B2(n_112),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_121),
.B1(n_169),
.B2(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_86),
.B(n_80),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_98),
.B(n_95),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_161),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_78),
.B(n_117),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_155),
.B1(n_153),
.B2(n_168),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_196),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_144),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_181),
.A2(n_157),
.B1(n_167),
.B2(n_189),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_184),
.A2(n_198),
.B1(n_179),
.B2(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_190),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_132),
.A2(n_148),
.B1(n_136),
.B2(n_159),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_187),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_201),
.B1(n_176),
.B2(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_130),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_150),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_140),
.B(n_132),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_146),
.A2(n_137),
.B(n_128),
.C(n_168),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

INVx3_ASAP7_75t_SL g218 ( 
.A(n_197),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_140),
.A2(n_159),
.B1(n_136),
.B2(n_145),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_184),
.B1(n_183),
.B2(n_179),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_145),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_193),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_143),
.A2(n_152),
.B1(n_158),
.B2(n_163),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_223),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_170),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_214),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_167),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_208),
.B(n_220),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_181),
.A2(n_175),
.B1(n_171),
.B2(n_199),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_206),
.Y(n_247)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_174),
.C(n_171),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_224),
.C(n_226),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_221),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_190),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_176),
.A2(n_196),
.B1(n_195),
.B2(n_185),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_183),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_221),
.B1(n_212),
.B2(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_173),
.C(n_197),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_173),
.C(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_242),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_219),
.A2(n_192),
.B(n_180),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_233),
.B(n_241),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_180),
.B(n_192),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_207),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_238),
.A2(n_218),
.B1(n_246),
.B2(n_247),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_210),
.B(n_204),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_222),
.C(n_224),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_182),
.A3(n_173),
.B1(n_220),
.B2(n_50),
.C1(n_111),
.C2(n_185),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_245),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_226),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_218),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_206),
.A2(n_212),
.B(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_252),
.Y(n_264)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_242),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_241),
.A2(n_246),
.B1(n_234),
.B2(n_245),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_262),
.A2(n_256),
.B1(n_252),
.B2(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g267 ( 
.A(n_263),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_253),
.B(n_229),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_244),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_269),
.A2(n_248),
.B1(n_273),
.B2(n_272),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_228),
.C(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_257),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_229),
.C(n_231),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_255),
.C(n_261),
.Y(n_277)
);

BUFx12_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_275),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_268),
.C(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_282),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_280),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_253),
.C(n_259),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_228),
.B1(n_254),
.B2(n_258),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_269),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_289),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_230),
.A3(n_275),
.B1(n_262),
.B2(n_270),
.C1(n_276),
.C2(n_267),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_275),
.A3(n_230),
.B1(n_276),
.B2(n_280),
.C1(n_279),
.C2(n_267),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_233),
.B(n_232),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_296),
.A2(n_290),
.B(n_287),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_285),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_297),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_295),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_302),
.B(n_301),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_303),
.Y(n_304)
);


endmodule