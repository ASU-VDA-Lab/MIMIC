module fake_jpeg_18620_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_7),
.B(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND4xp25_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.C(n_1),
.D(n_2),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_34),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_29),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_13),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_12),
.B(n_4),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_16),
.B(n_20),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_34),
.B1(n_28),
.B2(n_11),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_47),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_61),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_46),
.B1(n_42),
.B2(n_39),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_29),
.C(n_26),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.C(n_37),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_29),
.C(n_26),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_11),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_71),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_41),
.B(n_49),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_38),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_74),
.B1(n_46),
.B2(n_42),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_49),
.B1(n_39),
.B2(n_42),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_51),
.B1(n_58),
.B2(n_57),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_37),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_80),
.C(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_52),
.B1(n_51),
.B2(n_59),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_63),
.C(n_55),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_74),
.C(n_68),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_65),
.B1(n_15),
.B2(n_16),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_89),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_77),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_77),
.C(n_83),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_75),
.B(n_72),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_6),
.B(n_10),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_93),
.C(n_10),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_93),
.B(n_90),
.C(n_92),
.D(n_38),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_102),
.B(n_100),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_100),
.Y(n_104)
);


endmodule