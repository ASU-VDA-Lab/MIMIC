module fake_netlist_1_12040_n_666 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_666);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_666;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_393;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g76 ( .A(n_27), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_8), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_30), .Y(n_78) );
INVx1_ASAP7_75t_SL g79 ( .A(n_57), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_75), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_36), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_62), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_11), .Y(n_84) );
BUFx5_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_58), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_11), .Y(n_88) );
BUFx2_ASAP7_75t_L g89 ( .A(n_52), .Y(n_89) );
BUFx5_ASAP7_75t_L g90 ( .A(n_33), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_1), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_67), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_74), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_16), .Y(n_94) );
OR2x2_ASAP7_75t_L g95 ( .A(n_56), .B(n_20), .Y(n_95) );
NOR2xp33_ASAP7_75t_L g96 ( .A(n_29), .B(n_50), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_72), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_54), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_63), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_8), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_24), .B(n_68), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_64), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_49), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_35), .Y(n_104) );
BUFx8_ASAP7_75t_SL g105 ( .A(n_55), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_53), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_28), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_48), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_31), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_25), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_23), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_32), .Y(n_113) );
BUFx5_ASAP7_75t_L g114 ( .A(n_7), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_44), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_45), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_70), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_6), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_10), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_46), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_15), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_114), .Y(n_122) );
NOR2x1_ASAP7_75t_L g123 ( .A(n_80), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_114), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_85), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_114), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_76), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_114), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_114), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_114), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_89), .B(n_0), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_92), .B(n_1), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_77), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_83), .B(n_2), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_85), .B(n_3), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_93), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_85), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_105), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_87), .B(n_4), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_94), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_90), .Y(n_147) );
BUFx12f_ASAP7_75t_L g148 ( .A(n_78), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_102), .B(n_5), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_90), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_97), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_106), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_90), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_110), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_88), .B(n_7), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_90), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_112), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_113), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_90), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_120), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_111), .Y(n_161) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_91), .A2(n_119), .B(n_109), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_90), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_124), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_137), .B(n_115), .Y(n_165) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_134), .B(n_95), .Y(n_166) );
AO22x2_ASAP7_75t_L g167 ( .A1(n_149), .A2(n_101), .B1(n_79), .B2(n_118), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_128), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_162), .A2(n_100), .B1(n_81), .B2(n_108), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_122), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_135), .B(n_121), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_122), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_124), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_162), .A2(n_117), .B1(n_116), .B2(n_107), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_122), .Y(n_177) );
BUFx10_ASAP7_75t_L g178 ( .A(n_126), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_122), .Y(n_179) );
AND3x1_ASAP7_75t_L g180 ( .A(n_141), .B(n_101), .C(n_96), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_128), .Y(n_182) );
NAND3xp33_ASAP7_75t_L g183 ( .A(n_134), .B(n_104), .C(n_103), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
AO22x2_ASAP7_75t_L g185 ( .A1(n_149), .A2(n_9), .B1(n_10), .B2(n_12), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_128), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_137), .B(n_99), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_132), .B(n_98), .Y(n_190) );
INVxp67_ASAP7_75t_SL g191 ( .A(n_127), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_127), .Y(n_192) );
OR2x6_ASAP7_75t_L g193 ( .A(n_132), .B(n_12), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_138), .B(n_13), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_127), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g196 ( .A(n_127), .B(n_40), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_138), .B(n_13), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_146), .B(n_41), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_154), .B(n_14), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_128), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_154), .B(n_14), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_159), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_129), .Y(n_203) );
CKINVDCx6p67_ASAP7_75t_R g204 ( .A(n_148), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_129), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_159), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_129), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_129), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_130), .Y(n_209) );
OR2x6_ASAP7_75t_L g210 ( .A(n_123), .B(n_17), .Y(n_210) );
INVxp33_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_130), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_157), .B(n_158), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_157), .B(n_18), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_130), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_130), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_158), .B(n_19), .Y(n_217) );
OAI21xp33_ASAP7_75t_SL g218 ( .A1(n_160), .A2(n_21), .B(n_22), .Y(n_218) );
BUFx10_ASAP7_75t_L g219 ( .A(n_144), .Y(n_219) );
INVx4_ASAP7_75t_L g220 ( .A(n_193), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_197), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_197), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_193), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_197), .A2(n_162), .B1(n_160), .B2(n_123), .Y(n_224) );
NOR2x2_ASAP7_75t_L g225 ( .A(n_193), .B(n_148), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_165), .B(n_139), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_172), .B(n_187), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_172), .B(n_145), .Y(n_228) );
NAND2x1_ASAP7_75t_L g229 ( .A(n_199), .B(n_125), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_179), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_183), .B(n_155), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_190), .B(n_125), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_179), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_217), .B(n_199), .Y(n_234) );
AND2x6_ASAP7_75t_SL g235 ( .A(n_193), .B(n_140), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_213), .A2(n_163), .B(n_156), .C(n_153), .Y(n_236) );
AND2x6_ASAP7_75t_L g237 ( .A(n_217), .B(n_163), .Y(n_237) );
INVx5_ASAP7_75t_L g238 ( .A(n_174), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_190), .B(n_146), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_199), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_217), .B(n_146), .Y(n_241) );
NOR2xp67_ASAP7_75t_L g242 ( .A(n_218), .B(n_163), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_166), .B(n_146), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_188), .B(n_125), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_189), .B(n_156), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_201), .B(n_146), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_211), .A2(n_156), .B(n_153), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_166), .B(n_133), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_211), .A2(n_153), .B(n_133), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_194), .A2(n_143), .B(n_133), .C(n_150), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_178), .B(n_146), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_191), .B(n_143), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_179), .B(n_143), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_180), .A2(n_152), .B1(n_151), .B2(n_150), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_201), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_201), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_204), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_214), .B(n_150), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_214), .B(n_147), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_192), .B(n_147), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_192), .B(n_147), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_192), .B(n_142), .Y(n_263) );
NOR2xp67_ASAP7_75t_L g264 ( .A(n_194), .B(n_142), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_212), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_167), .A2(n_152), .B1(n_151), .B2(n_142), .Y(n_266) );
NAND3xp33_ASAP7_75t_SL g267 ( .A(n_169), .B(n_136), .C(n_152), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_210), .A2(n_152), .B1(n_151), .B2(n_136), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_176), .B(n_152), .Y(n_269) );
INVxp67_ASAP7_75t_L g270 ( .A(n_178), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_210), .A2(n_152), .B1(n_151), .B2(n_136), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_185), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_178), .B(n_151), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_167), .A2(n_151), .B1(n_128), .B2(n_37), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_210), .A2(n_26), .B1(n_34), .B2(n_38), .Y(n_275) );
INVx5_ASAP7_75t_L g276 ( .A(n_174), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_167), .A2(n_39), .B1(n_42), .B2(n_43), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_202), .A2(n_47), .B(n_51), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_212), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_234), .A2(n_167), .B1(n_185), .B2(n_210), .Y(n_280) );
OR2x6_ASAP7_75t_SL g281 ( .A(n_225), .B(n_219), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_220), .B(n_174), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_240), .A2(n_185), .B1(n_212), .B2(n_215), .Y(n_284) );
CKINVDCx16_ASAP7_75t_R g285 ( .A(n_247), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_226), .B(n_184), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_249), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_228), .B(n_164), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
BUFx12f_ASAP7_75t_L g290 ( .A(n_258), .Y(n_290) );
INVx4_ASAP7_75t_L g291 ( .A(n_223), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_270), .B(n_219), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_230), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_232), .Y(n_294) );
BUFx12f_ASAP7_75t_L g295 ( .A(n_235), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_272), .A2(n_196), .B(n_181), .C(n_175), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_248), .A2(n_203), .B(n_216), .Y(n_297) );
AOI22xp33_ASAP7_75t_SL g298 ( .A1(n_237), .A2(n_185), .B1(n_196), .B2(n_219), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_250), .A2(n_207), .B(n_205), .Y(n_299) );
NOR2xp33_ASAP7_75t_R g300 ( .A(n_267), .B(n_59), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_227), .B(n_206), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_231), .B(n_206), .Y(n_302) );
NOR2xp67_ASAP7_75t_SL g303 ( .A(n_221), .B(n_202), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_250), .A2(n_173), .B(n_208), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_229), .A2(n_198), .B(n_209), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_255), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_238), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_236), .A2(n_198), .B(n_209), .C(n_177), .Y(n_308) );
BUFx12f_ASAP7_75t_L g309 ( .A(n_238), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_264), .B(n_171), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_238), .B(n_171), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_221), .B(n_208), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_222), .A2(n_195), .B1(n_177), .B2(n_173), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_233), .Y(n_314) );
OAI21xp33_ASAP7_75t_SL g315 ( .A1(n_256), .A2(n_195), .B(n_65), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_222), .B(n_200), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_273), .B(n_200), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_257), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_252), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_259), .A2(n_170), .B(n_186), .Y(n_320) );
BUFx10_ASAP7_75t_L g321 ( .A(n_243), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_269), .A2(n_170), .B(n_66), .C(n_69), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_239), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_246), .B(n_168), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_266), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_238), .B(n_168), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_318), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_304), .A2(n_241), .B(n_260), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_305), .A2(n_278), .B(n_242), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_312), .Y(n_331) );
INVx2_ASAP7_75t_SL g332 ( .A(n_309), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_289), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_280), .A2(n_251), .B(n_259), .C(n_260), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_286), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_294), .B(n_288), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_290), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_284), .A2(n_237), .B1(n_274), .B2(n_224), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_304), .A2(n_261), .B(n_263), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_323), .A2(n_245), .B(n_244), .C(n_261), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_322), .A2(n_275), .B(n_271), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_287), .B(n_253), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
OAI222xp33_ASAP7_75t_L g345 ( .A1(n_298), .A2(n_277), .B1(n_268), .B2(n_279), .C1(n_262), .C2(n_254), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_320), .A2(n_276), .B(n_237), .Y(n_346) );
O2A1O1Ixp33_ASAP7_75t_L g347 ( .A1(n_301), .A2(n_237), .B(n_276), .C(n_182), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_325), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_283), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_298), .A2(n_237), .B1(n_276), .B2(n_182), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_289), .B(n_276), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_291), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_326), .A2(n_168), .B(n_182), .C(n_186), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_293), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_299), .A2(n_168), .B(n_182), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_320), .A2(n_186), .A3(n_71), .B(n_73), .Y(n_357) );
AOI21xp33_ASAP7_75t_L g358 ( .A1(n_296), .A2(n_186), .B(n_61), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_338), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_336), .B(n_291), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_336), .B(n_307), .Y(n_361) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_351), .B(n_297), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_335), .A2(n_296), .B(n_302), .C(n_315), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g364 ( .A(n_335), .B(n_303), .Y(n_364) );
OAI21x1_ASAP7_75t_SL g365 ( .A1(n_351), .A2(n_322), .B(n_308), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_348), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_343), .A2(n_295), .B1(n_306), .B2(n_321), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_348), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_356), .A2(n_297), .B(n_308), .Y(n_369) );
OA21x2_ASAP7_75t_L g370 ( .A1(n_358), .A2(n_299), .B(n_310), .Y(n_370) );
OAI21x1_ASAP7_75t_SL g371 ( .A1(n_341), .A2(n_314), .B(n_313), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_333), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_343), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_328), .B(n_292), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_333), .A2(n_281), .B1(n_300), .B2(n_321), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_328), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_329), .A2(n_324), .B(n_327), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_355), .B(n_319), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_349), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_355), .Y(n_380) );
AOI21x1_ASAP7_75t_L g381 ( .A1(n_330), .A2(n_311), .B(n_282), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_331), .B(n_316), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_338), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_331), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_344), .Y(n_385) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_362), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_372), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_376), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_366), .B(n_357), .Y(n_389) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_365), .A2(n_358), .B(n_345), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_372), .Y(n_391) );
AO21x2_ASAP7_75t_L g392 ( .A1(n_365), .A2(n_354), .B(n_346), .Y(n_392) );
OA21x2_ASAP7_75t_L g393 ( .A1(n_369), .A2(n_330), .B(n_342), .Y(n_393) );
OAI322xp33_ASAP7_75t_L g394 ( .A1(n_373), .A2(n_344), .A3(n_332), .B1(n_353), .B2(n_334), .C1(n_337), .C2(n_340), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_376), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_380), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_373), .B(n_339), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_380), .Y(n_400) );
OR2x6_ASAP7_75t_L g401 ( .A(n_362), .B(n_346), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_363), .A2(n_347), .B(n_342), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_368), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_384), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_377), .A2(n_357), .B(n_317), .Y(n_407) );
OA21x2_ASAP7_75t_L g408 ( .A1(n_381), .A2(n_357), .B(n_352), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_384), .B(n_357), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_385), .B(n_350), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_385), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_360), .B(n_357), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_374), .B(n_332), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_361), .B(n_350), .Y(n_415) );
INVx4_ASAP7_75t_L g416 ( .A(n_364), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_370), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_370), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_388), .B(n_378), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_388), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_417), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_417), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_413), .B(n_378), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_413), .B(n_361), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_395), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_413), .B(n_361), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_409), .B(n_350), .Y(n_427) );
AO21x2_ASAP7_75t_L g428 ( .A1(n_403), .A2(n_371), .B(n_382), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_406), .B(n_370), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_405), .B(n_397), .Y(n_430) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_387), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_417), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_418), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_402), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_402), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_418), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_406), .B(n_370), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_405), .B(n_379), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_416), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_406), .B(n_367), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_391), .B(n_364), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_391), .B(n_364), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_409), .B(n_375), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_397), .B(n_353), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_402), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_400), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_409), .B(n_352), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_400), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_404), .B(n_316), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_404), .B(n_371), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_398), .B(n_359), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_396), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_414), .B(n_383), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_389), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_414), .A2(n_398), .B1(n_402), .B2(n_390), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_396), .B(n_399), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_402), .B(n_399), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_396), .B(n_399), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_410), .B(n_389), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_441), .B(n_386), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_432), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_454), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_423), .B(n_415), .Y(n_469) );
AND2x4_ASAP7_75t_SL g470 ( .A(n_441), .B(n_416), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_454), .Y(n_471) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_458), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_423), .B(n_410), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_456), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_456), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_424), .B(n_415), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_465), .B(n_410), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_419), .B(n_389), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_420), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_420), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_458), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_424), .B(n_415), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_421), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_465), .B(n_416), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_425), .Y(n_486) );
OAI211xp5_ASAP7_75t_L g487 ( .A1(n_461), .A2(n_386), .B(n_416), .C(n_403), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_416), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_425), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_443), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_443), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_441), .B(n_415), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_419), .B(n_415), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_442), .B(n_390), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_449), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_426), .B(n_408), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_426), .B(n_450), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_449), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_450), .B(n_408), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_463), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_451), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_439), .B(n_408), .Y(n_503) );
AND2x4_ASAP7_75t_SL g504 ( .A(n_441), .B(n_401), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_430), .B(n_408), .Y(n_505) );
NOR4xp25_ASAP7_75t_SL g506 ( .A(n_431), .B(n_394), .C(n_407), .D(n_390), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_442), .B(n_390), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_460), .B(n_401), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_460), .B(n_401), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_427), .B(n_401), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_459), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_451), .B(n_446), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_457), .B(n_408), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_463), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_427), .B(n_446), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_440), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_447), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_427), .B(n_401), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_457), .B(n_401), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_444), .A2(n_407), .B1(n_412), .B2(n_394), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_447), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_478), .B(n_435), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_468), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_471), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_500), .B(n_429), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_497), .B(n_429), .Y(n_526) );
AND2x4_ASAP7_75t_SL g527 ( .A(n_510), .B(n_448), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_512), .B(n_461), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_492), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_473), .B(n_435), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_475), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_474), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_498), .B(n_427), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_517), .B(n_453), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_476), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_521), .B(n_453), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g537 ( .A(n_506), .B(n_445), .C(n_444), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_501), .B(n_438), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_485), .B(n_458), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_508), .B(n_438), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_501), .B(n_514), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_480), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_481), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_514), .B(n_469), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_508), .B(n_434), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_486), .B(n_464), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_489), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_490), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_491), .B(n_464), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_494), .B(n_433), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_511), .A2(n_452), .B1(n_428), .B2(n_392), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_496), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_499), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_509), .B(n_433), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_509), .B(n_433), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_488), .B(n_434), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_502), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_515), .B(n_462), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_516), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_519), .B(n_445), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_516), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_467), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_474), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_484), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_509), .B(n_455), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_515), .B(n_455), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_467), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_513), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_479), .B(n_462), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_505), .B(n_455), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_570), .B(n_507), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_563), .B(n_495), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_528), .B(n_477), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_564), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_541), .B(n_472), .Y(n_577) );
AOI21xp33_ASAP7_75t_SL g578 ( .A1(n_529), .A2(n_493), .B(n_466), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_560), .Y(n_579) );
INVxp33_ASAP7_75t_L g580 ( .A(n_529), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_562), .B(n_483), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_527), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_533), .B(n_518), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_525), .B(n_472), .Y(n_584) );
AOI322xp5_ASAP7_75t_L g585 ( .A1(n_525), .A2(n_518), .A3(n_510), .B1(n_482), .B2(n_466), .C1(n_484), .C2(n_436), .Y(n_585) );
OAI21xp33_ASAP7_75t_L g586 ( .A1(n_551), .A2(n_487), .B(n_510), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_527), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_526), .B(n_482), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_526), .B(n_504), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_523), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_544), .B(n_437), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_539), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_524), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_540), .B(n_504), .Y(n_594) );
OAI31xp33_ASAP7_75t_L g595 ( .A1(n_537), .A2(n_470), .A3(n_493), .B(n_466), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_540), .B(n_520), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_559), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_568), .B(n_437), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_538), .B(n_437), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_571), .B(n_422), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_559), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_532), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_534), .B(n_422), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_536), .B(n_422), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_532), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_531), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_565), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_535), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_596), .A2(n_561), .B1(n_569), .B2(n_551), .C(n_548), .Y(n_609) );
AOI211xp5_ASAP7_75t_L g610 ( .A1(n_595), .A2(n_561), .B(n_522), .C(n_530), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_586), .A2(n_547), .B1(n_543), .B2(n_542), .C(n_552), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_578), .B(n_572), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_597), .Y(n_613) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_580), .A2(n_553), .B(n_557), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_579), .B(n_558), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_590), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_582), .A2(n_567), .B1(n_555), .B2(n_554), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_582), .A2(n_567), .B1(n_555), .B2(n_554), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_587), .B(n_470), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_593), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_573), .B(n_568), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_574), .B(n_545), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_588), .B(n_545), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_SL g624 ( .A1(n_602), .A2(n_566), .B(n_565), .C(n_421), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_585), .A2(n_549), .B1(n_546), .B2(n_550), .C(n_556), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_608), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_606), .Y(n_627) );
AOI211xp5_ASAP7_75t_SL g628 ( .A1(n_589), .A2(n_452), .B(n_566), .C(n_434), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_588), .B(n_589), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_574), .Y(n_630) );
NAND4xp25_ASAP7_75t_SL g631 ( .A(n_610), .B(n_594), .C(n_584), .D(n_592), .Y(n_631) );
AND4x1_ASAP7_75t_L g632 ( .A(n_628), .B(n_583), .C(n_594), .D(n_575), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_630), .B(n_599), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_616), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_620), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_611), .B(n_576), .C(n_583), .D(n_581), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_625), .A2(n_587), .B1(n_576), .B2(n_601), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_619), .A2(n_580), .B(n_601), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_626), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_612), .A2(n_577), .B(n_599), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_629), .B(n_598), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_623), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_613), .A2(n_607), .B(n_605), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_631), .B(n_613), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_SL g645 ( .A1(n_640), .A2(n_624), .B(n_609), .C(n_614), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_642), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_636), .A2(n_615), .B1(n_627), .B2(n_621), .C(n_622), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_637), .A2(n_618), .B1(n_617), .B2(n_615), .Y(n_648) );
NAND4xp75_ASAP7_75t_L g649 ( .A(n_638), .B(n_600), .C(n_604), .D(n_603), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_636), .A2(n_598), .B1(n_591), .B2(n_602), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_632), .A2(n_607), .B1(n_605), .B2(n_436), .C(n_407), .Y(n_651) );
NAND4xp25_ASAP7_75t_SL g652 ( .A(n_651), .B(n_643), .C(n_633), .D(n_639), .Y(n_652) );
XOR2xp5_ASAP7_75t_L g653 ( .A(n_648), .B(n_635), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_650), .B(n_634), .Y(n_654) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_645), .B(n_641), .C(n_436), .Y(n_655) );
NOR3xp33_ASAP7_75t_SL g656 ( .A(n_652), .B(n_644), .C(n_649), .Y(n_656) );
AO211x2_ASAP7_75t_L g657 ( .A1(n_655), .A2(n_647), .B(n_646), .C(n_407), .Y(n_657) );
INVxp33_ASAP7_75t_SL g658 ( .A(n_653), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_658), .Y(n_659) );
NOR2x1p5_ASAP7_75t_L g660 ( .A(n_656), .B(n_654), .Y(n_660) );
OAI22x1_ASAP7_75t_L g661 ( .A1(n_660), .A2(n_657), .B1(n_407), .B2(n_393), .Y(n_661) );
XNOR2x1_ASAP7_75t_L g662 ( .A(n_661), .B(n_659), .Y(n_662) );
OAI22xp5_ASAP7_75t_SL g663 ( .A1(n_662), .A2(n_393), .B1(n_412), .B2(n_392), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_392), .B1(n_428), .B2(n_393), .Y(n_664) );
OA211x2_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_392), .B(n_428), .C(n_393), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_665), .A2(n_428), .B1(n_393), .B2(n_412), .Y(n_666) );
endmodule