module real_jpeg_14599_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_312, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_312;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_2),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_42),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_2),
.A2(n_42),
.B1(n_58),
.B2(n_62),
.Y(n_234)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_4),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_96),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_4),
.A2(n_58),
.B1(n_62),
.B2(n_96),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_96),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_6),
.A2(n_29),
.B1(n_58),
.B2(n_62),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_6),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_58),
.B1(n_62),
.B2(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_67),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_10),
.A2(n_37),
.B1(n_58),
.B2(n_62),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_10),
.A2(n_37),
.B1(n_48),
.B2(n_49),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_11),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_11),
.A2(n_58),
.B1(n_62),
.B2(n_137),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_137),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_137),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g230 ( 
.A(n_12),
.B(n_33),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_13),
.A2(n_58),
.B1(n_62),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_13),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_142),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_142),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_142),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_14),
.A2(n_53),
.B1(n_58),
.B2(n_62),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_15),
.A2(n_48),
.B1(n_49),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_15),
.B(n_58),
.C(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_47),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_15),
.A2(n_140),
.B(n_143),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_15),
.A2(n_32),
.B(n_46),
.C(n_171),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_15),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_15),
.B(n_25),
.Y(n_217)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_110),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_20),
.B(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_70),
.C(n_78),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_21),
.B(n_70),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_38),
.B2(n_69),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_22),
.A2(n_23),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_23),
.B(n_39),
.C(n_55),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_24),
.A2(n_31),
.B(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_26),
.A2(n_30),
.B(n_125),
.C(n_216),
.Y(n_215)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_26),
.A2(n_32),
.A3(n_34),
.B1(n_217),
.B2(n_230),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_30),
.A2(n_31),
.B1(n_244),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_30),
.A2(n_264),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_31),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_31),
.B(n_95),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_31),
.A2(n_92),
.B(n_244),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_54),
.B1(n_55),
.B2(n_68),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_47),
.B2(n_51),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_43),
.B(n_178),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_45),
.A2(n_48),
.B(n_125),
.Y(n_171)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_47),
.B(n_178),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_64)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_49),
.B(n_129),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_52),
.A2(n_72),
.B1(n_74),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_55),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B(n_65),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_63),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_56),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_56),
.A2(n_63),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_56),
.A2(n_63),
.B1(n_223),
.B2(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_56),
.A2(n_63),
.B1(n_89),
.B2(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_57),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_57),
.B(n_125),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_57),
.A2(n_138),
.B(n_222),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_62),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_63),
.B(n_127),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_70),
.A2(n_71),
.B(n_75),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_72),
.A2(n_176),
.B(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_72),
.A2(n_74),
.B1(n_191),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_72),
.A2(n_177),
.B(n_220),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_266),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_74),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_74),
.A2(n_192),
.B(n_266),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_76),
.A2(n_126),
.B(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_78),
.B(n_308),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B(n_91),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_79),
.A2(n_80),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_81),
.A2(n_82),
.B1(n_91),
.B2(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_83),
.A2(n_84),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_83),
.B(n_144),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_83),
.A2(n_84),
.B1(n_234),
.B2(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_84),
.B(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_86),
.A2(n_140),
.B1(n_157),
.B2(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_91),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_306),
.B(n_310),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_293),
.B(n_305),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_276),
.B(n_292),
.Y(n_114)
);

OAI321xp33_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_236),
.A3(n_269),
.B1(n_274),
.B2(n_275),
.C(n_312),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_208),
.B(n_235),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_185),
.B(n_207),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_166),
.B(n_184),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_145),
.B(n_165),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_130),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_121),
.B(n_130),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_128),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_123),
.B1(n_128),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_157),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_139),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_135),
.C(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B(n_143),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_140),
.A2(n_157),
.B1(n_173),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_140),
.A2(n_157),
.B1(n_199),
.B2(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_153),
.B(n_164),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_151),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_159),
.B(n_163),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_156),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_158),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_168),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_179),
.C(n_183),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_172),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_174)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_186),
.B(n_187),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_200),
.B2(n_201),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_203),
.C(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_194),
.C(n_198),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_209),
.B(n_210),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_225),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_226),
.C(n_227),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_218),
.B2(n_224),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_219),
.C(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_253),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_247),
.C(n_252),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_238),
.A2(n_239),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_245),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_245),
.C(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_247),
.B(n_252),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_250),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_268),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_261),
.C(n_268),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_259),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_267),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_265),
.C(n_267),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_291),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_291),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_289),
.B2(n_290),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_287),
.C(n_290),
.Y(n_304)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_295),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_304),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_299),
.C(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_309),
.Y(n_310)
);


endmodule