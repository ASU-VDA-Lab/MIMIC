module real_jpeg_9878_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_41;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_63),
.B1(n_69),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_72),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_72),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_5),
.A2(n_63),
.B1(n_69),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_5),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_90),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_90),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_90),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_70),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_12),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_12),
.A2(n_53),
.B(n_65),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_12),
.A2(n_63),
.B1(n_69),
.B2(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_12),
.B(n_166),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_12),
.A2(n_38),
.B(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_12),
.B(n_38),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_217),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_12),
.A2(n_52),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_52),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_58),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_13),
.A2(n_58),
.B1(n_63),
.B2(n_69),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_58),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_15),
.A2(n_63),
.B1(n_69),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_15),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_139),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_139),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_139),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_16),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_16),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_17),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_94),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_21),
.B(n_94),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_80),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_22),
.A2(n_23),
.B1(n_74),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_60),
.C(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_25),
.B(n_36),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_26),
.A2(n_33),
.B(n_34),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_26),
.A2(n_33),
.B1(n_83),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_26),
.A2(n_33),
.B1(n_200),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_26),
.A2(n_33),
.B1(n_202),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_26),
.A2(n_33),
.B1(n_233),
.B2(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_27),
.A2(n_28),
.B1(n_147),
.B2(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_27),
.A2(n_28),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_30),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_29),
.B(n_45),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_29),
.B(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_30),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_33),
.B(n_143),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_41),
.B1(n_44),
.B2(n_85),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_39),
.B1(n_51),
.B2(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_38),
.B(n_56),
.Y(n_246)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_39),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_44),
.B1(n_46),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_41),
.A2(n_44),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_41),
.A2(n_44),
.B1(n_208),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_41),
.A2(n_44),
.B1(n_231),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_41),
.A2(n_44),
.B1(n_169),
.B2(n_239),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_43),
.Y(n_212)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_44),
.B(n_143),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_60),
.B1(n_61),
.B2(n_73),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_55),
.B1(n_57),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_50),
.A2(n_55),
.B1(n_93),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_50),
.A2(n_55),
.B1(n_134),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_50),
.A2(n_55),
.B1(n_162),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_50),
.A2(n_55),
.B1(n_186),
.B2(n_241),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_54),
.C(n_55),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_67)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_54),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_55),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_55),
.B(n_143),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_59),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_62),
.A2(n_67),
.B1(n_71),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_62),
.A2(n_67),
.B1(n_89),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.C(n_67),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_64),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_63),
.A2(n_64),
.B(n_143),
.C(n_144),
.Y(n_142)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_67),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_74),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_76),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_80),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.C(n_91),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_82),
.B(n_84),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_86),
.A2(n_101),
.B1(n_104),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_120),
.B2(n_121),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_111),
.B2(n_112),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_105),
.B(n_110),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_105),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_120),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_151),
.B(n_273),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_148),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_126),
.B(n_148),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.C(n_130),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_129),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_131),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_135),
.C(n_140),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_140),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_191),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_173),
.B(n_190),
.Y(n_153)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_154),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_170),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_155),
.B(n_170),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_167),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_161),
.B1(n_167),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_174),
.B(n_176),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.C(n_182),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_177),
.B(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_180),
.A2(n_182),
.B1(n_183),
.B2(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_180),
.Y(n_269)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_188),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_184),
.A2(n_185),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_187),
.B(n_188),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_189),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_271),
.C(n_272),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_265),
.B(n_270),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_251),
.B(n_264),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_235),
.B(n_250),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_225),
.B(n_234),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_214),
.B(n_224),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_198),
.B(n_203),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_209),
.B2(n_213),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_213),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_207),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_209),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_219),
.B(n_223),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_218),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_226),
.B(n_227),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_230),
.C(n_232),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_237),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_237),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.CI(n_243),
.CON(n_237),
.SN(n_237)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_261),
.C(n_262),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_260),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_261),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);


endmodule