module fake_jpeg_18464_n_300 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_265;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_40),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_15),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_23),
.B1(n_31),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_15),
.B1(n_40),
.B2(n_25),
.Y(n_75)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_23),
.B1(n_31),
.B2(n_33),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_36),
.B1(n_25),
.B2(n_14),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_44),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_59),
.B(n_60),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_15),
.B1(n_24),
.B2(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_90),
.B1(n_98),
.B2(n_25),
.Y(n_103)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_31),
.B1(n_33),
.B2(n_15),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_74),
.B1(n_75),
.B2(n_91),
.Y(n_104)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_86),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_44),
.C(n_36),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_72),
.C(n_37),
.Y(n_108)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_44),
.C(n_36),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_38),
.B1(n_40),
.B2(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_76),
.B(n_81),
.Y(n_119)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_77),
.Y(n_123)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_87),
.Y(n_120)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_88),
.B(n_92),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_24),
.B1(n_29),
.B2(n_14),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_100),
.C(n_101),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_24),
.B1(n_29),
.B2(n_21),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_26),
.B1(n_16),
.B2(n_27),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_21),
.B1(n_27),
.B2(n_16),
.Y(n_130)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_0),
.B(n_1),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_115),
.B(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_82),
.B1(n_87),
.B2(n_100),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_74),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_2),
.B(n_3),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_2),
.B(n_3),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_62),
.A2(n_2),
.B(n_4),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_126),
.B(n_131),
.C(n_17),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_4),
.B(n_17),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_16),
.B1(n_21),
.B2(n_27),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_4),
.B(n_17),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_134),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_135),
.B1(n_129),
.B2(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2x1p5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_138),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_142),
.B1(n_146),
.B2(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_145),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_123),
.C(n_28),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_80),
.B1(n_37),
.B2(n_35),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_80),
.B1(n_37),
.B2(n_35),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_149),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_39),
.B1(n_24),
.B2(n_29),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_89),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_102),
.A2(n_39),
.B1(n_41),
.B2(n_79),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_154),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_39),
.B1(n_29),
.B2(n_41),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_157),
.B1(n_114),
.B2(n_122),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_96),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_19),
.B1(n_73),
.B2(n_17),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_109),
.B1(n_113),
.B2(n_17),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_85),
.B1(n_68),
.B2(n_19),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_121),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_109),
.A2(n_17),
.B1(n_20),
.B2(n_6),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_163),
.B(n_169),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_171),
.B(n_181),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_129),
.B1(n_114),
.B2(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_115),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_124),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_174),
.B(n_185),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_145),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_28),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_156),
.C(n_142),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_122),
.B1(n_113),
.B2(n_112),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_140),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_189),
.B(n_18),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_111),
.B(n_4),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_207),
.C(n_164),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_206),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_196),
.B1(n_209),
.B2(n_213),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_148),
.B1(n_144),
.B2(n_111),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_202),
.B1(n_208),
.B2(n_180),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_159),
.A2(n_19),
.B1(n_18),
.B2(n_30),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_30),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_178),
.B(n_30),
.Y(n_205)
);

AOI31xp67_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_20),
.A3(n_32),
.B(n_18),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_20),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_159),
.A2(n_18),
.B1(n_32),
.B2(n_20),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_32),
.B1(n_18),
.B2(n_8),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_206),
.B(n_211),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_32),
.B(n_7),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_222),
.B(n_210),
.Y(n_236)
);

OAI22x1_ASAP7_75t_SL g219 ( 
.A1(n_201),
.A2(n_189),
.B1(n_161),
.B2(n_171),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_223),
.B1(n_228),
.B2(n_229),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_176),
.B1(n_167),
.B2(n_168),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_230),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_160),
.B(n_163),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_169),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_214),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_168),
.B1(n_187),
.B2(n_166),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_182),
.C(n_173),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_162),
.Y(n_233)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_236),
.A2(n_216),
.B1(n_164),
.B2(n_171),
.Y(n_264)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_217),
.A2(n_196),
.B1(n_197),
.B2(n_191),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_245),
.B1(n_252),
.B2(n_218),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_244),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_198),
.B1(n_190),
.B2(n_166),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_162),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_190),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_202),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_208),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_205),
.CI(n_232),
.CON(n_253),
.SN(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_221),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_257),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_260),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_230),
.C(n_164),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_266),
.C(n_249),
.Y(n_275)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_237),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_207),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_226),
.C(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_273),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_272),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_237),
.C(n_241),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_252),
.C(n_244),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_276),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_257),
.C(n_262),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_226),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_260),
.B1(n_265),
.B2(n_275),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_267),
.A2(n_254),
.B1(n_248),
.B2(n_239),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_282),
.B(n_283),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_271),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_264),
.B(n_256),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_174),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_248),
.B(n_224),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_287),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_281),
.A2(n_256),
.B(n_227),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_284),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_280),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_279),
.B(n_289),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_253),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_295),
.A2(n_294),
.B(n_227),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_297),
.A2(n_250),
.B(n_251),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_171),
.B(n_188),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_183),
.Y(n_300)
);


endmodule