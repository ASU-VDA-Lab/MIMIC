module real_jpeg_3726_n_31 (n_17, n_8, n_0, n_21, n_168, n_2, n_29, n_10, n_175, n_9, n_12, n_24, n_166, n_170, n_6, n_176, n_28, n_171, n_169, n_167, n_23, n_11, n_14, n_172, n_25, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_1, n_26, n_27, n_20, n_19, n_30, n_16, n_15, n_13, n_31);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_29;
input n_10;
input n_175;
input n_9;
input n_12;
input n_24;
input n_166;
input n_170;
input n_6;
input n_176;
input n_28;
input n_171;
input n_169;
input n_167;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_30;
input n_16;
input n_15;
input n_13;

output n_31;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_80;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_1),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_2),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_3),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_4),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_5),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_6),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_9),
.B(n_54),
.Y(n_138)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_10),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_11),
.A2(n_72),
.B1(n_104),
.B2(n_107),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_12),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_14),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_15),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_16),
.B(n_67),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_17),
.A2(n_81),
.B(n_85),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_74),
.C(n_98),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_19),
.B(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_19),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_20),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_22),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_23),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_24),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_25),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_82),
.Y(n_81)
);

AO22x1_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_77),
.B1(n_79),
.B2(n_90),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_76),
.C(n_91),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_35),
.B1(n_145),
.B2(n_148),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_30),
.B(n_37),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_30),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_30),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_30),
.B(n_151),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_30),
.A2(n_146),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_160),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_154),
.B(n_159),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_150),
.B(n_153),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_44),
.B(n_144),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_39),
.B(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_40),
.B(n_143),
.Y(n_142)
);

BUFx4f_ASAP7_75t_SL g158 ( 
.A(n_40),
.Y(n_158)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_43),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_140),
.C(n_141),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_51),
.B(n_139),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_47),
.B(n_50),
.Y(n_139)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_57),
.C(n_138),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_56),
.B(n_152),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_134),
.C(n_135),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_65),
.B(n_133),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_60),
.B(n_64),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_108),
.Y(n_107)
);

OAI221xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_109),
.C(n_123),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_68),
.B(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_100),
.C(n_101),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_93),
.C(n_94),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.C(n_89),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_88),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_124),
.A3(n_125),
.B1(n_128),
.B2(n_129),
.C1(n_132),
.C2(n_176),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.C(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_166),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_167),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_168),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_169),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_170),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_171),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_172),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_173),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_174),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_175),
.Y(n_122)
);


endmodule