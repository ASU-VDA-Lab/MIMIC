module fake_jpeg_27542_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_29),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_27),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_11),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_22),
.B1(n_14),
.B2(n_11),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_44)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_25),
.B1(n_14),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_32),
.B1(n_23),
.B2(n_16),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_50),
.B1(n_33),
.B2(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_24),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_34),
.B(n_35),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_48),
.B(n_42),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_32),
.B1(n_40),
.B2(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_61),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

AO21x1_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_43),
.B(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_58),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_51),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_52),
.B(n_55),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

OAI22x1_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_69),
.B1(n_67),
.B2(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_20),
.B1(n_18),
.B2(n_5),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_63),
.B1(n_45),
.B2(n_46),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_80),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_60),
.A3(n_54),
.B1(n_61),
.B2(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_65),
.B1(n_72),
.B2(n_46),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_65),
.B(n_2),
.C(n_3),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_73),
.C(n_20),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_92),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_7),
.B(n_10),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_18),
.C(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_1),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_84),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_9),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_93),
.B(n_86),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_1),
.A3(n_2),
.B1(n_5),
.B2(n_6),
.C1(n_86),
.C2(n_98),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_100),
.C(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_2),
.Y(n_103)
);


endmodule