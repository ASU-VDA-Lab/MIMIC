module real_jpeg_9506_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx24_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_1),
.A2(n_26),
.B1(n_29),
.B2(n_48),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_3),
.A2(n_53),
.B1(n_62),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_3),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_102),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_3),
.A2(n_26),
.B1(n_29),
.B2(n_102),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_102),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_SL g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_9),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_9),
.A2(n_55),
.B(n_59),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_9),
.A2(n_53),
.B1(n_62),
.B2(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_66),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_9),
.A2(n_37),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_9),
.B(n_37),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_9),
.A2(n_82),
.B1(n_83),
.B2(n_226),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_10),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_10),
.A2(n_34),
.B1(n_53),
.B2(n_62),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_10),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_11),
.A2(n_28),
.B1(n_58),
.B2(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_11),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_11),
.A2(n_28),
.B1(n_53),
.B2(n_62),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_13),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_13),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_13),
.A2(n_26),
.B1(n_29),
.B2(n_63),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_63),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_14),
.A2(n_26),
.B1(n_29),
.B2(n_41),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_15),
.A2(n_53),
.B1(n_62),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_15),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_146),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_15),
.A2(n_37),
.B1(n_38),
.B2(n_146),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_15),
.A2(n_26),
.B1(n_29),
.B2(n_146),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_19),
.B(n_106),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_79),
.C(n_90),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_20),
.A2(n_21),
.B1(n_79),
.B2(n_156),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_50),
.C(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_23),
.B(n_35),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_24),
.A2(n_83),
.B(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_31),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_26),
.A2(n_29),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_26),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_217)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_29),
.B(n_46),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_29),
.B(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_30),
.A2(n_31),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_31),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_32),
.A2(n_82),
.B(n_210),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_36),
.A2(n_45),
.B(n_96),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_43),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_38),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_37),
.B(n_70),
.Y(n_254)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_38),
.A2(n_75),
.B1(n_249),
.B2(n_254),
.Y(n_253)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_47),
.B(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_42),
.A2(n_45),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_42),
.A2(n_45),
.B1(n_216),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_42),
.A2(n_45),
.B1(n_239),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_42),
.A2(n_122),
.B(n_247),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_44),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_45),
.B(n_150),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_67),
.B2(n_78),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_61),
.B(n_64),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_57),
.B1(n_61),
.B2(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_52),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_52),
.A2(n_57),
.B1(n_101),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_52),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B(n_56),
.C(n_57),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_53),
.A2(n_54),
.B(n_150),
.C(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_69),
.B(n_70),
.C(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_70),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g249 ( 
.A(n_59),
.B(n_150),
.CON(n_249),
.SN(n_249)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_66),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_73),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_77),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_68),
.A2(n_140),
.B1(n_141),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_68),
.A2(n_140),
.B1(n_171),
.B2(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_68),
.B(n_150),
.Y(n_237)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_74),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_69),
.B(n_104),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_69),
.A2(n_74),
.B1(n_194),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_74),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_79),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_89),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_81),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_85),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_82),
.A2(n_83),
.B1(n_208),
.B2(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_82),
.A2(n_84),
.B(n_94),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_83),
.B(n_150),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_87),
.A2(n_98),
.B(n_124),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_90),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.C(n_103),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_95),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_106),
.Y(n_281)
);

FAx1_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.CI(n_126),
.CON(n_106),
.SN(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_115),
.B2(n_116),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_115),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B(n_125),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_157),
.B(n_280),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_154),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_131),
.B(n_154),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_136),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_135),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_136),
.A2(n_137),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.C(n_147),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B(n_142),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_199),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_180),
.B(n_198),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_200),
.C(n_279),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_177),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_177),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_176),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_170),
.B1(n_176),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_181),
.B(n_183),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_184),
.B(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_187),
.A2(n_189),
.B1(n_190),
.B2(n_277),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_187),
.Y(n_277)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.C(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_191),
.A2(n_192),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_195),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_273),
.B(n_278),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_258),
.B(n_272),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_242),
.B(n_257),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_233),
.B(n_241),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_222),
.B(n_232),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_211),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_217),
.B2(n_221),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_212),
.B(n_221),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_217),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_227),
.B(n_231),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_225),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_243),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.CI(n_240),
.CON(n_236),
.SN(n_236)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_252),
.B2(n_256),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_251),
.C(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_252),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_260),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_266),
.B2(n_267),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_269),
.C(n_270),
.Y(n_274)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_268),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_269),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);


endmodule