module fake_jpeg_11176_n_578 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_578);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_578;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_65),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_32),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_73),
.B(n_86),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_32),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_75),
.B(n_106),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_76),
.Y(n_174)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_101),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_35),
.B(n_17),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_34),
.Y(n_103)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_35),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_27),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_1),
.Y(n_150)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_47),
.B1(n_51),
.B2(n_28),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_118),
.A2(n_132),
.B1(n_136),
.B2(n_145),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_53),
.B1(n_54),
.B2(n_34),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_119),
.A2(n_151),
.B1(n_170),
.B2(n_19),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_81),
.A2(n_28),
.B1(n_34),
.B2(n_54),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_27),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_134),
.B(n_142),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_87),
.A2(n_54),
.B1(n_53),
.B2(n_27),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_37),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_58),
.A2(n_79),
.B1(n_68),
.B2(n_102),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_159),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_61),
.A2(n_53),
.B1(n_48),
.B2(n_46),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_57),
.B(n_37),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_66),
.A2(n_53),
.B1(n_52),
.B2(n_49),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_25),
.B1(n_21),
.B2(n_26),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_74),
.A2(n_38),
.B1(n_48),
.B2(n_46),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_67),
.B(n_38),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_80),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_76),
.B(n_45),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_45),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_131),
.B(n_143),
.C(n_122),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_176),
.B(n_189),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_39),
.B1(n_24),
.B2(n_60),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_96),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_178),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_179),
.B(n_203),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_78),
.B1(n_83),
.B2(n_98),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_181),
.A2(n_182),
.B1(n_220),
.B2(n_227),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_200),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_92),
.B1(n_91),
.B2(n_95),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_185),
.A2(n_152),
.B1(n_168),
.B2(n_138),
.Y(n_268)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_186),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_187),
.B(n_228),
.Y(n_241)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_188),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_113),
.A2(n_39),
.B(n_49),
.C(n_19),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_191),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_111),
.B(n_19),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_193),
.B(n_196),
.Y(n_289)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_112),
.B(n_36),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_114),
.Y(n_197)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_197),
.Y(n_249)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_123),
.B(n_90),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_225),
.C(n_230),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_89),
.B1(n_93),
.B2(n_52),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_202),
.A2(n_212),
.B1(n_156),
.B2(n_161),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_126),
.B(n_36),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_128),
.B(n_36),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_204),
.B(n_206),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_146),
.B(n_52),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_207),
.Y(n_271)
);

INVx5_ASAP7_75t_SL g208 ( 
.A(n_130),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_208),
.Y(n_283)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_211),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_119),
.A2(n_69),
.B1(n_21),
.B2(n_49),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_130),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g214 ( 
.A1(n_149),
.A2(n_71),
.B1(n_33),
.B2(n_26),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_214),
.A2(n_167),
.B(n_133),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_137),
.Y(n_216)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_217),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_124),
.A2(n_33),
.B1(n_21),
.B2(n_25),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_33),
.B1(n_26),
.B2(n_25),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_141),
.B(n_109),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_223),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_127),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_171),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g226 ( 
.A(n_175),
.Y(n_226)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_132),
.A2(n_109),
.B1(n_110),
.B2(n_4),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_115),
.B(n_2),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_162),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_235),
.Y(n_253)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_153),
.Y(n_232)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_139),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_234),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_175),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_125),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_238),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_129),
.B(n_3),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_120),
.C(n_5),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_133),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_180),
.A2(n_118),
.B(n_167),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_244),
.A2(n_279),
.B(n_178),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_248),
.A2(n_280),
.B(n_214),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_266),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_187),
.A2(n_125),
.B1(n_156),
.B2(n_117),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_263),
.A2(n_269),
.B1(n_178),
.B2(n_229),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_193),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_181),
.A2(n_162),
.B1(n_117),
.B2(n_174),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_L g325 ( 
.A1(n_267),
.A2(n_268),
.B1(n_286),
.B2(n_191),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_7),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_194),
.B(n_161),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_285),
.Y(n_314)
);

AOI22x1_ASAP7_75t_L g279 ( 
.A1(n_230),
.A2(n_168),
.B1(n_152),
.B2(n_138),
.Y(n_279)
);

AOI32xp33_ASAP7_75t_L g280 ( 
.A1(n_237),
.A2(n_174),
.A3(n_129),
.B1(n_6),
.B2(n_7),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_196),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_281),
.B(n_192),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_220),
.A2(n_206),
.B1(n_204),
.B2(n_203),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_294),
.B1(n_212),
.B2(n_225),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_201),
.B(n_3),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_226),
.A2(n_195),
.B1(n_190),
.B2(n_232),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_179),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_291),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_295),
.B(n_297),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_296),
.A2(n_303),
.B1(n_308),
.B2(n_315),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_309),
.B1(n_310),
.B2(n_317),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_300),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_189),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_323),
.Y(n_348)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_282),
.A2(n_214),
.B1(n_176),
.B2(n_211),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_248),
.A2(n_215),
.B(n_208),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_304),
.A2(n_275),
.B(n_274),
.Y(n_356)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_222),
.B1(n_210),
.B2(n_198),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_241),
.A2(n_269),
.B1(n_262),
.B2(n_289),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_241),
.A2(n_197),
.B1(n_199),
.B2(n_224),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_199),
.C(n_228),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_318),
.C(n_332),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_291),
.Y(n_312)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_255),
.Y(n_313)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_272),
.A2(n_236),
.B1(n_186),
.B2(n_209),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_241),
.B(n_217),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_316),
.A2(n_287),
.B(n_284),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_262),
.A2(n_216),
.B1(n_233),
.B2(n_219),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_289),
.C(n_242),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_246),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_324),
.Y(n_351)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_255),
.Y(n_320)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_320),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_321),
.B(n_341),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_238),
.B(n_207),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_322),
.A2(n_271),
.B(n_258),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_246),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_325),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_188),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_327),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_242),
.B(n_8),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_251),
.B(n_245),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_328),
.B(n_331),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_244),
.A2(n_183),
.B1(n_9),
.B2(n_10),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_329),
.A2(n_340),
.B1(n_283),
.B2(n_292),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_250),
.B(n_8),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_336),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_250),
.B(n_183),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_253),
.B(n_183),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_246),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_239),
.B(n_8),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_334),
.Y(n_345)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_335),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_290),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_260),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_339),
.Y(n_361)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_277),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_260),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_268),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_276),
.B(n_17),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_342),
.Y(n_363)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_275),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_273),
.B(n_9),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_274),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_299),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_353),
.B(n_366),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_311),
.C(n_332),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_380),
.C(n_384),
.Y(n_399)
);

AO22x1_ASAP7_75t_L g392 ( 
.A1(n_356),
.A2(n_385),
.B1(n_381),
.B2(n_351),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_323),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_371),
.Y(n_397)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_334),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_316),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_382),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_374),
.A2(n_387),
.B1(n_388),
.B2(n_310),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_301),
.B(n_294),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_309),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_314),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_304),
.A2(n_279),
.B(n_264),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_379),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_279),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_316),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_326),
.B(n_287),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_300),
.A2(n_284),
.B(n_243),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_308),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_297),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_296),
.A2(n_315),
.B1(n_303),
.B2(n_329),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_298),
.A2(n_292),
.B1(n_243),
.B2(n_254),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_324),
.B1(n_333),
.B2(n_319),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_390),
.A2(n_413),
.B1(n_414),
.B2(n_421),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_356),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_391),
.A2(n_360),
.B(n_378),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_392),
.A2(n_360),
.B(n_375),
.Y(n_436)
);

XOR2x2_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_330),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_394),
.B(n_271),
.Y(n_458)
);

FAx1_ASAP7_75t_SL g395 ( 
.A(n_348),
.B(n_312),
.CI(n_295),
.CON(n_395),
.SN(n_395)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_424),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_422),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_321),
.C(n_342),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_401),
.B(n_404),
.C(n_411),
.Y(n_456)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_343),
.C(n_339),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_361),
.Y(n_407)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_408),
.A2(n_419),
.B1(n_420),
.B2(n_381),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_254),
.Y(n_454)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_302),
.C(n_337),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_348),
.B(n_376),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_412),
.B(n_423),
.C(n_425),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_386),
.A2(n_362),
.B1(n_353),
.B2(n_381),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_365),
.A2(n_322),
.B1(n_317),
.B2(n_313),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_369),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_415),
.B(n_417),
.Y(n_438)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_368),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_365),
.A2(n_387),
.B1(n_346),
.B2(n_362),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_379),
.A2(n_307),
.B1(n_320),
.B2(n_336),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_374),
.A2(n_335),
.B1(n_305),
.B2(n_340),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_349),
.B(n_265),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_349),
.B(n_261),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_265),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_426),
.B(n_306),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_390),
.A2(n_388),
.B1(n_358),
.B2(n_382),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_429),
.A2(n_432),
.B1(n_440),
.B2(n_448),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_400),
.A2(n_377),
.B1(n_371),
.B2(n_363),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_433),
.A2(n_429),
.B1(n_437),
.B2(n_405),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_434),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_412),
.B(n_363),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_435),
.B(n_454),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_436),
.A2(n_444),
.B(n_405),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_418),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_443),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_419),
.A2(n_359),
.B1(n_378),
.B2(n_357),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_397),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_441),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_391),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_393),
.B(n_372),
.Y(n_445)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_445),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_393),
.B(n_410),
.Y(n_446)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_391),
.A2(n_359),
.B1(n_372),
.B2(n_357),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_391),
.A2(n_380),
.B1(n_383),
.B2(n_350),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_449),
.A2(n_450),
.B1(n_407),
.B2(n_396),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_420),
.A2(n_383),
.B1(n_350),
.B2(n_352),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_402),
.A2(n_264),
.B(n_338),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_452),
.A2(n_396),
.B(n_402),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_406),
.A2(n_306),
.B1(n_257),
.B2(n_261),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_457),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_455),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_389),
.Y(n_457)
);

XNOR2x2_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_392),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_399),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_394),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_463),
.A2(n_452),
.B(n_436),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_404),
.C(n_411),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_466),
.C(n_475),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_399),
.C(n_401),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_445),
.Y(n_468)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_470),
.A2(n_442),
.B1(n_430),
.B2(n_447),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_423),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g502 ( 
.A1(n_472),
.A2(n_449),
.B(n_448),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_425),
.C(n_409),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_422),
.Y(n_476)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_476),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_446),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_478),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_444),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_428),
.B(n_430),
.Y(n_479)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_479),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_438),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_480),
.B(n_439),
.Y(n_489)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_454),
.B(n_435),
.C(n_458),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_457),
.C(n_442),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_483),
.A2(n_487),
.B(n_433),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_392),
.Y(n_493)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_451),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_485),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_466),
.C(n_486),
.Y(n_512)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_489),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_475),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_494),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_492),
.A2(n_474),
.B(n_479),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_502),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_469),
.B(n_431),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_498),
.B(n_511),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_461),
.B(n_427),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_499),
.B(n_471),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_483),
.A2(n_427),
.B1(n_440),
.B2(n_432),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_501),
.A2(n_507),
.B1(n_465),
.B2(n_474),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_504),
.A2(n_510),
.B1(n_485),
.B2(n_481),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_486),
.B(n_395),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_508),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_462),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_477),
.A2(n_447),
.B1(n_450),
.B2(n_426),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_395),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_473),
.A2(n_453),
.B1(n_258),
.B2(n_271),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_464),
.B(n_259),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_521),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_491),
.Y(n_517)
);

BUFx24_ASAP7_75t_SL g533 ( 
.A(n_517),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_510),
.A2(n_467),
.B1(n_468),
.B2(n_465),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_520),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_478),
.C(n_472),
.Y(n_520)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_522),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_500),
.B(n_472),
.C(n_487),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_528),
.C(n_252),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_506),
.B(n_461),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_524),
.B(n_526),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_462),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_525),
.B(n_247),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_496),
.B(n_467),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_527),
.A2(n_490),
.B1(n_497),
.B2(n_504),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_488),
.B(n_484),
.C(n_463),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_529),
.A2(n_502),
.B(n_509),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_530),
.A2(n_503),
.B1(n_495),
.B2(n_471),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_SL g549 ( 
.A(n_531),
.B(n_542),
.C(n_516),
.Y(n_549)
);

OAI321xp33_ASAP7_75t_L g532 ( 
.A1(n_519),
.A2(n_490),
.A3(n_509),
.B1(n_497),
.B2(n_476),
.C(n_503),
.Y(n_532)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_532),
.Y(n_547)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_535),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_538),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_SL g538 ( 
.A1(n_525),
.A2(n_492),
.B1(n_493),
.B2(n_505),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_513),
.A2(n_508),
.B1(n_258),
.B2(n_259),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_514),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_515),
.A2(n_247),
.B1(n_252),
.B2(n_277),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_540),
.A2(n_543),
.B1(n_16),
.B2(n_14),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_541),
.B(n_545),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_523),
.A2(n_520),
.B(n_528),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_515),
.A2(n_516),
.B1(n_514),
.B2(n_521),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_548),
.B(n_549),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_512),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_550),
.B(n_556),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_544),
.A2(n_277),
.B(n_15),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_551),
.A2(n_554),
.B(n_555),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_L g554 ( 
.A(n_534),
.B(n_277),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_537),
.B(n_14),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_537),
.B(n_14),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_557),
.A2(n_545),
.B1(n_531),
.B2(n_540),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_547),
.B(n_533),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_562),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_536),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_551),
.Y(n_563)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_563),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_564),
.A2(n_553),
.B(n_543),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_567),
.B(n_568),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_560),
.A2(n_553),
.B(n_561),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_565),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_570),
.B(n_572),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_566),
.B(n_558),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_571),
.A2(n_557),
.B(n_558),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_541),
.B(n_15),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_575),
.A2(n_573),
.B(n_15),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_576),
.B(n_15),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_577),
.B(n_16),
.Y(n_578)
);


endmodule