module fake_jpeg_19332_n_155 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_30),
.B(n_10),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_15),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_76),
.Y(n_82)
);

INVx11_ASAP7_75t_SL g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_80),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_65),
.B1(n_68),
.B2(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_52),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_88),
.C(n_72),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_65),
.B1(n_54),
.B2(n_47),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_87),
.B1(n_91),
.B2(n_53),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_66),
.B1(n_59),
.B2(n_71),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_66),
.B1(n_72),
.B2(n_70),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_73),
.B1(n_64),
.B2(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_105),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_90),
.B1(n_88),
.B2(n_51),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_89),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_84),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_116),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_117),
.B1(n_67),
.B2(n_3),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_50),
.B1(n_69),
.B2(n_57),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_5),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_96),
.B1(n_103),
.B2(n_104),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

AO21x2_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_62),
.B(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_7),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_63),
.C(n_62),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_7),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_16),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_132),
.B(n_20),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_6),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_8),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_28),
.B1(n_43),
.B2(n_42),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_118),
.B(n_115),
.Y(n_134)
);

OAI211xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_25),
.B(n_40),
.C(n_39),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_119),
.B(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_135),
.A2(n_139),
.B1(n_127),
.B2(n_130),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_138),
.C(n_8),
.Y(n_144)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_135),
.C(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_133),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_143),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_14),
.B1(n_38),
.B2(n_33),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_29),
.B(n_46),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_9),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_9),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_11),
.Y(n_155)
);


endmodule