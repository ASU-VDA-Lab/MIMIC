module fake_jpeg_27693_n_356 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_34),
.Y(n_60)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_27),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_17),
.B(n_32),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_57),
.A2(n_17),
.B1(n_49),
.B2(n_29),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_18),
.B1(n_19),
.B2(n_26),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_61),
.B1(n_75),
.B2(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_60),
.B(n_62),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_18),
.B1(n_19),
.B2(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_72),
.Y(n_93)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_74),
.B(n_83),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_33),
.B1(n_30),
.B2(n_27),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_84),
.B1(n_49),
.B2(n_17),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_33),
.B1(n_35),
.B2(n_23),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_35),
.B1(n_17),
.B2(n_32),
.Y(n_107)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_82),
.Y(n_109)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_33),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_27),
.B1(n_32),
.B2(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_11),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_31),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_48),
.B(n_42),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_106),
.B1(n_119),
.B2(n_101),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_47),
.B(n_42),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_92),
.A2(n_110),
.B(n_117),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_99),
.Y(n_153)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_47),
.B1(n_50),
.B2(n_32),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_39),
.B1(n_35),
.B2(n_51),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_97),
.A2(n_107),
.B1(n_79),
.B2(n_82),
.Y(n_144)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_98),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_118),
.Y(n_141)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_113),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_104),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_31),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_35),
.B1(n_29),
.B2(n_21),
.Y(n_106)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_88),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_67),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_49),
.C(n_68),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_64),
.B(n_29),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_64),
.A2(n_49),
.B(n_15),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_21),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_125),
.Y(n_129)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_21),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_134),
.A2(n_144),
.B1(n_78),
.B2(n_65),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_136),
.B(n_151),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_111),
.B(n_97),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_142),
.Y(n_160)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_139),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_83),
.Y(n_142)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_62),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_147),
.Y(n_174)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_102),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_60),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_87),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_87),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_116),
.C(n_126),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_100),
.A2(n_95),
.B1(n_107),
.B2(n_120),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_158),
.A2(n_110),
.B1(n_117),
.B2(n_106),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_163),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_156),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_184),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_170),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_175),
.B1(n_193),
.B2(n_153),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_13),
.B(n_14),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_123),
.B1(n_122),
.B2(n_94),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_185),
.B1(n_189),
.B2(n_191),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_118),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_85),
.CI(n_71),
.CON(n_171),
.SN(n_171)
);

XOR2x2_ASAP7_75t_SL g217 ( 
.A(n_171),
.B(n_36),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_115),
.B(n_91),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_173),
.A2(n_180),
.B(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_137),
.A2(n_85),
.B1(n_86),
.B2(n_81),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_178),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_96),
.Y(n_179)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_65),
.B(n_66),
.C(n_69),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_181),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_108),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_127),
.C(n_115),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_195),
.C(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_132),
.B(n_91),
.Y(n_198)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_124),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_138),
.Y(n_207)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_133),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_36),
.C(n_127),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_197),
.A2(n_209),
.B(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_207),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_164),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_129),
.B1(n_128),
.B2(n_147),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_201),
.A2(n_203),
.B1(n_205),
.B2(n_216),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_175),
.B1(n_183),
.B2(n_167),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_211),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_167),
.A2(n_129),
.B1(n_142),
.B2(n_138),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_155),
.C(n_154),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_208),
.B(n_212),
.C(n_143),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_130),
.B(n_146),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_135),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_152),
.C(n_130),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_165),
.A2(n_150),
.B1(n_139),
.B2(n_70),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_180),
.B(n_194),
.C(n_161),
.D(n_163),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_177),
.A2(n_1),
.B(n_2),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_12),
.B(n_14),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_152),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_227),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_176),
.A2(n_150),
.B1(n_82),
.B2(n_79),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_176),
.B1(n_186),
.B2(n_188),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_121),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_226),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_185),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g225 ( 
.A1(n_171),
.A2(n_150),
.B1(n_121),
.B2(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_79),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_160),
.B(n_190),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_161),
.B1(n_215),
.B2(n_222),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_257),
.B1(n_218),
.B2(n_196),
.Y(n_271)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_199),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_243),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_228),
.B(n_178),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_237),
.B(n_238),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_240),
.B(n_12),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_214),
.B1(n_205),
.B2(n_217),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_191),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_253),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_162),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_193),
.Y(n_250)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_210),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_189),
.Y(n_252)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_224),
.B(n_13),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_255),
.A2(n_200),
.B1(n_203),
.B2(n_225),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_208),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_172),
.C(n_13),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_256),
.C(n_269),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_260),
.A2(n_267),
.B1(n_269),
.B2(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_197),
.B1(n_209),
.B2(n_206),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_226),
.B1(n_204),
.B2(n_212),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_232),
.A2(n_207),
.B1(n_211),
.B2(n_223),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_276),
.B1(n_279),
.B2(n_230),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_232),
.A2(n_172),
.B1(n_143),
.B2(n_5),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_253),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_278),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_242),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_284),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_268),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_250),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_233),
.C(n_239),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_289),
.C(n_292),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_233),
.C(n_239),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_242),
.B(n_230),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_298),
.B(n_275),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_235),
.C(n_245),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_295),
.B(n_296),
.Y(n_306)
);

BUFx12_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_231),
.B(n_245),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_235),
.C(n_252),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_299),
.B(n_301),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_248),
.B1(n_246),
.B2(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_265),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_312),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_258),
.B(n_266),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_309),
.B(n_314),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_294),
.A2(n_267),
.B(n_260),
.Y(n_309)
);

XNOR2x1_ASAP7_75t_SL g310 ( 
.A(n_291),
.B(n_295),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_310),
.B(n_313),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_298),
.Y(n_328)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_262),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_288),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_284),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_319),
.A2(n_3),
.B(n_6),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_290),
.B1(n_282),
.B2(n_261),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_330),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_285),
.C(n_287),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_327),
.C(n_328),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_319),
.B(n_264),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_290),
.B1(n_307),
.B2(n_297),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_326),
.A2(n_329),
.B1(n_313),
.B2(n_302),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_289),
.C(n_292),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_303),
.A2(n_264),
.B1(n_263),
.B2(n_270),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_280),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_302),
.B1(n_314),
.B2(n_312),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_333),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_334),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_323),
.A2(n_315),
.B1(n_306),
.B2(n_309),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_320),
.A2(n_240),
.B1(n_276),
.B2(n_277),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_336),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_324),
.B(n_7),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_3),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_338),
.B(n_340),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_330),
.B(n_3),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_342),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_335),
.A2(n_339),
.B(n_331),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_324),
.B(n_327),
.Y(n_346)
);

AOI322xp5_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_322),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_6),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_SL g348 ( 
.A1(n_343),
.A2(n_336),
.B(n_337),
.C(n_339),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

AOI322xp5_ASAP7_75t_L g352 ( 
.A1(n_349),
.A2(n_351),
.A3(n_344),
.B1(n_345),
.B2(n_7),
.C1(n_10),
.C2(n_347),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_343),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_351)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_352),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_350),
.B(n_353),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_10),
.Y(n_356)
);


endmodule