module fake_jpeg_11279_n_143 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_42),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_9),
.B(n_44),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_2),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_22),
.B1(n_38),
.B2(n_37),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_52),
.B1(n_46),
.B2(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_4),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_61),
.B(n_53),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_94),
.B(n_8),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_55),
.B(n_59),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_23),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_60),
.B(n_56),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_64),
.B1(n_59),
.B2(n_55),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_63),
.B1(n_9),
.B2(n_10),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_63),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_63),
.B1(n_5),
.B2(n_7),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_102),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_4),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_118),
.B1(n_29),
.B2(n_30),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_24),
.C(n_11),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_40),
.C(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_25),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_115),
.B(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_91),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_12),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_13),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_15),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_16),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_123),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_127),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_128),
.Y(n_132)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_133),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_SL g137 ( 
.A(n_131),
.B(n_106),
.C(n_122),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_138),
.B1(n_108),
.B2(n_135),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_122),
.B(n_116),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_136),
.B(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g142 ( 
.A(n_141),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_132),
.Y(n_143)
);


endmodule