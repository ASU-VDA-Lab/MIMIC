module fake_jpeg_28867_n_321 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_49),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_13),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_0),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_21),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_56),
.B(n_96),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_16),
.B1(n_35),
.B2(n_20),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_57),
.A2(n_91),
.B1(n_92),
.B2(n_24),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_21),
.B1(n_22),
.B2(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_58),
.A2(n_69),
.B1(n_73),
.B2(n_80),
.Y(n_135)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_54),
.B1(n_46),
.B2(n_35),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_22),
.B1(n_31),
.B2(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_77),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_31),
.B1(n_23),
.B2(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_37),
.B(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_26),
.Y(n_83)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_43),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_10),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_35),
.B1(n_20),
.B2(n_32),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_27),
.B1(n_25),
.B2(n_19),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_43),
.B(n_34),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_34),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_39),
.A2(n_31),
.B1(n_19),
.B2(n_27),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_32),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_25),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_45),
.A2(n_27),
.B1(n_25),
.B2(n_19),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_SL g105 ( 
.A(n_68),
.B(n_26),
.C(n_24),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_121),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_17),
.B1(n_28),
.B2(n_25),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_123),
.B1(n_129),
.B2(n_130),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_17),
.B(n_9),
.C(n_13),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_5),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_133),
.B1(n_134),
.B2(n_6),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_28),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_61),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_28),
.B(n_24),
.C(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_72),
.B(n_28),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_90),
.B(n_28),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_131),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_62),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_5),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_134),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_70),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_103),
.B(n_90),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_140),
.B(n_151),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_56),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_147),
.C(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_132),
.B1(n_130),
.B2(n_133),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_56),
.C(n_85),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_76),
.C(n_86),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_76),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_85),
.C(n_61),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_70),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_96),
.B(n_95),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_161),
.B(n_66),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_86),
.C(n_93),
.Y(n_158)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_112),
.A2(n_63),
.B(n_71),
.Y(n_161)
);

BUFx4f_ASAP7_75t_SL g162 ( 
.A(n_122),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_67),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_104),
.B(n_67),
.Y(n_164)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_167),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_63),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_170),
.Y(n_198)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_111),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_120),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_195),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_115),
.B1(n_129),
.B2(n_118),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_196),
.B1(n_203),
.B2(n_150),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_120),
.C(n_115),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_200),
.C(n_206),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_192),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_193),
.A2(n_199),
.B(n_143),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_120),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_120),
.B(n_130),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_130),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_138),
.B(n_122),
.C(n_123),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_159),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_202),
.B(n_204),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_157),
.A2(n_111),
.B1(n_59),
.B2(n_87),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_111),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_147),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_109),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_145),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_207),
.Y(n_213)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_210),
.A2(n_126),
.B(n_108),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_219),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_227),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_148),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_222),
.C(n_182),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_150),
.B1(n_158),
.B2(n_141),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_168),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_150),
.B1(n_171),
.B2(n_152),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_226),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_228),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_192),
.A2(n_175),
.B1(n_203),
.B2(n_181),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_178),
.B1(n_198),
.B2(n_206),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_172),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_169),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_236),
.Y(n_255)
);

NOR2x1_ASAP7_75t_R g235 ( 
.A(n_201),
.B(n_165),
.Y(n_235)
);

AOI221xp5_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_184),
.B1(n_180),
.B2(n_190),
.C(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

AOI211xp5_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_197),
.B(n_178),
.C(n_180),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_239),
.B1(n_226),
.B2(n_229),
.Y(n_261)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_184),
.B1(n_188),
.B2(n_177),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_247),
.C(n_252),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_253),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_185),
.A3(n_191),
.B1(n_183),
.B2(n_188),
.C1(n_208),
.C2(n_189),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_254),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_183),
.C(n_208),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_174),
.C(n_189),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_223),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_160),
.C(n_177),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_109),
.C(n_108),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_215),
.B(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_213),
.B(n_6),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_257),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_224),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_264),
.B1(n_267),
.B2(n_275),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_230),
.B1(n_227),
.B2(n_212),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_228),
.B1(n_225),
.B2(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_270),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_219),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_214),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_272),
.A2(n_274),
.B1(n_257),
.B2(n_250),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_276),
.Y(n_283)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_232),
.B1(n_214),
.B2(n_101),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_6),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_247),
.C(n_252),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_241),
.C(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_238),
.C(n_244),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_284),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_238),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_261),
.A2(n_259),
.B1(n_258),
.B2(n_254),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_285),
.A2(n_264),
.B1(n_275),
.B2(n_240),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_244),
.C(n_246),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_262),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_296),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_295),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_268),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_294),
.C(n_281),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_265),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_273),
.B1(n_237),
.B2(n_255),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_239),
.B(n_267),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_305),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_289),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_300),
.B(n_293),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_290),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_SL g307 ( 
.A1(n_291),
.A2(n_239),
.B(n_282),
.C(n_287),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_278),
.C(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_306),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_250),
.B1(n_295),
.B2(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_313),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_307),
.B(n_74),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_304),
.C(n_303),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_316),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_311),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_311),
.C(n_65),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_318),
.B(n_74),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_98),
.Y(n_321)
);


endmodule