module fake_jpeg_25359_n_356 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_40),
.B(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_41),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_51),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_55),
.Y(n_75)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_58),
.Y(n_86)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_0),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_62),
.B1(n_80),
.B2(n_97),
.Y(n_100)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_74),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_85),
.B1(n_96),
.B2(n_81),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_66),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_67),
.Y(n_128)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_72),
.B(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_87),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_23),
.B1(n_26),
.B2(n_20),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_25),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_39),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_42),
.B(n_34),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_89),
.B(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_19),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_37),
.B1(n_28),
.B2(n_32),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_19),
.B1(n_36),
.B2(n_32),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_62),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_111),
.C(n_118),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_57),
.B1(n_37),
.B2(n_32),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_103),
.A2(n_107),
.B1(n_123),
.B2(n_22),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_119),
.Y(n_149)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_57),
.B1(n_37),
.B2(n_32),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_45),
.B1(n_44),
.B2(n_28),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_108),
.A2(n_135),
.B1(n_60),
.B2(n_61),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_92),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_55),
.C(n_18),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_51),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_125),
.Y(n_148)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_114),
.B(n_132),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_45),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_1),
.B(n_2),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_1),
.B(n_2),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_71),
.A2(n_36),
.B1(n_19),
.B2(n_28),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_126),
.Y(n_168)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_36),
.B1(n_37),
.B2(n_13),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_44),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_34),
.B1(n_22),
.B2(n_18),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_34),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_134),
.Y(n_150)
);

BUFx10_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_73),
.B(n_35),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_34),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_95),
.A2(n_93),
.B1(n_18),
.B2(n_22),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_33),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_83),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_2),
.B(n_3),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_167),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_83),
.B1(n_70),
.B2(n_69),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_35),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_130),
.C(n_137),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_152),
.Y(n_173)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_154),
.Y(n_172)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_158),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_73),
.B1(n_22),
.B2(n_35),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_160),
.B1(n_165),
.B2(n_118),
.Y(n_175)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_163),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_12),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_100),
.B1(n_120),
.B2(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_33),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_33),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_102),
.A2(n_77),
.B1(n_35),
.B2(n_33),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_100),
.B1(n_121),
.B2(n_111),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_116),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_163),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_175),
.A2(n_195),
.B(n_201),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_184),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_102),
.B1(n_122),
.B2(n_124),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_138),
.B1(n_126),
.B2(n_117),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_126),
.B1(n_115),
.B2(n_101),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_128),
.B1(n_142),
.B2(n_101),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_126),
.B1(n_128),
.B2(n_106),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_193),
.B1(n_202),
.B2(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_192),
.Y(n_214)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_205),
.Y(n_225)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_189),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_168),
.B(n_158),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_148),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_167),
.A2(n_77),
.B1(n_130),
.B2(n_136),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_137),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_136),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_204),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_146),
.Y(n_210)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_200),
.B(n_203),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_130),
.B(n_4),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_171),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_140),
.B(n_3),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_155),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_143),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_147),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_211),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_147),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_149),
.C(n_161),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_213),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_149),
.C(n_168),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_216),
.B(n_217),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_4),
.B(n_142),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_190),
.B(n_178),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_151),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_221),
.B(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_180),
.B(n_151),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_154),
.A3(n_153),
.B1(n_8),
.B2(n_10),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_239),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_162),
.B1(n_7),
.B2(n_8),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_176),
.B1(n_173),
.B2(n_188),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_162),
.C(n_11),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_236),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_174),
.A2(n_6),
.B(n_11),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_232),
.Y(n_251)
);

A2O1A1O1Ixp25_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_6),
.B(n_13),
.C(n_14),
.D(n_15),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_191),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_174),
.A2(n_14),
.B(n_15),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_240),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_254),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_233),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_250),
.A2(n_253),
.B(n_256),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_264),
.C(n_232),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_187),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_260),
.Y(n_270)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_261),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_219),
.A2(n_175),
.B1(n_186),
.B2(n_179),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_184),
.B1(n_219),
.B2(n_226),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_216),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_182),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_265),
.Y(n_286)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_209),
.C(n_213),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_279),
.C(n_280),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_210),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_269),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_227),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_227),
.B(n_238),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_275),
.B1(n_254),
.B2(n_243),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_212),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_278),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_247),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_220),
.C(n_234),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_234),
.C(n_217),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_252),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_215),
.B(n_240),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_255),
.C(n_242),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_242),
.A2(n_238),
.B(n_231),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_251),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_236),
.C(n_207),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_224),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_261),
.C(n_265),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_299),
.C(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_293),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_292),
.B1(n_304),
.B2(n_281),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_274),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_244),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_263),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_224),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_303),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_259),
.C(n_248),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_272),
.A2(n_243),
.B1(n_249),
.B2(n_266),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_302),
.B1(n_283),
.B2(n_251),
.Y(n_314)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_255),
.B1(n_286),
.B2(n_259),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_273),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_306),
.B(n_315),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_278),
.C(n_269),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_319),
.C(n_315),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_299),
.C(n_301),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_313),
.Y(n_330)
);

A2O1A1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_271),
.B(n_287),
.C(n_280),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_257),
.B(n_241),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_253),
.Y(n_324)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_305),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_285),
.C(n_250),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_320),
.A2(n_307),
.B1(n_308),
.B2(n_316),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_293),
.B1(n_288),
.B2(n_296),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_294),
.B1(n_270),
.B2(n_256),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_257),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_327),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_260),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_199),
.B(n_189),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_241),
.Y(n_327)
);

INVx11_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_202),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_181),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_329),
.B(n_14),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_294),
.B(n_206),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_336),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_333),
.A2(n_334),
.B(n_339),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_338),
.B(n_340),
.C(n_324),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_326),
.A2(n_260),
.B(n_199),
.Y(n_336)
);

AOI322xp5_ASAP7_75t_L g350 ( 
.A1(n_343),
.A2(n_16),
.A3(n_196),
.B1(n_323),
.B2(n_325),
.C1(n_344),
.C2(n_342),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_335),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_344),
.A2(n_345),
.B(n_196),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_339),
.A2(n_330),
.B(n_321),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_337),
.B(n_331),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_347),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_323),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_328),
.C(n_325),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_351),
.C(n_16),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_350),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_352),
.A2(n_349),
.B(n_16),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_353),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_355),
.Y(n_356)
);


endmodule