module fake_jpeg_17053_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVxp33_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_29),
.Y(n_56)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_59),
.B(n_62),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_61),
.B(n_29),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_66),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_37),
.B1(n_28),
.B2(n_35),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_35),
.B1(n_28),
.B2(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_53),
.B1(n_23),
.B2(n_27),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_84),
.A2(n_88),
.B1(n_96),
.B2(n_44),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_82),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_93),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_28),
.B1(n_51),
.B2(n_23),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_110),
.B1(n_75),
.B2(n_50),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_51),
.B1(n_53),
.B2(n_32),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g89 ( 
.A(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_51),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_27),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_81),
.B1(n_77),
.B2(n_75),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_67),
.B1(n_83),
.B2(n_63),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_27),
.A3(n_17),
.B1(n_39),
.B2(n_36),
.Y(n_97)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_24),
.A3(n_26),
.B1(n_22),
.B2(n_25),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_34),
.C(n_32),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_50),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_66),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_32),
.B1(n_38),
.B2(n_36),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_67),
.A2(n_27),
.B1(n_16),
.B2(n_18),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_117),
.A2(n_135),
.B(n_95),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_134),
.B(n_107),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_85),
.B(n_16),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_130),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_129),
.B1(n_137),
.B2(n_88),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_103),
.B1(n_95),
.B2(n_109),
.Y(n_158)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_18),
.B1(n_24),
.B2(n_26),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_50),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_94),
.A2(n_26),
.B1(n_24),
.B2(n_22),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_44),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_44),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_139),
.B(n_107),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_105),
.CI(n_102),
.CON(n_140),
.SN(n_140)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_145),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_151),
.B1(n_157),
.B2(n_167),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_111),
.C(n_96),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_160),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_104),
.B(n_25),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_117),
.A2(n_96),
.B1(n_101),
.B2(n_100),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_120),
.C(n_128),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_164),
.C(n_170),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_165),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_108),
.B(n_103),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_163),
.B(n_171),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_96),
.B1(n_101),
.B2(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_169),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_25),
.B(n_21),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_104),
.C(n_38),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_34),
.B1(n_98),
.B2(n_19),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_127),
.B1(n_14),
.B2(n_13),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_11),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_25),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_21),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_185),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_180),
.B1(n_184),
.B2(n_204),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_160),
.B(n_147),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_188),
.B(n_203),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_114),
.B1(n_122),
.B2(n_125),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_170),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_202),
.C(n_21),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_114),
.B1(n_126),
.B2(n_124),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_131),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_189),
.B(n_195),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_162),
.B1(n_166),
.B2(n_143),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_104),
.Y(n_192)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_21),
.Y(n_193)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_150),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_150),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_198),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_155),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_140),
.C(n_113),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_26),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_113),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_0),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_1),
.B(n_2),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_157),
.B1(n_168),
.B2(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_158),
.B1(n_171),
.B2(n_143),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_224),
.B(n_204),
.C(n_175),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_167),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_218),
.C(n_221),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_177),
.A2(n_30),
.B1(n_19),
.B2(n_24),
.Y(n_216)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_174),
.A2(n_181),
.B1(n_186),
.B2(n_176),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_219),
.B(n_30),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_21),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_178),
.C(n_202),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_192),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_174),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_178),
.B(n_22),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_194),
.Y(n_234)
);

FAx1_ASAP7_75t_SL g231 ( 
.A(n_221),
.B(n_194),
.CI(n_203),
.CON(n_231),
.SN(n_231)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_183),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_239),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_251),
.B1(n_224),
.B2(n_212),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_234),
.B(n_250),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_188),
.B(n_203),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_246),
.B(n_214),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_180),
.B(n_172),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_236),
.A2(n_247),
.B1(n_235),
.B2(n_242),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_244),
.B1(n_248),
.B2(n_208),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_241),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_219),
.Y(n_261)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_217),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_187),
.B1(n_181),
.B2(n_201),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_193),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_226),
.C(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_261),
.C(n_264),
.Y(n_271)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_231),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_213),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_266),
.C(n_3),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_30),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_236),
.A2(n_223),
.B1(n_215),
.B2(n_248),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_262),
.A2(n_265),
.B1(n_233),
.B2(n_2),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_211),
.B1(n_225),
.B2(n_206),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_263),
.A2(n_233),
.B1(n_248),
.B2(n_210),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_207),
.C(n_216),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_210),
.B1(n_30),
.B2(n_19),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_234),
.C(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_275),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g274 ( 
.A(n_254),
.B(n_233),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_260),
.B1(n_262),
.B2(n_268),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_12),
.C(n_10),
.Y(n_278)
);

BUFx12f_ASAP7_75t_SL g290 ( 
.A(n_278),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_282),
.Y(n_295)
);

FAx1_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_1),
.CI(n_2),
.CON(n_280),
.SN(n_280)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_281),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_21),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_3),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_266),
.C(n_264),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_271),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_259),
.C(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_9),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_265),
.B1(n_255),
.B2(n_6),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_276),
.B1(n_277),
.B2(n_280),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_301),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_274),
.B(n_283),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_305),
.B(n_293),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_304),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_280),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_302),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_4),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_303),
.Y(n_311)
);

XNOR2x1_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_4),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_306),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_291),
.B(n_290),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_295),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_295),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_312),
.B(n_305),
.C(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_314),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_313),
.B(n_307),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_309),
.B(n_284),
.Y(n_319)
);

OAI221xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_288),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_7),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_8),
.B(n_302),
.Y(n_323)
);


endmodule