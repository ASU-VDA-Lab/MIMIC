module fake_netlist_5_264_n_935 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_935);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_935;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_284;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_433;
wire n_368;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_624;
wire n_252;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_929;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_399;
wire n_341;
wire n_394;
wire n_204;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_795;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_917;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_513;
wire n_425;
wire n_407;
wire n_527;
wire n_707;
wire n_679;
wire n_710;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_868;
wire n_803;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_927;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

INVx2_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_111),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_60),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_31),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_30),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_18),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_51),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_54),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_31),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_63),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_58),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_97),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_13),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_8),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_70),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_47),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_179),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_28),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_181),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_35),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_130),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_62),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_15),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_112),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_14),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_28),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_90),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_34),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_106),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_48),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_133),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_88),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_87),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_25),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_43),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_143),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_153),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_177),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_37),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_144),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_10),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_93),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_119),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_21),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_59),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_23),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_183),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_56),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_77),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_91),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_98),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_3),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_20),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_84),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_1),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_20),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_105),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_26),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_32),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_109),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_178),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_167),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_115),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_44),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_141),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_37),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_34),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_120),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_81),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_36),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_13),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_149),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_180),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_24),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_139),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_35),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_22),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_184),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_127),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_50),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_107),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_225),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_0),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_190),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_209),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_229),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_229),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_210),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_229),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_194),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_198),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_193),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_215),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_220),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_226),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_198),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_212),
.B(n_0),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_193),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_195),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_195),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_200),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_230),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_217),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_232),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_233),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_238),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_217),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_240),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_218),
.B(n_2),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_207),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_219),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_222),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_227),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_236),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_244),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_255),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_265),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_222),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_250),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_239),
.B(n_2),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_214),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_247),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_250),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_267),
.Y(n_335)
);

BUFx2_ASAP7_75t_SL g336 ( 
.A(n_242),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_249),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_259),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_273),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_245),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_234),
.B(n_3),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_241),
.B(n_4),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_260),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_271),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_272),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_275),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_274),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_245),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_277),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_279),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_191),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_292),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_293),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_304),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_300),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_298),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_301),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_309),
.B(n_188),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_300),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_332),
.B(n_246),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_307),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_305),
.B(n_191),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_287),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_337),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_310),
.B(n_311),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_302),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_306),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_313),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_315),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_299),
.A2(n_263),
.B1(n_256),
.B2(n_282),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_307),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_316),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_196),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_317),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_319),
.B(n_196),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_213),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_299),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_291),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_326),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_331),
.B(n_231),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_320),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_328),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_308),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_359),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_360),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_364),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_394),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_364),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_354),
.Y(n_421)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_383),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_408),
.B(n_234),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_408),
.B(n_383),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_410),
.A2(n_350),
.B1(n_347),
.B2(n_216),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_290),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_408),
.B(n_248),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_231),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_389),
.Y(n_433)
);

AO21x2_ASAP7_75t_L g434 ( 
.A1(n_391),
.A2(n_192),
.B(n_189),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_286),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_383),
.Y(n_437)
);

AND2x6_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_248),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_404),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_365),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_394),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_354),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_411),
.B(n_197),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_278),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_389),
.B(n_199),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_405),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_358),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_401),
.B(n_294),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_386),
.B(n_327),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_374),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_358),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_361),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_410),
.B(n_202),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_407),
.B(n_204),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_206),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_407),
.B(n_211),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_357),
.B(n_340),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_401),
.A2(n_188),
.B1(n_208),
.B2(n_223),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_266),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_361),
.B(n_224),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_361),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_361),
.Y(n_469)
);

NAND2x1p5_ASAP7_75t_L g470 ( 
.A(n_367),
.B(n_228),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_369),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g472 ( 
.A(n_384),
.B(n_208),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_403),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_366),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_366),
.B(n_235),
.Y(n_475)
);

NAND2x1p5_ASAP7_75t_L g476 ( 
.A(n_367),
.B(n_237),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_372),
.A2(n_349),
.B1(n_340),
.B2(n_201),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_369),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_376),
.Y(n_479)
);

NAND2x1p5_ASAP7_75t_L g480 ( 
.A(n_376),
.B(n_251),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_378),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_370),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_362),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_421),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_472),
.B(n_355),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_430),
.B(n_356),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_472),
.B(n_382),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_462),
.A2(n_466),
.B1(n_433),
.B2(n_464),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_412),
.B(n_385),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_428),
.B(n_390),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_403),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_474),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_423),
.A2(n_253),
.B1(n_257),
.B2(n_268),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_479),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_421),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_413),
.B(n_406),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_426),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_433),
.B(n_409),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_426),
.Y(n_500)
);

NOR2x2_ASAP7_75t_L g501 ( 
.A(n_436),
.B(n_314),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_417),
.B(n_420),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_447),
.B(n_388),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_445),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_449),
.B(n_443),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_415),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_429),
.B(n_377),
.Y(n_507)
);

INVx8_ASAP7_75t_L g508 ( 
.A(n_447),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_L g509 ( 
.A(n_447),
.B(n_201),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_473),
.B(n_377),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_471),
.Y(n_511)
);

O2A1O1Ixp5_ASAP7_75t_L g512 ( 
.A1(n_423),
.A2(n_280),
.B(n_261),
.C(n_399),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_432),
.B(n_378),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_433),
.B(n_381),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_457),
.Y(n_515)
);

NAND2x1p5_ASAP7_75t_L g516 ( 
.A(n_414),
.B(n_379),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_414),
.B(n_379),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_455),
.B(n_349),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_456),
.B(n_392),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_446),
.B(n_455),
.Y(n_521)
);

A2O1A1Ixp33_ASAP7_75t_L g522 ( 
.A1(n_462),
.A2(n_396),
.B(n_392),
.C(n_399),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_478),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_478),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_456),
.B(n_440),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_429),
.B(n_395),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_458),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_458),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_446),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_452),
.B(n_395),
.Y(n_531)
);

OAI221xp5_ASAP7_75t_L g532 ( 
.A1(n_465),
.A2(n_397),
.B1(n_396),
.B2(n_400),
.C(n_393),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_469),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_427),
.A2(n_397),
.B(n_371),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_418),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_418),
.B(n_370),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_431),
.B(n_371),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_462),
.B(n_393),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_451),
.A2(n_447),
.B1(n_461),
.B2(n_463),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_450),
.B(n_400),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_471),
.B(n_381),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_477),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_482),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_447),
.A2(n_314),
.B1(n_318),
.B2(n_323),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_454),
.B(n_203),
.Y(n_546)
);

OAI22x1_ASAP7_75t_SL g547 ( 
.A1(n_436),
.A2(n_330),
.B1(n_318),
.B2(n_323),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_450),
.B(n_482),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_482),
.B(n_475),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_471),
.B(n_381),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_203),
.Y(n_551)
);

AND3x1_ASAP7_75t_L g552 ( 
.A(n_467),
.B(n_402),
.C(n_330),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_450),
.B(n_205),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_484),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_528),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_492),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_483),
.B(n_461),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_486),
.B(n_460),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_492),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_506),
.B(n_463),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_484),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_488),
.A2(n_447),
.B1(n_434),
.B2(n_427),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_513),
.B(n_431),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_SL g565 ( 
.A(n_543),
.B(n_263),
.C(n_256),
.Y(n_565)
);

NOR3xp33_ASAP7_75t_SL g566 ( 
.A(n_515),
.B(n_487),
.C(n_485),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_511),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_528),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_548),
.B(n_444),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_520),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_511),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_491),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_529),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_541),
.B(n_434),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_529),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_496),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_516),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_533),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_520),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_498),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_R g582 ( 
.A(n_490),
.B(n_368),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_526),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_540),
.B(n_505),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_510),
.B(n_329),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_527),
.B(n_434),
.Y(n_586)
);

NOR3xp33_ASAP7_75t_SL g587 ( 
.A(n_490),
.B(n_243),
.C(n_221),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_R g588 ( 
.A(n_503),
.B(n_373),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_508),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_545),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_521),
.B(n_470),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_519),
.B(n_470),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_499),
.A2(n_538),
.B1(n_527),
.B2(n_494),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_495),
.B(n_476),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_518),
.B(n_476),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_502),
.B(n_425),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_547),
.B(n_387),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_551),
.A2(n_438),
.B1(n_453),
.B2(n_468),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_531),
.B(n_329),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_549),
.B(n_489),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_531),
.B(n_439),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_520),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_535),
.B(n_471),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_551),
.B(n_441),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_526),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_539),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_542),
.B(n_550),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_507),
.B(n_334),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_558),
.B(n_497),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_567),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_558),
.B(n_553),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_602),
.B(n_526),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_570),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_606),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_560),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_567),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_584),
.A2(n_444),
.B(n_437),
.Y(n_621)
);

AO32x2_ASAP7_75t_L g622 ( 
.A1(n_609),
.A2(n_444),
.A3(n_437),
.B1(n_501),
.B2(n_534),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_566),
.B(n_546),
.C(n_381),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_604),
.B(n_546),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_584),
.A2(n_437),
.B(n_499),
.Y(n_625)
);

AO21x1_ASAP7_75t_L g626 ( 
.A1(n_586),
.A2(n_550),
.B(n_542),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_574),
.A2(n_536),
.B(n_525),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_572),
.B(n_580),
.Y(n_628)
);

AOI21x1_ASAP7_75t_SL g629 ( 
.A1(n_611),
.A2(n_517),
.B(n_512),
.Y(n_629)
);

AO31x2_ASAP7_75t_L g630 ( 
.A1(n_564),
.A2(n_522),
.A3(n_500),
.B(n_504),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_590),
.B(n_493),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_573),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_585),
.B(n_514),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g634 ( 
.A1(n_569),
.A2(n_555),
.B(n_562),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_567),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_556),
.B(n_559),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_569),
.A2(n_555),
.B(n_554),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_555),
.A2(n_537),
.B(n_516),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_554),
.A2(n_537),
.B(n_500),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_612),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_611),
.B(n_498),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_557),
.A2(n_524),
.B(n_504),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

NOR2x1_ASAP7_75t_L g644 ( 
.A(n_594),
.B(n_514),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_603),
.A2(n_416),
.B(n_509),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_601),
.A2(n_524),
.B(n_523),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_603),
.A2(n_416),
.B(n_448),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_595),
.B(n_334),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_599),
.B(n_544),
.Y(n_649)
);

O2A1O1Ixp5_ASAP7_75t_L g650 ( 
.A1(n_608),
.A2(n_459),
.B(n_442),
.C(n_419),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_592),
.B(n_552),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_593),
.B(n_493),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_561),
.A2(n_424),
.B(n_419),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_583),
.Y(n_654)
);

AO22x2_ASAP7_75t_L g655 ( 
.A1(n_611),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_593),
.B(n_480),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_596),
.B(n_480),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_471),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_643),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_556),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_615),
.A2(n_601),
.B(n_577),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_643),
.Y(n_662)
);

NAND2x1_ASAP7_75t_L g663 ( 
.A(n_614),
.B(n_571),
.Y(n_663)
);

OAI222xp33_ASAP7_75t_L g664 ( 
.A1(n_648),
.A2(n_624),
.B1(n_633),
.B2(n_652),
.C1(n_600),
.C2(n_644),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_639),
.A2(n_578),
.B(n_576),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_614),
.Y(n_666)
);

OA21x2_ASAP7_75t_L g667 ( 
.A1(n_650),
.A2(n_579),
.B(n_575),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_632),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_619),
.B(n_556),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_642),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_653),
.A2(n_578),
.B(n_576),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_636),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_649),
.B(n_556),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_640),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_656),
.A2(n_559),
.B1(n_563),
.B2(n_571),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_620),
.Y(n_676)
);

CKINVDCx8_ASAP7_75t_R g677 ( 
.A(n_636),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_636),
.B(n_559),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_653),
.A2(n_581),
.B(n_589),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_616),
.B(n_654),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_641),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_622),
.B(n_581),
.Y(n_682)
);

AOI21x1_ASAP7_75t_L g683 ( 
.A1(n_627),
.A2(n_610),
.B(n_597),
.Y(n_683)
);

BUFx12f_ASAP7_75t_L g684 ( 
.A(n_617),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_641),
.Y(n_685)
);

OA21x2_ASAP7_75t_L g686 ( 
.A1(n_650),
.A2(n_532),
.B(n_607),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_634),
.A2(n_637),
.B(n_638),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_654),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_637),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_638),
.B(n_590),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_618),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_630),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_630),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_625),
.B(n_591),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_634),
.A2(n_568),
.B(n_424),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_640),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_655),
.A2(n_582),
.B1(n_588),
.B2(n_612),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_620),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_657),
.A2(n_587),
.B(n_565),
.C(n_607),
.Y(n_699)
);

OAI221xp5_ASAP7_75t_L g700 ( 
.A1(n_623),
.A2(n_264),
.B1(n_582),
.B2(n_559),
.C(n_252),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_R g701 ( 
.A(n_674),
.B(n_588),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_688),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_660),
.B(n_658),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_659),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_697),
.A2(n_651),
.B1(n_655),
.B2(n_626),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_668),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_677),
.A2(n_655),
.B1(n_646),
.B2(n_635),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_664),
.A2(n_645),
.B(n_621),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_684),
.Y(n_709)
);

NOR2x1_ASAP7_75t_SL g710 ( 
.A(n_676),
.B(n_590),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_659),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_696),
.B(n_680),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_668),
.Y(n_713)
);

AOI221xp5_ASAP7_75t_L g714 ( 
.A1(n_700),
.A2(n_205),
.B1(n_252),
.B2(n_285),
.C(n_254),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_699),
.A2(n_631),
.B(n_628),
.C(n_647),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_681),
.A2(n_438),
.B1(n_242),
.B2(n_607),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_661),
.A2(n_631),
.B(n_635),
.C(n_568),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_674),
.A2(n_571),
.B1(n_254),
.B2(n_258),
.Y(n_718)
);

OAI221xp5_ASAP7_75t_L g719 ( 
.A1(n_688),
.A2(n_262),
.B1(n_285),
.B2(n_270),
.C(n_269),
.Y(n_719)
);

AO21x2_ASAP7_75t_L g720 ( 
.A1(n_683),
.A2(n_622),
.B(n_629),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_694),
.A2(n_605),
.B(n_590),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_673),
.B(n_438),
.Y(n_722)
);

AND2x2_ASAP7_75t_SL g723 ( 
.A(n_681),
.B(n_591),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_669),
.B(n_605),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_672),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_684),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_691),
.A2(n_270),
.B1(n_258),
.B2(n_262),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_678),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_677),
.A2(n_685),
.B1(n_676),
.B2(n_670),
.Y(n_729)
);

AOI211xp5_ASAP7_75t_L g730 ( 
.A1(n_675),
.A2(n_269),
.B(n_284),
.C(n_242),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_685),
.A2(n_605),
.B1(n_591),
.B2(n_622),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_678),
.B(n_284),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_691),
.A2(n_438),
.B1(n_605),
.B2(n_622),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_672),
.A2(n_629),
.B1(n_448),
.B2(n_424),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_678),
.B(n_438),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_678),
.Y(n_736)
);

AND2x2_ASAP7_75t_SL g737 ( 
.A(n_666),
.B(n_630),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_SL g738 ( 
.A1(n_670),
.A2(n_419),
.B(n_630),
.C(n_438),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_662),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_676),
.A2(n_448),
.B1(n_416),
.B2(n_422),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_662),
.B(n_5),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_698),
.B(n_6),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_698),
.B(n_7),
.Y(n_743)
);

CKINVDCx16_ASAP7_75t_R g744 ( 
.A(n_682),
.Y(n_744)
);

OAI221xp5_ASAP7_75t_L g745 ( 
.A1(n_694),
.A2(n_422),
.B1(n_448),
.B2(n_416),
.C(n_11),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_676),
.A2(n_448),
.B1(n_422),
.B2(n_416),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_676),
.A2(n_422),
.B1(n_9),
.B2(n_10),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_682),
.B(n_8),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_693),
.B(n_9),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_SL g750 ( 
.A(n_701),
.B(n_693),
.C(n_11),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_706),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_705),
.A2(n_676),
.B1(n_666),
.B2(n_663),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_745),
.A2(n_686),
.B1(n_692),
.B2(n_667),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_SL g754 ( 
.A1(n_712),
.A2(n_694),
.B1(n_663),
.B2(n_666),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_747),
.A2(n_686),
.B1(n_692),
.B2(n_667),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_713),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_702),
.B(n_666),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_747),
.A2(n_694),
.B1(n_686),
.B2(n_683),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_714),
.A2(n_686),
.B1(n_667),
.B2(n_694),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_728),
.B(n_667),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_748),
.B(n_40),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_SL g762 ( 
.A1(n_707),
.A2(n_690),
.B1(n_689),
.B2(n_687),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_725),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_744),
.B(n_689),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_704),
.Y(n_765)
);

OAI221xp5_ASAP7_75t_L g766 ( 
.A1(n_708),
.A2(n_690),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_711),
.Y(n_767)
);

OAI332xp33_ASAP7_75t_L g768 ( 
.A1(n_719),
.A2(n_12),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.B3(n_19),
.C1(n_21),
.C2(n_22),
.Y(n_768)
);

BUFx6f_ASAP7_75t_SL g769 ( 
.A(n_709),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_741),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_707),
.A2(n_665),
.B1(n_679),
.B2(n_671),
.Y(n_771)
);

NOR2x1_ASAP7_75t_L g772 ( 
.A(n_726),
.B(n_690),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_730),
.A2(n_687),
.B1(n_695),
.B2(n_23),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_749),
.A2(n_17),
.B1(n_19),
.B2(n_24),
.Y(n_774)
);

OAI211xp5_ASAP7_75t_L g775 ( 
.A1(n_742),
.A2(n_695),
.B(n_26),
.C(n_27),
.Y(n_775)
);

OR2x2_ASAP7_75t_SL g776 ( 
.A(n_725),
.B(n_25),
.Y(n_776)
);

OAI211xp5_ASAP7_75t_L g777 ( 
.A1(n_743),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_739),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_L g779 ( 
.A1(n_715),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.C(n_36),
.Y(n_779)
);

OAI211xp5_ASAP7_75t_SL g780 ( 
.A1(n_727),
.A2(n_33),
.B(n_38),
.C(n_39),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_718),
.A2(n_38),
.B1(n_39),
.B2(n_679),
.Y(n_781)
);

OAI33xp33_ASAP7_75t_L g782 ( 
.A1(n_731),
.A2(n_41),
.A3(n_42),
.B1(n_45),
.B2(n_46),
.B3(n_49),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_703),
.B(n_665),
.Y(n_783)
);

AOI221xp5_ASAP7_75t_L g784 ( 
.A1(n_732),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.C(n_57),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_723),
.A2(n_671),
.B1(n_64),
.B2(n_65),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_736),
.Y(n_786)
);

AOI222xp33_ASAP7_75t_L g787 ( 
.A1(n_703),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.C1(n_68),
.C2(n_69),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_760),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_751),
.B(n_737),
.Y(n_789)
);

OAI211xp5_ASAP7_75t_L g790 ( 
.A1(n_779),
.A2(n_733),
.B(n_726),
.C(n_729),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_756),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_783),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_764),
.B(n_720),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_762),
.B(n_720),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_765),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_770),
.B(n_729),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_767),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_758),
.B(n_731),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_758),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_778),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_755),
.B(n_717),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_757),
.B(n_738),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_755),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_753),
.B(n_725),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_753),
.B(n_722),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_771),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_786),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_771),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_754),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_759),
.B(n_734),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_759),
.B(n_735),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_772),
.Y(n_812)
);

AO21x2_ASAP7_75t_L g813 ( 
.A1(n_766),
.A2(n_740),
.B(n_721),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_768),
.A2(n_774),
.B1(n_773),
.B2(n_784),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_763),
.B(n_757),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_791),
.Y(n_816)
);

OAI211xp5_ASAP7_75t_SL g817 ( 
.A1(n_814),
.A2(n_750),
.B(n_787),
.C(n_777),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_809),
.A2(n_780),
.B1(n_774),
.B2(n_750),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_811),
.A2(n_782),
.B1(n_781),
.B2(n_752),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_815),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_800),
.Y(n_821)
);

AOI221xp5_ASAP7_75t_L g822 ( 
.A1(n_799),
.A2(n_775),
.B1(n_761),
.B2(n_769),
.C(n_785),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_811),
.A2(n_769),
.B1(n_716),
.B2(n_763),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_SL g824 ( 
.A1(n_809),
.A2(n_776),
.B1(n_746),
.B2(n_724),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_815),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_800),
.B(n_71),
.Y(n_826)
);

OAI31xp33_ASAP7_75t_L g827 ( 
.A1(n_790),
.A2(n_746),
.A3(n_73),
.B(n_74),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_806),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_791),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_SL g830 ( 
.A1(n_790),
.A2(n_710),
.B(n_79),
.C(n_80),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_810),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_801),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_796),
.Y(n_833)
);

NAND4xp25_ASAP7_75t_L g834 ( 
.A(n_796),
.B(n_92),
.C(n_94),
.D(n_95),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_816),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_820),
.B(n_788),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_825),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_829),
.Y(n_838)
);

OA211x2_ASAP7_75t_L g839 ( 
.A1(n_822),
.A2(n_802),
.B(n_813),
.C(n_799),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_821),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_833),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_825),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_826),
.Y(n_843)
);

NOR2x1_ASAP7_75t_L g844 ( 
.A(n_834),
.B(n_812),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_818),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_824),
.B(n_788),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_846),
.B(n_837),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_841),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_838),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_843),
.B(n_806),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_835),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_846),
.B(n_837),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_849),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_848),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_847),
.B(n_852),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_850),
.B(n_845),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_850),
.B(n_843),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_847),
.B(n_842),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_855),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_856),
.B(n_852),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_855),
.B(n_852),
.Y(n_861)
);

OAI321xp33_ASAP7_75t_L g862 ( 
.A1(n_854),
.A2(n_817),
.A3(n_819),
.B1(n_832),
.B2(n_828),
.C(n_831),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_858),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_859),
.B(n_858),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_L g865 ( 
.A1(n_862),
.A2(n_844),
.B1(n_839),
.B2(n_857),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_863),
.A2(n_819),
.B1(n_853),
.B2(n_823),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_860),
.A2(n_861),
.B(n_863),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_864),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_866),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_867),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_865),
.B(n_851),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_867),
.B(n_851),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_870),
.A2(n_815),
.B1(n_808),
.B2(n_830),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_869),
.B(n_868),
.Y(n_874)
);

NOR3x1_ASAP7_75t_L g875 ( 
.A(n_871),
.B(n_802),
.C(n_838),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_SL g876 ( 
.A1(n_872),
.A2(n_828),
.B(n_827),
.C(n_812),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_SL g877 ( 
.A(n_870),
.B(n_823),
.C(n_842),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_870),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_870),
.B(n_835),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_870),
.A2(n_800),
.B(n_812),
.Y(n_880)
);

OAI32xp33_ASAP7_75t_L g881 ( 
.A1(n_878),
.A2(n_798),
.A3(n_808),
.B1(n_803),
.B2(n_810),
.Y(n_881)
);

OAI21xp5_ASAP7_75t_L g882 ( 
.A1(n_876),
.A2(n_840),
.B(n_803),
.Y(n_882)
);

AOI211xp5_ASAP7_75t_L g883 ( 
.A1(n_874),
.A2(n_794),
.B(n_801),
.C(n_798),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_L g884 ( 
.A1(n_879),
.A2(n_815),
.B(n_794),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_875),
.B(n_836),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_880),
.B(n_836),
.Y(n_886)
);

AOI211xp5_ASAP7_75t_L g887 ( 
.A1(n_877),
.A2(n_804),
.B(n_797),
.C(n_795),
.Y(n_887)
);

OAI211xp5_ASAP7_75t_L g888 ( 
.A1(n_873),
.A2(n_804),
.B(n_795),
.C(n_797),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_SL g889 ( 
.A(n_874),
.B(n_96),
.C(n_100),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_879),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_886),
.Y(n_891)
);

OAI322xp33_ASAP7_75t_L g892 ( 
.A1(n_890),
.A2(n_807),
.A3(n_792),
.B1(n_788),
.B2(n_789),
.C1(n_805),
.C2(n_793),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_883),
.B(n_789),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_889),
.B(n_807),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_R g895 ( 
.A(n_885),
.B(n_101),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_881),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_SL g897 ( 
.A1(n_887),
.A2(n_807),
.B(n_792),
.C(n_113),
.Y(n_897)
);

AOI21xp33_ASAP7_75t_L g898 ( 
.A1(n_888),
.A2(n_882),
.B(n_884),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_889),
.Y(n_899)
);

NOR4xp75_ASAP7_75t_L g900 ( 
.A(n_891),
.B(n_793),
.C(n_805),
.D(n_114),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_891),
.Y(n_901)
);

XNOR2x1_ASAP7_75t_L g902 ( 
.A(n_899),
.B(n_103),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_894),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_896),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_893),
.Y(n_905)
);

OR5x1_ASAP7_75t_L g906 ( 
.A(n_895),
.B(n_813),
.C(n_116),
.D(n_118),
.E(n_122),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_897),
.Y(n_907)
);

NOR4xp25_ASAP7_75t_L g908 ( 
.A(n_904),
.B(n_898),
.C(n_892),
.D(n_792),
.Y(n_908)
);

NAND5xp2_ASAP7_75t_L g909 ( 
.A(n_904),
.B(n_110),
.C(n_123),
.D(n_124),
.E(n_125),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_SL g910 ( 
.A(n_901),
.B(n_126),
.C(n_128),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_SL g911 ( 
.A(n_900),
.B(n_131),
.C(n_132),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_907),
.B(n_134),
.Y(n_912)
);

AOI21xp33_ASAP7_75t_SL g913 ( 
.A1(n_902),
.A2(n_135),
.B(n_136),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_903),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_905),
.Y(n_915)
);

XNOR2x1_ASAP7_75t_L g916 ( 
.A(n_915),
.B(n_906),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_914),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_912),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_909),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_SL g920 ( 
.A1(n_908),
.A2(n_813),
.B1(n_788),
.B2(n_140),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_919),
.B(n_913),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_918),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_917),
.B(n_911),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_922),
.B(n_920),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_921),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_925),
.B(n_921),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_924),
.A2(n_916),
.B(n_923),
.Y(n_927)
);

AOI31xp67_ASAP7_75t_L g928 ( 
.A1(n_926),
.A2(n_910),
.A3(n_138),
.B(n_142),
.Y(n_928)
);

AOI222xp33_ASAP7_75t_SL g929 ( 
.A1(n_927),
.A2(n_137),
.B1(n_145),
.B2(n_146),
.C1(n_147),
.C2(n_148),
.Y(n_929)
);

AOI221x1_ASAP7_75t_L g930 ( 
.A1(n_927),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_930)
);

AOI222xp33_ASAP7_75t_SL g931 ( 
.A1(n_928),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.C1(n_158),
.C2(n_159),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_929),
.A2(n_813),
.B1(n_788),
.B2(n_162),
.Y(n_932)
);

AOI322xp5_ASAP7_75t_L g933 ( 
.A1(n_932),
.A2(n_930),
.A3(n_788),
.B1(n_164),
.B2(n_165),
.C1(n_166),
.C2(n_168),
.Y(n_933)
);

OAI221xp5_ASAP7_75t_R g934 ( 
.A1(n_933),
.A2(n_931),
.B1(n_161),
.B2(n_169),
.C(n_170),
.Y(n_934)
);

AOI211xp5_ASAP7_75t_L g935 ( 
.A1(n_934),
.A2(n_160),
.B(n_171),
.C(n_172),
.Y(n_935)
);


endmodule