module fake_jpeg_28896_n_366 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_366);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_366;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_9),
.C(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_19),
.B(n_10),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_57),
.B(n_58),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_10),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_65),
.B(n_73),
.Y(n_149)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_70),
.Y(n_128)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_21),
.B(n_8),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_28),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g118 ( 
.A(n_82),
.Y(n_118)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_86),
.Y(n_144)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_88),
.Y(n_114)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_89),
.B(n_90),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_11),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx24_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_24),
.B(n_7),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

CKINVDCx11_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_141),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_1),
.B(n_2),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_39),
.C(n_33),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_46),
.B1(n_43),
.B2(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_124),
.B1(n_148),
.B2(n_93),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_52),
.A2(n_27),
.B1(n_44),
.B2(n_41),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_134),
.B1(n_142),
.B2(n_33),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_67),
.A2(n_46),
.B1(n_43),
.B2(n_32),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_72),
.A2(n_68),
.B1(n_64),
.B2(n_60),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_140),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_95),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_79),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_56),
.A2(n_25),
.B1(n_44),
.B2(n_41),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_49),
.A2(n_22),
.B1(n_38),
.B2(n_27),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_156),
.Y(n_193)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_157),
.Y(n_208)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_158),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_166),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_106),
.A2(n_47),
.B(n_38),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_161),
.B(n_184),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_50),
.B1(n_51),
.B2(n_74),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_165),
.B1(n_124),
.B2(n_111),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_47),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_164),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_75),
.B1(n_76),
.B2(n_71),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g206 ( 
.A(n_167),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_189),
.B1(n_133),
.B2(n_109),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_91),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_188),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_17),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_173),
.Y(n_190)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

BUFx4f_ASAP7_75t_SL g173 ( 
.A(n_118),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_182),
.B1(n_108),
.B2(n_137),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_17),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_177),
.Y(n_197)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_108),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_185),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_112),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_178),
.B(n_179),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_25),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_180),
.B(n_181),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_146),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_127),
.A2(n_22),
.B(n_66),
.C(n_80),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_116),
.B(n_96),
.CI(n_13),
.CON(n_184),
.SN(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_1),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_126),
.B(n_14),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_186),
.B(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_15),
.C(n_2),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_133),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_202),
.B1(n_204),
.B2(n_178),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_176),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_137),
.B1(n_147),
.B2(n_143),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_199),
.A2(n_143),
.B1(n_147),
.B2(n_102),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_98),
.B1(n_99),
.B2(n_125),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_98),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_214),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_15),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_212),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_135),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_99),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_169),
.B(n_123),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_152),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_169),
.A2(n_128),
.B(n_109),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_219),
.C(n_218),
.Y(n_225)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_206),
.B1(n_208),
.B2(n_220),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_226),
.B1(n_243),
.B2(n_215),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_237),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_156),
.B1(n_151),
.B2(n_125),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_212),
.A2(n_183),
.B(n_160),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_227),
.A2(n_241),
.B(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_153),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_207),
.B(n_164),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_233),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_182),
.B(n_173),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_154),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_188),
.CI(n_123),
.CON(n_235),
.SN(n_235)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_190),
.B(n_172),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_197),
.B(n_107),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_240),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_211),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_167),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_200),
.A2(n_128),
.B(n_173),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_158),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_201),
.Y(n_259)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_203),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_241),
.A2(n_206),
.B1(n_192),
.B2(n_193),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_258),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_241),
.A2(n_213),
.B1(n_202),
.B2(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx3_ASAP7_75t_SL g254 ( 
.A(n_223),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_213),
.B1(n_200),
.B2(n_210),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_255),
.A2(n_267),
.B1(n_245),
.B2(n_233),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_213),
.C(n_216),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_235),
.C(n_240),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_215),
.B1(n_198),
.B2(n_220),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_261),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_198),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

OR2x2_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_118),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_236),
.B(n_238),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_271),
.Y(n_303)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_235),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_287),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_266),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_101),
.B(n_135),
.Y(n_297)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_237),
.CI(n_227),
.CON(n_275),
.SN(n_275)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_283),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_264),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_206),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_281),
.C(n_282),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_201),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_224),
.B1(n_232),
.B2(n_234),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_279),
.A2(n_286),
.B1(n_258),
.B2(n_247),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_229),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_256),
.C(n_251),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_254),
.A2(n_247),
.B(n_251),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_249),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_233),
.B1(n_236),
.B2(n_231),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_222),
.C(n_209),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_280),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_290),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_285),
.B1(n_273),
.B2(n_279),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_291),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_255),
.B1(n_267),
.B2(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_263),
.B1(n_260),
.B2(n_233),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_294),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_263),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_246),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_304),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_273),
.B(n_287),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_280),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_246),
.B(n_101),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_283),
.B(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_305),
.B(n_290),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_282),
.C(n_302),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_314),
.C(n_318),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_275),
.CI(n_269),
.CON(n_309),
.SN(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_303),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_303),
.B1(n_295),
.B2(n_296),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_281),
.C(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_316),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_275),
.C(n_270),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_300),
.B(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_320),
.A2(n_316),
.B(n_308),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_321),
.A2(n_327),
.B1(n_312),
.B2(n_311),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_322),
.A2(n_328),
.B1(n_331),
.B2(n_311),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_288),
.C(n_289),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_329),
.C(n_330),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_318),
.B(n_269),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_315),
.A2(n_299),
.B1(n_243),
.B2(n_205),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_299),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_299),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_205),
.B1(n_208),
.B2(n_155),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_307),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_209),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_334),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_319),
.B(n_313),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_335),
.A2(n_340),
.B1(n_323),
.B2(n_317),
.Y(n_343)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_338),
.Y(n_347)
);

AO221x1_ASAP7_75t_L g338 ( 
.A1(n_331),
.A2(n_312),
.B1(n_308),
.B2(n_309),
.C(n_329),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_328),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_339),
.B(n_341),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_310),
.B1(n_313),
.B2(n_309),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_330),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_342),
.B(n_343),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_336),
.A2(n_323),
.B(n_317),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_344),
.A2(n_345),
.B(n_335),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_332),
.A2(n_208),
.B1(n_157),
.B2(n_196),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_345),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_353),
.Y(n_359)
);

AOI21x1_ASAP7_75t_L g352 ( 
.A1(n_346),
.A2(n_349),
.B(n_347),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_355),
.B(n_138),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_159),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_354),
.B(n_135),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_342),
.A2(n_138),
.B(n_170),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_119),
.C(n_103),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_356),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_357),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_359),
.C(n_358),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_363),
.B(n_101),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_360),
.B(n_119),
.C(n_120),
.Y(n_363)
);

AO21x2_ASAP7_75t_L g365 ( 
.A1(n_364),
.A2(n_100),
.B(n_120),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_365),
.A2(n_102),
.B(n_100),
.Y(n_366)
);


endmodule