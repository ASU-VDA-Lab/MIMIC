module fake_jpeg_467_n_515 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_52),
.B(n_53),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_30),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_56),
.B(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_18),
.A2(n_17),
.B1(n_14),
.B2(n_2),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_58),
.A2(n_51),
.B1(n_46),
.B2(n_45),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_68),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_13),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_60),
.A2(n_62),
.B(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_13),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_13),
.C(n_2),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_29),
.C(n_47),
.Y(n_126)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_77),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_78),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_2),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_92),
.Y(n_139)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_42),
.B(n_3),
.Y(n_88)
);

HAxp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_26),
.CON(n_113),
.SN(n_113)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_3),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_27),
.B(n_12),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_27),
.B(n_12),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_27),
.Y(n_117)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_57),
.B1(n_54),
.B2(n_36),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_106),
.A2(n_107),
.B1(n_118),
.B2(n_121),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_33),
.B1(n_43),
.B2(n_19),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_29),
.B1(n_47),
.B2(n_46),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_108),
.A2(n_73),
.B1(n_94),
.B2(n_86),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_113),
.A2(n_138),
.B(n_22),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_41),
.B1(n_43),
.B2(n_19),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_83),
.B1(n_75),
.B2(n_99),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_80),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_136),
.A2(n_141),
.B1(n_70),
.B2(n_85),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_52),
.B(n_51),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_152),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_88),
.A2(n_22),
.B(n_45),
.C(n_44),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_60),
.A2(n_21),
.B1(n_44),
.B2(n_40),
.Y(n_141)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_63),
.B(n_40),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_148),
.B(n_21),
.Y(n_197)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_69),
.B(n_37),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_37),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_62),
.Y(n_165)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_62),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_160),
.B(n_172),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_43),
.B1(n_98),
.B2(n_79),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_163),
.A2(n_185),
.B1(n_205),
.B2(n_50),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_188),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_104),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_167),
.B(n_184),
.Y(n_226)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_105),
.A2(n_93),
.B1(n_97),
.B2(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_65),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_93),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_97),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_183),
.Y(n_219)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_178),
.A2(n_195),
.B(n_199),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_198),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_103),
.A2(n_20),
.B1(n_32),
.B2(n_156),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_181),
.A2(n_107),
.B1(n_118),
.B2(n_102),
.Y(n_215)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_125),
.B(n_84),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_64),
.Y(n_184)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_134),
.B(n_32),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_105),
.B(n_89),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_189),
.B(n_50),
.C(n_34),
.Y(n_251)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_134),
.B(n_20),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_193),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_115),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_115),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_197),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_123),
.B(n_87),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_116),
.B(n_21),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_201),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_91),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_146),
.Y(n_223)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_123),
.A2(n_96),
.B1(n_95),
.B2(n_26),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_149),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_211),
.Y(n_246)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_208),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_124),
.B(n_4),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_34),
.Y(n_257)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_113),
.A2(n_6),
.B(n_8),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_6),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_106),
.B(n_121),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_213),
.A2(n_220),
.B(n_229),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_215),
.B(n_228),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_132),
.B(n_149),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_112),
.B1(n_143),
.B2(n_145),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_222),
.A2(n_237),
.B1(n_243),
.B2(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_223),
.B(n_260),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_227),
.A2(n_253),
.B1(n_208),
.B2(n_182),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_187),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_160),
.A2(n_157),
.B(n_129),
.C(n_124),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_157),
.B(n_129),
.C(n_100),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_233),
.B(n_252),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_180),
.A2(n_146),
.B(n_100),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_180),
.A2(n_199),
.B1(n_183),
.B2(n_172),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_189),
.A2(n_145),
.B1(n_143),
.B2(n_112),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_198),
.B1(n_200),
.B2(n_195),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_199),
.A2(n_109),
.B1(n_50),
.B2(n_34),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_170),
.A2(n_109),
.B1(n_50),
.B2(n_34),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_257),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_170),
.A2(n_6),
.B(n_8),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_176),
.B(n_6),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_259),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_210),
.A2(n_34),
.B1(n_50),
.B2(n_10),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_187),
.B1(n_211),
.B2(n_171),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_257),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_169),
.B(n_8),
.C(n_9),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_189),
.C(n_206),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_159),
.B(n_9),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_169),
.B(n_9),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_261),
.B(n_262),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_173),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_264),
.A2(n_249),
.B(n_243),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_231),
.A2(n_210),
.B1(n_168),
.B2(n_162),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_265),
.A2(n_290),
.B1(n_242),
.B2(n_244),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_191),
.C(n_209),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_273),
.C(n_291),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_272),
.Y(n_322)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_245),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_209),
.C(n_177),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_274),
.A2(n_279),
.B1(n_284),
.B2(n_242),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_257),
.Y(n_339)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_238),
.A2(n_164),
.B1(n_174),
.B2(n_166),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_203),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_281),
.B(n_282),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_247),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_232),
.B(n_204),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_283),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_238),
.A2(n_164),
.B1(n_166),
.B2(n_174),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_179),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_295),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_179),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_287),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_214),
.B(n_207),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_289),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_190),
.C(n_186),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_246),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_296),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_214),
.B(n_161),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_299),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_219),
.B(n_195),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_239),
.Y(n_302)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_241),
.B(n_185),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_246),
.Y(n_332)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

AOI32xp33_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_231),
.A3(n_235),
.B1(n_223),
.B2(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_306),
.B(n_332),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_263),
.A2(n_220),
.B(n_248),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_313),
.A2(n_316),
.B(n_320),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_213),
.B(n_229),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_263),
.B(n_227),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_331),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_230),
.B(n_233),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_268),
.B(n_219),
.C(n_224),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_334),
.C(n_337),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_327),
.A2(n_342),
.B(n_293),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_224),
.C(n_251),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_267),
.A2(n_222),
.B1(n_258),
.B2(n_224),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_335),
.A2(n_343),
.B1(n_344),
.B2(n_266),
.Y(n_377)
);

OA22x2_ASAP7_75t_L g336 ( 
.A1(n_274),
.A2(n_250),
.B1(n_215),
.B2(n_256),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_290),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g337 ( 
.A(n_273),
.B(n_255),
.C(n_257),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_340),
.C(n_278),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_257),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_285),
.A2(n_240),
.B1(n_218),
.B2(n_252),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_341),
.A2(n_272),
.B1(n_270),
.B2(n_295),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_276),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_267),
.A2(n_218),
.B1(n_244),
.B2(n_228),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_345),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_286),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_352),
.C(n_367),
.Y(n_401)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_316),
.A2(n_285),
.B1(n_280),
.B2(n_264),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_348),
.A2(n_325),
.B1(n_319),
.B2(n_312),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_349),
.A2(n_350),
.B1(n_353),
.B2(n_359),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_341),
.A2(n_280),
.B1(n_265),
.B2(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_315),
.Y(n_351)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_261),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_333),
.B(n_300),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_360),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_342),
.A2(n_300),
.B1(n_271),
.B2(n_297),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_358),
.A2(n_340),
.B1(n_305),
.B2(n_336),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_342),
.A2(n_297),
.B1(n_282),
.B2(n_304),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_338),
.B(n_312),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_329),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_371),
.Y(n_394)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_318),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_365),
.B(n_366),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_311),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_292),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_370),
.C(n_339),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_301),
.C(n_294),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_326),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_373),
.A2(n_377),
.B1(n_336),
.B2(n_330),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_311),
.B(n_302),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_375),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_313),
.A2(n_296),
.B(n_217),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_324),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_376),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_390),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_349),
.A2(n_344),
.B1(n_320),
.B2(n_325),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_384),
.A2(n_397),
.B1(n_354),
.B2(n_368),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_386),
.A2(n_402),
.B1(n_407),
.B2(n_408),
.Y(n_412)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_389),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_374),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_324),
.Y(n_393)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_393),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_332),
.Y(n_396)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_396),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_353),
.A2(n_319),
.B1(n_336),
.B2(n_328),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_310),
.Y(n_399)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_399),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_346),
.B(n_337),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_406),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_L g402 ( 
.A1(n_356),
.A2(n_358),
.B(n_348),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_355),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_405),
.A2(n_359),
.B1(n_327),
.B2(n_307),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_369),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_375),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_408),
.A2(n_350),
.B1(n_354),
.B2(n_373),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_413),
.B1(n_418),
.B2(n_398),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_385),
.A2(n_368),
.B(n_354),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_414),
.A2(n_422),
.B(n_430),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_417),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_370),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_382),
.A2(n_355),
.B1(n_365),
.B2(n_364),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_305),
.Y(n_419)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_386),
.A2(n_307),
.B(n_367),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_309),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_425),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_266),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_379),
.B(n_277),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_429),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_217),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_380),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_389),
.B(n_277),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_385),
.A2(n_10),
.B(n_11),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_391),
.A2(n_10),
.B1(n_12),
.B2(n_394),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_431),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_384),
.B(n_393),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_432),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_399),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_396),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_417),
.B(n_401),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_443),
.Y(n_459)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_414),
.A2(n_397),
.B(n_398),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_440),
.A2(n_415),
.B(n_413),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_404),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_446),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_416),
.B(n_403),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_442),
.B(n_449),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_392),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_410),
.A2(n_380),
.B1(n_395),
.B2(n_403),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_448),
.A2(n_409),
.B1(n_432),
.B2(n_426),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_400),
.C(n_381),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_433),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_412),
.B(n_387),
.Y(n_451)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_451),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_387),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_453),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_454),
.A2(n_463),
.B1(n_411),
.B2(n_421),
.Y(n_479)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_448),
.Y(n_458)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_466),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g462 ( 
.A(n_435),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_462),
.B(n_445),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_444),
.A2(n_409),
.B1(n_411),
.B2(n_426),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_434),
.Y(n_464)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_423),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_469),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_453),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_435),
.C(n_450),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_470),
.B(n_474),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_452),
.Y(n_471)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_457),
.A2(n_438),
.B1(n_415),
.B2(n_439),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_473),
.A2(n_466),
.B1(n_465),
.B2(n_463),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_449),
.C(n_440),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_438),
.C(n_423),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_475),
.B(n_478),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_468),
.B(n_383),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_476),
.B(n_461),
.Y(n_489)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_479),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_445),
.C(n_437),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_480),
.B(n_484),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_424),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_487),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_473),
.A2(n_421),
.B1(n_434),
.B2(n_425),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_491),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_427),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_392),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_492),
.B(n_496),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_419),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_477),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_470),
.B(n_395),
.Y(n_496)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_488),
.A2(n_482),
.B(n_480),
.C(n_475),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_498),
.B(n_502),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_493),
.A2(n_477),
.B(n_483),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_500),
.B(n_494),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_485),
.B(n_483),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_503),
.B(n_490),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_505),
.B(n_506),
.Y(n_508)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_499),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_507),
.A2(n_497),
.B(n_501),
.Y(n_509)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_510),
.B(n_495),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_507),
.A2(n_501),
.B(n_495),
.Y(n_510)
);

AO21x1_ASAP7_75t_L g513 ( 
.A1(n_511),
.A2(n_512),
.B(n_486),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_491),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_513),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_429),
.Y(n_515)
);


endmodule