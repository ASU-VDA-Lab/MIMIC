module fake_jpeg_18706_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_18),
.B1(n_29),
.B2(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_50),
.B1(n_16),
.B2(n_19),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_23),
.B(n_17),
.C(n_16),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_29),
.B1(n_22),
.B2(n_30),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_22),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_32),
.C(n_28),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_29),
.B1(n_19),
.B2(n_16),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_41),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_61),
.B(n_65),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_40),
.B1(n_42),
.B2(n_41),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_64),
.B1(n_73),
.B2(n_53),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_42),
.B1(n_40),
.B2(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_27),
.B1(n_19),
.B2(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR4xp25_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_78),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_32),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_79),
.B(n_78),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_86),
.B(n_88),
.C(n_76),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_45),
.B1(n_51),
.B2(n_46),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_97),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_12),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_48),
.Y(n_102)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_107),
.Y(n_126)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_48),
.B1(n_28),
.B2(n_25),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_80),
.C(n_77),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_68),
.C(n_82),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_120),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_66),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_98),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_103),
.B(n_26),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_26),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_104),
.B1(n_90),
.B2(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_121),
.B1(n_111),
.B2(n_86),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_153),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_64),
.B1(n_85),
.B2(n_62),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_93),
.B1(n_75),
.B2(n_101),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_149),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_75),
.B1(n_93),
.B2(n_63),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_21),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_21),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_110),
.C(n_113),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_14),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_163),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_2),
.B(n_3),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_161),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_135),
.B(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_113),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_101),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_123),
.B(n_117),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_138),
.B(n_142),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_118),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_146),
.C(n_150),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_180),
.B(n_170),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_131),
.B1(n_134),
.B2(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_179),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_185),
.C(n_168),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_143),
.B1(n_140),
.B2(n_148),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_144),
.B(n_133),
.C(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_124),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_168),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_159),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_187),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_184),
.A2(n_158),
.B(n_172),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_107),
.C(n_105),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_63),
.B1(n_48),
.B2(n_5),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_190),
.C(n_192),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_185),
.B(n_177),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_178),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_174),
.A2(n_170),
.B1(n_165),
.B2(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_160),
.B(n_161),
.C(n_169),
.D(n_154),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_199),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

OAI321xp33_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_156),
.A3(n_28),
.B1(n_25),
.B2(n_13),
.C(n_9),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_3),
.B(n_4),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_208),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_196),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_25),
.Y(n_214)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_192),
.B(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_189),
.B1(n_183),
.B2(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_211),
.B(n_213),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_195),
.B1(n_188),
.B2(n_186),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_214),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_190),
.C(n_28),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_215),
.A2(n_205),
.B1(n_204),
.B2(n_202),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_209),
.A2(n_201),
.B1(n_203),
.B2(n_208),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_209),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_25),
.C2(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_217),
.C(n_200),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_219),
.C(n_218),
.Y(n_224)
);

AOI31xp67_ASAP7_75t_SL g227 ( 
.A1(n_224),
.A2(n_6),
.A3(n_8),
.B(n_9),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_227),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_10),
.C(n_6),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_229),
.C(n_8),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_231),
.Y(n_232)
);


endmodule