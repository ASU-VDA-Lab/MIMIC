module fake_jpeg_21015_n_396 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_38),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_37),
.B(n_35),
.Y(n_71)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_46),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_51),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_21),
.B(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_55),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_26),
.B(n_29),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_62),
.Y(n_101)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_22),
.B1(n_33),
.B2(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_6),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_13),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_29),
.CON(n_69),
.SN(n_69)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_71),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_78),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_76),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_35),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_88),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_36),
.A2(n_35),
.B1(n_33),
.B2(n_28),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_60),
.B1(n_55),
.B2(n_65),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_33),
.B1(n_28),
.B2(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_59),
.B1(n_22),
.B2(n_17),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_32),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_39),
.B(n_16),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_47),
.B(n_27),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_40),
.A2(n_32),
.B1(n_17),
.B2(n_18),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_32),
.B1(n_17),
.B2(n_18),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_104),
.A2(n_132),
.B1(n_140),
.B2(n_142),
.Y(n_155)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_SL g162 ( 
.A(n_109),
.B(n_134),
.C(n_135),
.Y(n_162)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_114),
.B1(n_127),
.B2(n_130),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_70),
.A2(n_48),
.B1(n_62),
.B2(n_44),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_116),
.Y(n_153)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_15),
.B1(n_18),
.B2(n_54),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_52),
.B1(n_58),
.B2(n_56),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_78),
.A2(n_58),
.B1(n_43),
.B2(n_15),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_93),
.C(n_72),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_81),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_87),
.A2(n_31),
.B1(n_50),
.B2(n_42),
.Y(n_135)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_27),
.B1(n_63),
.B2(n_10),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_93),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_85),
.A2(n_24),
.B1(n_16),
.B2(n_27),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_85),
.B(n_95),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_144),
.A2(n_169),
.B(n_174),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_97),
.B(n_71),
.C(n_83),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_173),
.B(n_157),
.C(n_174),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_98),
.B(n_100),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_147),
.A2(n_170),
.B(n_129),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_95),
.C(n_101),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_148),
.B(n_145),
.C(n_162),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_124),
.B1(n_120),
.B2(n_113),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_72),
.B1(n_103),
.B2(n_115),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_173),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_104),
.A2(n_80),
.B1(n_86),
.B2(n_84),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_171),
.B1(n_172),
.B2(n_132),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_108),
.B(n_109),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_108),
.A2(n_100),
.B(n_123),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_86),
.B1(n_84),
.B2(n_92),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_92),
.B1(n_102),
.B2(n_73),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_106),
.B(n_97),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_111),
.A2(n_92),
.B(n_94),
.C(n_79),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_106),
.B(n_125),
.C(n_89),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_172),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_179),
.Y(n_226)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_183),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_182),
.B(n_191),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_119),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_119),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_187),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_190),
.B1(n_192),
.B2(n_205),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_195),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_123),
.B1(n_77),
.B2(n_126),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_117),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_77),
.B1(n_128),
.B2(n_107),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_176),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_103),
.B1(n_110),
.B2(n_116),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g240 ( 
.A1(n_194),
.A2(n_202),
.B(n_154),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_121),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_198),
.Y(n_243)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_121),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_24),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_212),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_67),
.B(n_137),
.C(n_139),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_150),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_67),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_214),
.C(n_201),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_105),
.B1(n_11),
.B2(n_14),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_24),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

BUFx24_ASAP7_75t_L g210 ( 
.A(n_149),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_131),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_154),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_158),
.A2(n_24),
.B1(n_112),
.B2(n_6),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_24),
.B1(n_112),
.B2(n_139),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_215),
.B1(n_151),
.B2(n_152),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_24),
.B1(n_139),
.B2(n_141),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_178),
.B(n_160),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_216),
.B(n_146),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_217),
.B(n_5),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_164),
.B(n_163),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_218),
.A2(n_244),
.B(n_246),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_223),
.B(n_228),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_164),
.C(n_177),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_179),
.C(n_206),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_225),
.A2(n_229),
.B1(n_233),
.B2(n_203),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_184),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_171),
.B1(n_154),
.B2(n_176),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_230),
.B1(n_244),
.B2(n_247),
.Y(n_258)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_249),
.B(n_250),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_150),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_242),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_198),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_146),
.B(n_152),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_143),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_251),
.Y(n_279)
);

AOI32xp33_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_143),
.A3(n_9),
.B1(n_10),
.B2(n_3),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_250),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_180),
.B(n_196),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_180),
.B(n_5),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_5),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_254),
.B(n_256),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_230),
.A2(n_239),
.B1(n_190),
.B2(n_236),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_260),
.B1(n_269),
.B2(n_270),
.Y(n_282)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_262),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_239),
.A2(n_192),
.B1(n_189),
.B2(n_200),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_268),
.C(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_264),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_221),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_281),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_227),
.B(n_251),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_267),
.A2(n_238),
.B1(n_228),
.B2(n_245),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_179),
.C(n_187),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_236),
.A2(n_216),
.B1(n_213),
.B2(n_205),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_226),
.A2(n_215),
.B1(n_199),
.B2(n_182),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_223),
.A2(n_210),
.B1(n_208),
.B2(n_207),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_273),
.B1(n_225),
.B2(n_233),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_226),
.A2(n_210),
.B1(n_197),
.B2(n_181),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_0),
.C(n_1),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_276),
.C(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_0),
.C(n_1),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_0),
.C(n_1),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_222),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_280),
.B(n_234),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_227),
.B(n_1),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_218),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_3),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_285),
.A2(n_296),
.B1(n_254),
.B2(n_256),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_288),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_243),
.B1(n_226),
.B2(n_220),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_302),
.B1(n_260),
.B2(n_270),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_263),
.B(n_249),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_261),
.B(n_243),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_291),
.B(n_259),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_222),
.Y(n_292)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_219),
.Y(n_294)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_238),
.B(n_232),
.Y(n_295)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_220),
.B1(n_229),
.B2(n_233),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_258),
.B(n_265),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_297),
.A2(n_298),
.B(n_257),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_300),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_279),
.B(n_232),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_238),
.C(n_221),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_275),
.C(n_274),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_245),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_307),
.B1(n_278),
.B2(n_276),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_279),
.B(n_231),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_308),
.A2(n_311),
.B(n_302),
.Y(n_335)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_310),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_259),
.B(n_255),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_315),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_313),
.A2(n_319),
.B1(n_282),
.B2(n_285),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_272),
.C(n_264),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_320),
.C(n_324),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_298),
.A2(n_253),
.B1(n_231),
.B2(n_248),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_1),
.C(n_2),
.Y(n_320)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_2),
.C(n_3),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_327),
.C(n_328),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_303),
.C(n_290),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_2),
.C(n_3),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_2),
.C(n_4),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_289),
.B1(n_282),
.B2(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_323),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_333),
.A2(n_338),
.B1(n_344),
.B2(n_310),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_346),
.Y(n_355)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_336),
.Y(n_352)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_340),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_311),
.B(n_326),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_342),
.B(n_343),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_319),
.A2(n_289),
.B(n_304),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_313),
.A2(n_287),
.B1(n_305),
.B2(n_286),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_325),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_322),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_316),
.C(n_327),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_350),
.C(n_358),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_353),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_315),
.C(n_312),
.Y(n_350)
);

AOI22x1_ASAP7_75t_SL g354 ( 
.A1(n_335),
.A2(n_288),
.B1(n_300),
.B2(n_309),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_354),
.A2(n_344),
.B1(n_345),
.B2(n_332),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_307),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_305),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_349),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_334),
.C(n_341),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_342),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_359),
.B(n_343),
.Y(n_365)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_365),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_362),
.B(n_369),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_341),
.C(n_339),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_366),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_352),
.B(n_332),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_370),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_338),
.C(n_320),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_355),
.B(n_328),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_371),
.A2(n_353),
.B(n_324),
.Y(n_376)
);

OAI322xp33_ASAP7_75t_L g372 ( 
.A1(n_361),
.A2(n_347),
.A3(n_351),
.B1(n_350),
.B2(n_356),
.C1(n_333),
.C2(n_360),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_301),
.Y(n_385)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_363),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_375),
.B(n_376),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_SL g378 ( 
.A(n_363),
.B(n_333),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_367),
.B(n_370),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_364),
.A2(n_301),
.B(n_11),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_4),
.B(n_11),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_381),
.A2(n_385),
.B(n_386),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_382),
.B(n_383),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_379),
.B(n_362),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_377),
.A2(n_4),
.B(n_12),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_12),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_387),
.A2(n_374),
.B(n_373),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_390),
.B(n_391),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_372),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_13),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_389),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_394),
.A2(n_392),
.B1(n_13),
.B2(n_14),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_395),
.B(n_14),
.Y(n_396)
);


endmodule