module fake_ariane_2517_n_381 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_117, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_112, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_108, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_381);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_117;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_112;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_108;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_381;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_347;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_245;
wire n_319;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_139;
wire n_130;
wire n_349;
wire n_346;
wire n_214;
wire n_348;
wire n_379;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_327;
wire n_372;
wire n_377;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_272;
wire n_339;
wire n_167;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_143;
wire n_152;
wire n_120;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_331;
wire n_267;
wire n_335;
wire n_350;
wire n_291;
wire n_344;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_301;
wire n_248;
wire n_277;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_303;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_333;
wire n_376;
wire n_221;
wire n_321;
wire n_361;
wire n_149;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_343;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_249;
wire n_212;
wire n_123;
wire n_355;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_216;
wire n_223;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_203;
wire n_378;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_159;
wire n_358;
wire n_131;
wire n_263;
wire n_360;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_118;
wire n_121;
wire n_353;
wire n_241;
wire n_357;
wire n_191;
wire n_211;
wire n_322;
wire n_251;
wire n_351;
wire n_359;
wire n_155;
wire n_127;

INVx1_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_66),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_7),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_5),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_1),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_24),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_92),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_44),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_77),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_11),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_29),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_32),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_83),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_18),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

BUFx8_ASAP7_75t_SL g149 ( 
.A(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_5),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_9),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_10),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_7),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_30),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_4),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_1),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

INVxp33_ASAP7_75t_SL g162 ( 
.A(n_79),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_67),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_112),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_47),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_21),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_49),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_2),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_73),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_80),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_31),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_118),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_0),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_3),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_129),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_192)
);

AND2x4_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_6),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_137),
.B(n_8),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_181),
.B(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_176),
.B1(n_175),
.B2(n_119),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_127),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_179),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_127),
.Y(n_207)
);

OR2x6_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_185),
.B(n_128),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_120),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_141),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_121),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_195),
.B(n_138),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_174),
.B1(n_161),
.B2(n_155),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_192),
.B1(n_188),
.B2(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_122),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_126),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_148),
.B(n_125),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_124),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_210),
.B(n_192),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_202),
.B1(n_210),
.B2(n_221),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_130),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_152),
.B1(n_171),
.B2(n_170),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_207),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_132),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_133),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_151),
.B1(n_169),
.B2(n_136),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_223),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_145),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_134),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_203),
.B(n_139),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_201),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

OR2x6_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_143),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_222),
.B(n_219),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_140),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_146),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_142),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_226),
.A2(n_166),
.B1(n_153),
.B2(n_147),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

NOR2x1p5_ASAP7_75t_SL g265 ( 
.A(n_231),
.B(n_144),
.Y(n_265)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_167),
.B(n_154),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_168),
.C(n_164),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_228),
.A2(n_163),
.B(n_159),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_234),
.A2(n_157),
.B1(n_225),
.B2(n_173),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_225),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_220),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_232),
.A2(n_220),
.B(n_13),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_220),
.B(n_14),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_12),
.B(n_15),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_230),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_241),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_281)
);

HB1xp67_ASAP7_75t_SL g282 ( 
.A(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_249),
.A2(n_20),
.B(n_22),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_117),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_241),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

BUFx8_ASAP7_75t_L g288 ( 
.A(n_283),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_242),
.B(n_239),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_269),
.B(n_263),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_259),
.A2(n_257),
.B(n_251),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_262),
.A2(n_239),
.B(n_246),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_245),
.B(n_227),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_245),
.B(n_25),
.C(n_26),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_245),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_267),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_258),
.B(n_27),
.C(n_28),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

AO32x2_ASAP7_75t_L g300 ( 
.A1(n_271),
.A2(n_258),
.A3(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_270),
.Y(n_301)
);

AO31x2_ASAP7_75t_L g302 ( 
.A1(n_264),
.A2(n_258),
.A3(n_36),
.B(n_37),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_261),
.A2(n_23),
.B(n_38),
.Y(n_303)
);

O2A1O1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_261),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_42),
.B(n_43),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_281),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

AO21x2_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_285),
.B(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_273),
.B(n_268),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_292),
.A2(n_264),
.B(n_279),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_303),
.B(n_298),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_277),
.B(n_280),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_293),
.A2(n_287),
.B(n_265),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_266),
.B(n_281),
.C(n_267),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

BUFx8_ASAP7_75t_SL g320 ( 
.A(n_297),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_54),
.B(n_55),
.Y(n_321)
);

AO21x2_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_296),
.B(n_302),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_299),
.Y(n_323)
);

AO21x2_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_302),
.B(n_300),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_309),
.A2(n_290),
.B1(n_307),
.B2(n_288),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_300),
.B(n_58),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_56),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_59),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_326),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_330),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_300),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_328),
.B(n_313),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_324),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_332),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_324),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_311),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_311),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_314),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_338),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_61),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_64),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_320),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_65),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_353),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_340),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_346),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_343),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_345),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_355),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_358),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_359),
.B(n_351),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_359),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_364),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_362),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_365),
.B(n_352),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_366),
.A2(n_363),
.B(n_343),
.Y(n_368)
);

O2A1O1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_368),
.A2(n_366),
.B(n_354),
.C(n_361),
.Y(n_369)
);

O2A1O1Ixp5_ASAP7_75t_L g370 ( 
.A1(n_367),
.A2(n_347),
.B(n_360),
.C(n_357),
.Y(n_370)
);

NOR4xp25_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_349),
.C(n_350),
.D(n_342),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_370),
.B(n_350),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_68),
.Y(n_373)
);

NAND4xp75_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_371),
.C(n_349),
.D(n_321),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_374),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_375),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_72),
.B(n_74),
.Y(n_377)
);

AOI222xp33_ASAP7_75t_SL g378 ( 
.A1(n_376),
.A2(n_75),
.B1(n_78),
.B2(n_81),
.C1(n_82),
.C2(n_87),
.Y(n_378)
);

OAI222xp33_ASAP7_75t_L g379 ( 
.A1(n_377),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.C1(n_101),
.C2(n_104),
.Y(n_379)
);

OAI22x1_ASAP7_75t_L g380 ( 
.A1(n_379),
.A2(n_378),
.B1(n_110),
.B2(n_113),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_109),
.B(n_115),
.Y(n_381)
);


endmodule