module fake_jpeg_23778_n_193 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_193);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_25),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_37),
.CON(n_50),
.SN(n_50)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_26),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_44),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_16),
.B1(n_25),
.B2(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_47),
.B1(n_48),
.B2(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_22),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_16),
.B1(n_25),
.B2(n_21),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_62),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_69),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_22),
.B1(n_27),
.B2(n_17),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_64),
.B1(n_71),
.B2(n_43),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_53),
.B1(n_42),
.B2(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_17),
.B1(n_15),
.B2(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_70),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_26),
.B1(n_17),
.B2(n_15),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_38),
.C(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_88),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_53),
.B(n_39),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_56),
.B(n_55),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_39),
.B1(n_41),
.B2(n_47),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_82),
.B1(n_87),
.B2(n_72),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_42),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_83),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_41),
.B1(n_47),
.B2(n_62),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_84),
.B1(n_89),
.B2(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_86),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_75),
.B1(n_80),
.B2(n_74),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_55),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_39),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_40),
.B1(n_46),
.B2(n_52),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_100),
.B(n_104),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_75),
.B1(n_74),
.B2(n_79),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_88),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_107),
.Y(n_112)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_101),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_0),
.B(n_17),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_70),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_37),
.B(n_54),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_0),
.B(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_111),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_123),
.B(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_92),
.B(n_35),
.CI(n_61),
.CON(n_115),
.SN(n_115)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_107),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_93),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_54),
.C(n_68),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_120),
.C(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_2),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_2),
.B(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_94),
.B1(n_106),
.B2(n_103),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_131),
.A2(n_138),
.B1(n_108),
.B2(n_115),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_136),
.B(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_101),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_91),
.C(n_95),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_137),
.B(n_110),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_93),
.B1(n_98),
.B2(n_95),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_119),
.C(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_151),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_132),
.B(n_111),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_146),
.C(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_124),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_126),
.B1(n_117),
.B2(n_5),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_95),
.C(n_110),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_3),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_112),
.C(n_109),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_112),
.C(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_134),
.C(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_152),
.A2(n_133),
.B1(n_130),
.B2(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_155),
.B(n_158),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_130),
.B1(n_116),
.B2(n_128),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_161),
.B1(n_6),
.B2(n_8),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_126),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_150),
.C(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

AOI31xp67_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_117),
.A3(n_5),
.B(n_6),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_141),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_167),
.C(n_172),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_161),
.A2(n_149),
.B1(n_146),
.B2(n_7),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_4),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_4),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_171),
.B(n_10),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_8),
.C(n_9),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_163),
.B1(n_159),
.B2(n_153),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_178),
.B1(n_172),
.B2(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_160),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_10),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_181),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_177),
.B(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_182),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_11),
.C(n_12),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_174),
.B(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_188),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_175),
.C(n_12),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_11),
.B(n_13),
.C(n_186),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_189),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_13),
.Y(n_193)
);


endmodule