module fake_jpeg_10552_n_272 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_59),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_22),
.B1(n_44),
.B2(n_27),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_70),
.B1(n_15),
.B2(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_27),
.B1(n_15),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_69),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_27),
.B1(n_15),
.B2(n_37),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_78),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_85),
.B1(n_89),
.B2(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_53),
.B1(n_41),
.B2(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_80),
.Y(n_106)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_35),
.B1(n_37),
.B2(n_52),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_38),
.B1(n_25),
.B2(n_16),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_37),
.B1(n_35),
.B2(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_90),
.B1(n_41),
.B2(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_31),
.B(n_28),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_72),
.B(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_28),
.B1(n_53),
.B2(n_41),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_50),
.B1(n_48),
.B2(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_47),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_103),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_68),
.B(n_65),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_102),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_114),
.B1(n_88),
.B2(n_84),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_31),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_110),
.B1(n_79),
.B2(n_81),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_72),
.B(n_63),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_111),
.B(n_115),
.C(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_74),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_36),
.B1(n_54),
.B2(n_49),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_43),
.B(n_25),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_94),
.B1(n_85),
.B2(n_38),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_81),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_16),
.B(n_25),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_120),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_76),
.B1(n_92),
.B2(n_91),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_137),
.B1(n_95),
.B2(n_67),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_76),
.C(n_82),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_34),
.C(n_29),
.Y(n_148)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_110),
.B1(n_98),
.B2(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_96),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_17),
.B1(n_24),
.B2(n_78),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_136),
.B(n_14),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_94),
.B1(n_24),
.B2(n_17),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_23),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_102),
.B(n_32),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_67),
.B1(n_32),
.B2(n_29),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_115),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_97),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_142),
.B(n_125),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_151),
.B1(n_154),
.B2(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_134),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_149),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_101),
.C(n_95),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_95),
.B1(n_32),
.B2(n_29),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_32),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_29),
.C(n_23),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_26),
.B1(n_18),
.B2(n_13),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_14),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_14),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_160),
.C(n_128),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_14),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_121),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_167),
.C(n_175),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_121),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_178),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_154),
.B1(n_144),
.B2(n_142),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_14),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_174),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_122),
.B1(n_120),
.B2(n_123),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_172),
.A2(n_157),
.B1(n_155),
.B2(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_132),
.C(n_129),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_132),
.C(n_23),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_21),
.C(n_14),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_173),
.B1(n_172),
.B2(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_199),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_26),
.B1(n_18),
.B2(n_13),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_26),
.B1(n_18),
.B2(n_2),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_193),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_26),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_200),
.B(n_21),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_21),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_166),
.C(n_171),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_190),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_164),
.C(n_167),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.C(n_205),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_164),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_166),
.C(n_177),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_0),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_1),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_216),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_21),
.C(n_3),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_218),
.C(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_214),
.B(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_5),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_197),
.B(n_192),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_6),
.B(n_8),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_5),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_226),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_185),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_218),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_192),
.B1(n_197),
.B2(n_193),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_190),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_200),
.C(n_189),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_210),
.C(n_215),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_214),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_6),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_206),
.C(n_211),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_244),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_237),
.Y(n_245)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_240),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_10),
.B1(n_11),
.B2(n_236),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_8),
.C(n_9),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_9),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_221),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_221),
.B1(n_229),
.B2(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_237),
.B1(n_244),
.B2(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_249),
.B(n_252),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_233),
.B(n_11),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_219),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_10),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_250),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_246),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_259),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_251),
.C(n_245),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_11),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_261),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_258),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_259),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_265),
.B(n_263),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_266),
.B(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_247),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_271),
.Y(n_272)
);


endmodule