module real_jpeg_4202_n_11 (n_5, n_4, n_8, n_0, n_1, n_51, n_53, n_2, n_6, n_7, n_52, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_51;
input n_53;
input n_2;
input n_6;
input n_7;
input n_52;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_49;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_48;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_3),
.A2(n_17),
.B(n_51),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_36),
.C(n_53),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_5),
.C(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_6),
.A2(n_7),
.B(n_25),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_7),
.C(n_20),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_10),
.C(n_14),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_10),
.B(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_22),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_18),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_15),
.A2(n_44),
.B(n_45),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_39),
.B(n_40),
.Y(n_38)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_43),
.B(n_46),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_42),
.Y(n_23)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_39),
.C(n_40),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_38),
.B(n_41),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B(n_35),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_52),
.Y(n_34)
);


endmodule