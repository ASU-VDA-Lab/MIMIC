module fake_jpeg_29977_n_481 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_481);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_481;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_50),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_16),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_62),
.Y(n_110)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_20),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_89),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_0),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_64),
.B(n_65),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx11_ASAP7_75t_SL g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_96),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_20),
.B(n_1),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_83),
.C(n_36),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_38),
.A2(n_2),
.B(n_3),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx2_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_86),
.B(n_37),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_23),
.B(n_2),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_23),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_24),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_27),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_117),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_36),
.B1(n_45),
.B2(n_48),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_111),
.A2(n_48),
.B1(n_29),
.B2(n_33),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_50),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_112),
.B(n_52),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_36),
.B1(n_26),
.B2(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_114),
.B1(n_120),
.B2(n_128),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_34),
.B1(n_47),
.B2(n_44),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_139),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_51),
.A2(n_56),
.B1(n_77),
.B2(n_60),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_47),
.B1(n_34),
.B2(n_29),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_57),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_129),
.A2(n_72),
.B1(n_79),
.B2(n_34),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_138),
.B(n_45),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_46),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_81),
.B(n_46),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_39),
.Y(n_156)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_156),
.B(n_162),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_70),
.B1(n_80),
.B2(n_94),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_158),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_37),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_159),
.B(n_171),
.C(n_193),
.Y(n_245)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_160),
.Y(n_219)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_165),
.Y(n_220)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_168),
.Y(n_255)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_100),
.B(n_75),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_172),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_102),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_178),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_110),
.A2(n_19),
.B(n_68),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_175),
.A2(n_30),
.B(n_28),
.Y(n_248)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_125),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_104),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_199),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_SL g180 ( 
.A1(n_111),
.A2(n_94),
.B(n_27),
.C(n_85),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_180),
.A2(n_113),
.B(n_128),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_110),
.B(n_32),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_189),
.Y(n_210)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_129),
.A2(n_78),
.B1(n_92),
.B2(n_71),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_202),
.B1(n_120),
.B2(n_114),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_195),
.Y(n_228)
);

INVx6_ASAP7_75t_SL g185 ( 
.A(n_151),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_61),
.B1(n_53),
.B2(n_55),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_186),
.A2(n_204),
.B1(n_206),
.B2(n_101),
.Y(n_238)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_150),
.B1(n_141),
.B2(n_147),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_99),
.B(n_98),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_103),
.B(n_39),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_200),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_109),
.B(n_97),
.C(n_88),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_121),
.Y(n_195)
);

NAND2x1p5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_27),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_208),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_134),
.B(n_32),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_203),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_141),
.A2(n_28),
.B1(n_45),
.B2(n_33),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

BUFx2_ASAP7_75t_SL g207 ( 
.A(n_101),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_145),
.B(n_87),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g244 ( 
.A(n_209),
.B(n_148),
.Y(n_244)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_158),
.A3(n_180),
.B1(n_155),
.B2(n_159),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_240),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_226),
.A2(n_231),
.B1(n_239),
.B2(n_165),
.Y(n_290)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_166),
.A2(n_29),
.B(n_33),
.Y(n_230)
);

OAI221xp5_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_202),
.B1(n_209),
.B2(n_183),
.C(n_203),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_171),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_234),
.B(n_195),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_235),
.A2(n_234),
.B1(n_242),
.B2(n_226),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_106),
.B(n_132),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_237),
.A2(n_243),
.B(n_4),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_171),
.A2(n_150),
.B1(n_147),
.B2(n_143),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_184),
.A2(n_30),
.A3(n_143),
.B1(n_27),
.B2(n_148),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_137),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_250),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_106),
.B(n_3),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_244),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_253),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_166),
.B(n_137),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_157),
.B(n_2),
.C(n_3),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_4),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_231),
.A2(n_196),
.B(n_186),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_257),
.A2(n_287),
.B(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_215),
.B(n_176),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_274),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_264),
.B(n_265),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_215),
.B(n_170),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_266),
.A2(n_271),
.B1(n_239),
.B2(n_244),
.Y(n_305)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_214),
.B(n_194),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_268),
.B(n_275),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_210),
.B(n_160),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_269),
.B(n_292),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_199),
.C(n_169),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_270),
.B(n_276),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_212),
.A2(n_182),
.B1(n_177),
.B2(n_197),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_272),
.Y(n_308)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_206),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_161),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_279),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_228),
.B(n_167),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_280),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_218),
.B(n_217),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_228),
.B(n_163),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_228),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_282),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_294),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_295),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_252),
.A2(n_5),
.B(n_6),
.Y(n_288)
);

AO21x2_ASAP7_75t_L g289 ( 
.A1(n_240),
.A2(n_191),
.B(n_204),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_289),
.A2(n_216),
.B1(n_241),
.B2(n_219),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_290),
.A2(n_291),
.B1(n_249),
.B2(n_216),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_244),
.A2(n_164),
.B1(n_191),
.B2(n_7),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_210),
.B(n_5),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_6),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_6),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_252),
.B(n_7),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_221),
.B(n_7),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_282),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_310),
.B1(n_311),
.B2(n_315),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_237),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_313),
.C(n_285),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_262),
.A2(n_249),
.B1(n_233),
.B2(n_213),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_301),
.A2(n_259),
.B(n_280),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_305),
.A2(n_316),
.B1(n_291),
.B2(n_283),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_290),
.A2(n_253),
.B1(n_248),
.B2(n_243),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_256),
.A2(n_253),
.B1(n_213),
.B2(n_223),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_225),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_258),
.A2(n_253),
.B1(n_232),
.B2(n_221),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_271),
.A2(n_223),
.B1(n_246),
.B2(n_241),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_258),
.A2(n_289),
.B1(n_262),
.B2(n_278),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_317),
.A2(n_319),
.B1(n_323),
.B2(n_327),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_251),
.B1(n_246),
.B2(n_220),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_328),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_289),
.A2(n_211),
.B1(n_220),
.B2(n_219),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_289),
.A2(n_211),
.B1(n_229),
.B2(n_222),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_286),
.A2(n_229),
.B1(n_222),
.B2(n_233),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_332),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_260),
.B(n_236),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_331),
.B(n_276),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_222),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_257),
.A2(n_236),
.B(n_9),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_288),
.B(n_286),
.Y(n_339)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_284),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_343),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_339),
.A2(n_344),
.B(n_359),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_318),
.A2(n_259),
.B(n_287),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_340),
.B(n_350),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_329),
.Y(n_365)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_314),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_333),
.A2(n_289),
.B(n_264),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_345),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_294),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_351),
.C(n_360),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_353),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_324),
.B(n_296),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_295),
.C(n_266),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_309),
.B(n_322),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_352),
.B(n_354),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_312),
.B(n_295),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_263),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_321),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_356),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_303),
.B(n_267),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_357),
.A2(n_319),
.B1(n_328),
.B2(n_327),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_273),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_364),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_275),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_298),
.C(n_329),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_298),
.B(n_272),
.C(n_9),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_350),
.C(n_352),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_306),
.A2(n_8),
.B(n_10),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_363),
.A2(n_307),
.B(n_320),
.Y(n_384)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_365),
.B(n_351),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_331),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_376),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_348),
.A2(n_305),
.B1(n_316),
.B2(n_310),
.Y(n_372)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_372),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_302),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_378),
.B(n_387),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_302),
.C(n_322),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_380),
.C(n_382),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_326),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_306),
.C(n_311),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_348),
.A2(n_307),
.B1(n_297),
.B2(n_304),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_362),
.B1(n_346),
.B2(n_334),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_338),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_386),
.A2(n_357),
.B1(n_339),
.B2(n_337),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_344),
.A2(n_320),
.B(n_308),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_359),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_390)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_390),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_359),
.A2(n_11),
.B1(n_14),
.B2(n_362),
.Y(n_391)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_391),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_397),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_371),
.C(n_367),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_402),
.C(n_367),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_395),
.A2(n_409),
.B1(n_372),
.B2(n_373),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_410),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_355),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_361),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_400),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_346),
.C(n_340),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_378),
.B(n_343),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_406),
.Y(n_424)
);

NOR3xp33_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_356),
.C(n_334),
.Y(n_404)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_343),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_335),
.Y(n_407)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_365),
.B(n_379),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_413),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_345),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_415),
.A2(n_426),
.B1(n_428),
.B2(n_430),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_392),
.A2(n_377),
.B(n_387),
.Y(n_416)
);

AOI21x1_ASAP7_75t_L g441 ( 
.A1(n_416),
.A2(n_408),
.B(n_405),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_376),
.C(n_382),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_417),
.B(n_418),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_380),
.C(n_366),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_431),
.C(n_396),
.Y(n_439)
);

INVx13_ASAP7_75t_L g420 ( 
.A(n_412),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_398),
.A2(n_386),
.B1(n_366),
.B2(n_390),
.Y(n_426)
);

INVx13_ASAP7_75t_L g427 ( 
.A(n_407),
.Y(n_427)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_427),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_398),
.A2(n_384),
.B1(n_388),
.B2(n_375),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_408),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_413),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_394),
.C(n_393),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_434),
.Y(n_456)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_433),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_421),
.B(n_401),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_421),
.B(n_393),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_436),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_410),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_438),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_409),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_440),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_405),
.Y(n_440)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_441),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_424),
.A2(n_375),
.B(n_363),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_443),
.A2(n_416),
.B(n_428),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_415),
.A2(n_364),
.B1(n_342),
.B2(n_14),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_444),
.B(n_414),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_455),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_441),
.A2(n_424),
.B(n_431),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_449),
.A2(n_450),
.B(n_438),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_445),
.A2(n_422),
.B(n_429),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_451),
.B(n_427),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_423),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_425),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_426),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_452),
.B(n_446),
.C(n_435),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_448),
.C(n_423),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_461),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_453),
.B(n_435),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_462),
.A2(n_450),
.B(n_451),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_463),
.B(n_465),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_456),
.A2(n_430),
.B1(n_422),
.B2(n_429),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_464),
.A2(n_466),
.B1(n_442),
.B2(n_14),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_439),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_454),
.A2(n_442),
.B1(n_420),
.B2(n_437),
.Y(n_466)
);

OA21x2_ASAP7_75t_SL g467 ( 
.A1(n_459),
.A2(n_455),
.B(n_446),
.Y(n_467)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_467),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_468),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_469),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_471),
.B(n_469),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_476),
.A2(n_477),
.B(n_475),
.Y(n_478)
);

OAI31xp33_ASAP7_75t_SL g477 ( 
.A1(n_474),
.A2(n_464),
.A3(n_472),
.B(n_470),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_462),
.C(n_458),
.Y(n_479)
);

XNOR2x1_ASAP7_75t_SL g480 ( 
.A(n_479),
.B(n_466),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_480),
.B(n_14),
.Y(n_481)
);


endmodule