module real_jpeg_6538_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_0),
.Y(n_531)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_1),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_1),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_1),
.Y(n_281)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_1),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_1),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_2),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_2),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_2),
.A2(n_51),
.B1(n_202),
.B2(n_272),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_2),
.A2(n_202),
.B1(n_283),
.B2(n_388),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_2),
.A2(n_202),
.B1(n_449),
.B2(n_451),
.Y(n_448)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_3),
.Y(n_188)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_3),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_3),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_4),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_46),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_4),
.A2(n_46),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_4),
.A2(n_46),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_5),
.A2(n_39),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_5),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_5),
.A2(n_187),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_5),
.A2(n_187),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_5),
.A2(n_187),
.B1(n_422),
.B2(n_425),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_7),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_8),
.Y(n_116)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_8),
.Y(n_382)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_10),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_11),
.A2(n_215),
.B1(n_217),
.B2(n_220),
.Y(n_214)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_11),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_11),
.A2(n_220),
.B1(n_258),
.B2(n_269),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_11),
.A2(n_179),
.B1(n_220),
.B2(n_303),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g362 ( 
.A1(n_11),
.A2(n_220),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_13),
.A2(n_160),
.B1(n_217),
.B2(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_13),
.B(n_382),
.C(n_383),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_13),
.B(n_88),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_13),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_13),
.B(n_130),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_13),
.B(n_210),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_14),
.A2(n_55),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_14),
.A2(n_73),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_14),
.A2(n_73),
.B1(n_216),
.B2(n_224),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_14),
.A2(n_73),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_16),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_16),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_16),
.A2(n_70),
.B1(n_167),
.B2(n_172),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_16),
.A2(n_70),
.B1(n_223),
.B2(n_228),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_16),
.A2(n_70),
.B1(n_207),
.B2(n_320),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_17),
.A2(n_50),
.B1(n_54),
.B2(n_57),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_17),
.A2(n_57),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_17),
.A2(n_57),
.B1(n_167),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_17),
.A2(n_57),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_18),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_18),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_18),
.A2(n_191),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_18),
.A2(n_191),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_18),
.A2(n_191),
.B1(n_304),
.B2(n_395),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_526),
.B(n_528),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_59),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_47),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B(n_41),
.Y(n_23)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_24),
.B(n_190),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_24),
.B(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_25),
.A2(n_48),
.B1(n_186),
.B2(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_25),
.B(n_160),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_30),
.Y(n_150)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_30),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_32),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_32),
.Y(n_204)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_32),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_32),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_34),
.B(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_34),
.A2(n_248),
.B(n_252),
.Y(n_247)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_38),
.Y(n_154)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_39),
.Y(n_192)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_40),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_40),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_47)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_47),
.B(n_62),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_58),
.B1(n_66),
.B2(n_71),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_48),
.A2(n_49),
.B1(n_58),
.B2(n_71),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_48),
.A2(n_253),
.B(n_271),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_48),
.A2(n_58),
.B1(n_66),
.B2(n_498),
.Y(n_497)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_53),
.Y(n_251)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_58),
.A2(n_186),
.B(n_189),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_139),
.B(n_525),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_135),
.C(n_136),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_63),
.A2(n_64),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.C(n_106),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_65),
.B(n_513),
.Y(n_512)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_74),
.A2(n_106),
.B1(n_107),
.B2(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_74),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_75),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_75),
.A2(n_102),
.B1(n_199),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_75),
.A2(n_102),
.B1(n_268),
.B2(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_75),
.A2(n_97),
.B1(n_102),
.B2(n_502),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_88),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_80),
.Y(n_462)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_82),
.Y(n_210)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_83),
.Y(n_350)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_86),
.Y(n_346)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_87),
.Y(n_201)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_87),
.Y(n_257)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_88),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

AOI22x1_ASAP7_75t_L g265 ( 
.A1(n_88),
.A2(n_137),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_88),
.A2(n_137),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_92),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_92),
.Y(n_244)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_92),
.Y(n_402)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_92),
.Y(n_465)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_111),
.B1(n_114),
.B2(n_117),
.Y(n_110)
);

INVx11_ASAP7_75t_L g400 ( 
.A(n_93),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_94),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_94),
.Y(n_231)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_95),
.Y(n_466)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_98),
.Y(n_258)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_102),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_102),
.A2(n_255),
.B(n_300),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_106),
.A2(n_107),
.B1(n_500),
.B2(n_501),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_106),
.B(n_497),
.C(n_500),
.Y(n_508)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_129),
.B(n_131),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_108),
.A2(n_129),
.B1(n_214),
.B2(n_221),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_108),
.A2(n_375),
.B(n_377),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_108),
.A2(n_129),
.B1(n_399),
.B2(n_448),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_108),
.A2(n_377),
.B(n_448),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_109),
.B(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_109),
.A2(n_130),
.B1(n_222),
.B2(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_109),
.A2(n_130),
.B1(n_277),
.B2(n_327),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_109),
.A2(n_130),
.B1(n_327),
.B2(n_353),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_120),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_120),
.A2(n_241),
.B(n_399),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_128),
.Y(n_120)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_124),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_125),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_127),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g426 ( 
.A(n_127),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_129),
.A2(n_214),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_130),
.B(n_242),
.Y(n_377)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_131),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_133),
.Y(n_330)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_133),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_135),
.B(n_136),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_198),
.B(n_205),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_137),
.B(n_266),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_137),
.A2(n_205),
.B(n_454),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_519),
.B(n_524),
.Y(n_139)
);

AOI21x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_491),
.B(n_516),
.Y(n_140)
);

OAI311xp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_312),
.A3(n_368),
.B1(n_485),
.C1(n_490),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_290),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_144),
.A2(n_487),
.B(n_488),
.Y(n_486)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_259),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_145),
.B(n_259),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_211),
.C(n_239),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_146),
.B(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_183),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_147),
.B(n_184),
.C(n_197),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_161),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_148),
.A2(n_161),
.B1(n_162),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_148),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_151),
.A3(n_152),
.B1(n_155),
.B2(n_159),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_SL g248 ( 
.A1(n_159),
.A2(n_160),
.B(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_160),
.A2(n_163),
.B(n_391),
.Y(n_418)
);

OAI21xp33_ASAP7_75t_SL g454 ( 
.A1(n_160),
.A2(n_320),
.B(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_170),
.B1(n_173),
.B2(n_176),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_163),
.A2(n_234),
.B1(n_279),
.B2(n_282),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_163),
.A2(n_282),
.B(n_332),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_163),
.A2(n_387),
.B(n_391),
.Y(n_386)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_164),
.A2(n_177),
.B1(n_233),
.B2(n_237),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_164),
.A2(n_171),
.B1(n_302),
.B2(n_307),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_164),
.B(n_394),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_164),
.A2(n_435),
.B1(n_436),
.B2(n_437),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_166),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_166),
.Y(n_417)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_166),
.Y(n_429)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_169),
.Y(n_287)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_169),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_169),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_182),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_196),
.B2(n_197),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_189),
.B(n_361),
.Y(n_360)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_211),
.A2(n_212),
.B1(n_239),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_232),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_213),
.B(n_232),
.Y(n_263)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_227),
.Y(n_380)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_231),
.Y(n_376)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_235),
.Y(n_395)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_236),
.Y(n_384)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.C(n_254),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_240),
.B(n_254),
.Y(n_293)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI32xp33_ASAP7_75t_L g460 ( 
.A1(n_244),
.A2(n_258),
.A3(n_456),
.B1(n_461),
.B2(n_463),
.Y(n_460)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_246),
.A2(n_247),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_260),
.B(n_275),
.C(n_288),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_275),
.B1(n_288),
.B2(n_289),
.Y(n_261)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_263),
.B(n_265),
.C(n_274),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_265),
.Y(n_273)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_278),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_309),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_291),
.B(n_309),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.C(n_298),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_292),
.B(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_295),
.A2(n_296),
.B1(n_298),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_298),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_308),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_299),
.B(n_476),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_301),
.B(n_308),
.Y(n_476)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_302),
.Y(n_459)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_365),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_SL g485 ( 
.A1(n_313),
.A2(n_365),
.B(n_486),
.C(n_489),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_337),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_314),
.B(n_337),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_324),
.C(n_336),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g367 ( 
.A(n_315),
.B(n_324),
.CI(n_336),
.CON(n_367),
.SN(n_367)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_318),
.C(n_323),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_331),
.B2(n_335),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_331),
.Y(n_357)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_331),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_331),
.A2(n_335),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_331),
.A2(n_357),
.B(n_360),
.Y(n_494)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_338),
.B(n_341),
.C(n_355),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_355),
.B2(n_356),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_351),
.B(n_354),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_343),
.B(n_352),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_345),
.Y(n_502)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g493 ( 
.A(n_354),
.B(n_494),
.CI(n_495),
.CON(n_493),
.SN(n_493)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_354),
.B(n_494),
.C(n_495),
.Y(n_515)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_362),
.Y(n_498)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_363),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_366),
.B(n_367),
.Y(n_489)
);

BUFx24_ASAP7_75t_SL g533 ( 
.A(n_367),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_479),
.B(n_484),
.Y(n_368)
);

AO21x1_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_468),
.B(n_478),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_442),
.B(n_467),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_405),
.B(n_441),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_385),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_373),
.B(n_385),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_378),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_374),
.A2(n_378),
.B1(n_379),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_396),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_386),
.B(n_397),
.C(n_404),
.Y(n_443)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_403),
.B2(n_404),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_400),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_433),
.B(n_440),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_419),
.B(n_432),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_418),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_415),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_416),
.Y(n_437)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_431),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_431),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_427),
.B(n_430),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_429),
.A2(n_430),
.B(n_459),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_438),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_434),
.B(n_438),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_444),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_457),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_452),
.B2(n_453),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_452),
.C(n_457),
.Y(n_469)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_460),
.Y(n_474)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_469),
.B(n_470),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_472),
.B1(n_475),
.B2(n_477),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_474),
.C(n_477),
.Y(n_480)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_475),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_480),
.B(n_481),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_505),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_504),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_504),
.Y(n_517)
);

BUFx24_ASAP7_75t_SL g534 ( 
.A(n_493),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_497),
.B1(n_499),
.B2(n_503),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_496),
.A2(n_497),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_496),
.B(n_507),
.C(n_511),
.Y(n_523)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_499),
.Y(n_503)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_505),
.A2(n_517),
.B(n_518),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_515),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_515),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_507),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_523),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_523),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_522),
.Y(n_521)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx13_ASAP7_75t_L g530 ( 
.A(n_527),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_531),
.Y(n_528)
);

BUFx12f_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);


endmodule