module fake_jpeg_26065_n_263 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_263);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_23),
.B1(n_17),
.B2(n_21),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_17),
.B1(n_23),
.B2(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_34),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_54),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_17),
.B1(n_23),
.B2(n_21),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_23),
.B1(n_17),
.B2(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_18),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_61),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_56),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_35),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_64),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_60),
.Y(n_81)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_30),
.C(n_34),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_37),
.B1(n_45),
.B2(n_28),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_19),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_37),
.B1(n_27),
.B2(n_45),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_55),
.B(n_51),
.C(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_79),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_69),
.A2(n_72),
.B1(n_58),
.B2(n_59),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_18),
.B(n_19),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_24),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_27),
.B1(n_32),
.B2(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_38),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_20),
.B1(n_14),
.B2(n_15),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_37),
.B1(n_26),
.B2(n_28),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_95),
.B(n_97),
.Y(n_102)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_88),
.B1(n_91),
.B2(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_89),
.Y(n_104)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_67),
.C(n_61),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_77),
.B1(n_72),
.B2(n_82),
.Y(n_111)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_24),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_33),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_101),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_59),
.B1(n_60),
.B2(n_48),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_33),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_76),
.A3(n_70),
.B1(n_78),
.B2(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_110),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_115),
.B1(n_117),
.B2(n_95),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_65),
.B1(n_76),
.B2(n_77),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_116),
.B(n_119),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_81),
.B1(n_66),
.B2(n_65),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_83),
.B(n_65),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_56),
.B(n_54),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_126),
.Y(n_151)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_105),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_110),
.B1(n_108),
.B2(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_134),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_101),
.C(n_99),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_141),
.C(n_129),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_140),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_139),
.A2(n_142),
.B(n_143),
.Y(n_147)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_97),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_33),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_86),
.B(n_91),
.Y(n_142)
);

AO21x1_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_97),
.B(n_91),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_146),
.B1(n_153),
.B2(n_124),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_135),
.A2(n_103),
.B1(n_114),
.B2(n_52),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_73),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_73),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_159),
.B(n_165),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_47),
.Y(n_152)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_32),
.B1(n_25),
.B2(n_51),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_154),
.B(n_164),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_14),
.B(n_20),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_47),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_133),
.C(n_131),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_13),
.C(n_15),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_16),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_75),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_14),
.B(n_20),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_169),
.C(n_181),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_133),
.C(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_162),
.B(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_182),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_165),
.B1(n_159),
.B2(n_75),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_166),
.A2(n_125),
.B1(n_143),
.B2(n_140),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_184),
.B1(n_149),
.B2(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_16),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_125),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_126),
.C(n_62),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_126),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_22),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_185),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_32),
.B1(n_75),
.B2(n_19),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_150),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_154),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_203),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_147),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_173),
.B(n_146),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_197),
.B(n_200),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_147),
.B1(n_157),
.B2(n_158),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_199),
.B1(n_197),
.B2(n_170),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_156),
.B1(n_149),
.B2(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_156),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_187),
.A2(n_168),
.B(n_169),
.C(n_178),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_215),
.C(n_193),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_22),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_167),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_214),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_178),
.C(n_176),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_172),
.B1(n_174),
.B2(n_168),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_191),
.B1(n_176),
.B2(n_184),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_220),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_211),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_183),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_62),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_212),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_62),
.C(n_34),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_227),
.C(n_229),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_237)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_31),
.C(n_75),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_31),
.C(n_22),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_232),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_228),
.A2(n_206),
.B(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_231),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_227),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_22),
.C(n_12),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_0),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_11),
.B(n_10),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_9),
.C(n_7),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_247),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_11),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_232),
.B(n_233),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_249),
.B(n_1),
.Y(n_255)
);

OAI221xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.C(n_7),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_252),
.A2(n_240),
.B1(n_246),
.B2(n_7),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_250),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_256),
.B(n_253),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_4),
.C(n_5),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_6),
.B(n_4),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_261),
.B(n_5),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_6),
.Y(n_263)
);


endmodule