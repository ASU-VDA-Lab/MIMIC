module real_jpeg_23734_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_0),
.B(n_13),
.CON(n_12),
.SN(n_12)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

AO21x1_ASAP7_75t_SL g17 ( 
.A1(n_2),
.A2(n_18),
.B(n_20),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_10),
.Y(n_9)
);

OR2x2_ASAP7_75t_SL g21 ( 
.A(n_3),
.B(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_19),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_25),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_11),
.B1(n_21),
.B2(n_22),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_10),
.B(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_14),
.Y(n_11)
);

BUFx24_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_13),
.B(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_20),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_34),
.Y(n_33)
);

OAI211xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_33),
.C(n_35),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);


endmodule