module fake_netlist_6_3459_n_1844 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1844);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1844;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_1697;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_458;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_924;
wire n_475;
wire n_1582;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_293),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_128),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_187),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_199),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_29),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_90),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_11),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_268),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_39),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_76),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_194),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_54),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_129),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_80),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_81),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_60),
.Y(n_326)
);

BUFx10_ASAP7_75t_L g327 ( 
.A(n_31),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_235),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_88),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_43),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_90),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_214),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_157),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_189),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_104),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_228),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_134),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_195),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_116),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_89),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_80),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_149),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_209),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_117),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_63),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_110),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_146),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_308),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_234),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_223),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_274),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_124),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_206),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_117),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_3),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_273),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_202),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_59),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_12),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_56),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_207),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_211),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_48),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_178),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_87),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_123),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_141),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_253),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_49),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_133),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_140),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_107),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_186),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_56),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_301),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_305),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_255),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_262),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_92),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_198),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_300),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_79),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_87),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_79),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_107),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_115),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_217),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_44),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_24),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_231),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_176),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_192),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_59),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_151),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_38),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_164),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_190),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_208),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_17),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_62),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_32),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_135),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_18),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_246),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_25),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_163),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_219),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_185),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_210),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_98),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_142),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_93),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_62),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_42),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_136),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_71),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_249),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_267),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_31),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_54),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_286),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_131),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_175),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_75),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_184),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_82),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_252),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_240),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_193),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_3),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_27),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_35),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_86),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_7),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_28),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_258),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_125),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_61),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_118),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_283),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_85),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_34),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_147),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_172),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_168),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_113),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_205),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_81),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_157),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_67),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_272),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_285),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_84),
.Y(n_455)
);

BUFx10_ASAP7_75t_L g456 ( 
.A(n_37),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_296),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_4),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_183),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_132),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_73),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_108),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_111),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_250),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_156),
.Y(n_465)
);

BUFx2_ASAP7_75t_SL g466 ( 
.A(n_271),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_30),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_265),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_68),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_139),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_135),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_85),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_196),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_34),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_65),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_11),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_182),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_1),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_241),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_226),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_105),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_19),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_82),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_144),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_74),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_83),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_26),
.Y(n_487)
);

BUFx8_ASAP7_75t_SL g488 ( 
.A(n_276),
.Y(n_488)
);

BUFx10_ASAP7_75t_L g489 ( 
.A(n_39),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_277),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_220),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_248),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_127),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_60),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_4),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_263),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_61),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_218),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_67),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_213),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_55),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_216),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_295),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_95),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_143),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_279),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_91),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_150),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_121),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_307),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_83),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_278),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_188),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_51),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_204),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_177),
.Y(n_516)
);

BUFx5_ASAP7_75t_L g517 ( 
.A(n_181),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_302),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_297),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_45),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_71),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_212),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_47),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_44),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_8),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_159),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_138),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_292),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_149),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_22),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_47),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_109),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_201),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_26),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_104),
.Y(n_535)
);

BUFx5_ASAP7_75t_L g536 ( 
.A(n_215),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_84),
.Y(n_537)
);

BUFx5_ASAP7_75t_L g538 ( 
.A(n_155),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_154),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_114),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_236),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_289),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_256),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_229),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_137),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_18),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_5),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_70),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_294),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_251),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_169),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_122),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_269),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_304),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_166),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_53),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_46),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_33),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_275),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_72),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_367),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_367),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_367),
.B(n_0),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_367),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_309),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_341),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_370),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_449),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_367),
.Y(n_569)
);

INVxp33_ASAP7_75t_SL g570 ( 
.A(n_461),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_422),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_367),
.Y(n_572)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_407),
.B(n_1),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_367),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_367),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_418),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_418),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_366),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_524),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_419),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_418),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_418),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_418),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_418),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_464),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_408),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_418),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_418),
.B(n_2),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_477),
.B(n_2),
.Y(n_589)
);

CKINVDCx16_ASAP7_75t_R g590 ( 
.A(n_379),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_372),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_374),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_518),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_538),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_315),
.B(n_319),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_376),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_384),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_533),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_538),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_385),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_R g602 ( 
.A(n_409),
.B(n_161),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_488),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_538),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g606 ( 
.A(n_345),
.B(n_5),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_538),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_395),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_396),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_403),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_405),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_310),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_333),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_412),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_413),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_512),
.B(n_6),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_417),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_377),
.Y(n_618)
);

INVxp33_ASAP7_75t_SL g619 ( 
.A(n_310),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_333),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_390),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_316),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_378),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_442),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_368),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_487),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_442),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_327),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_487),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_382),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_368),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_357),
.B(n_6),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_534),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_327),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_421),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_327),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_534),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_542),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_368),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_368),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_314),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_426),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_368),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_437),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_434),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_439),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_437),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_437),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_437),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_437),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_394),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_357),
.B(n_7),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_440),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_456),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_483),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_483),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_483),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_542),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_456),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_398),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_483),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_456),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_441),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_483),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_489),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_331),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_313),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_443),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_400),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_444),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_331),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_347),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_347),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_324),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_311),
.B(n_8),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_448),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_311),
.B(n_9),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_314),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_450),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_346),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_406),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_363),
.B(n_9),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_424),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_640),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_661),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_625),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_639),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_640),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_618),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_643),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_623),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_565),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_630),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_625),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_631),
.Y(n_695)
);

INVx6_ASAP7_75t_L g696 ( 
.A(n_595),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_631),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_667),
.B(n_363),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_644),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_624),
.B(n_476),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_581),
.Y(n_701)
);

INVxp67_ASAP7_75t_L g702 ( 
.A(n_571),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_581),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_566),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_647),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_627),
.B(n_392),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_578),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_648),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_649),
.Y(n_709)
);

OA21x2_ASAP7_75t_L g710 ( 
.A1(n_563),
.A2(n_490),
.B(n_392),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_566),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_650),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_651),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_655),
.B(n_490),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_656),
.Y(n_715)
);

XNOR2xp5_ASAP7_75t_L g716 ( 
.A(n_622),
.B(n_343),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_579),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_660),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_638),
.B(n_328),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_582),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_R g721 ( 
.A(n_603),
.B(n_411),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_657),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_669),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_681),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_664),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_582),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_561),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_580),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_585),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_658),
.B(n_335),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_593),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_599),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_613),
.B(n_476),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_674),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_590),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_567),
.B(n_358),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_579),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_620),
.B(n_514),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_662),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_583),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_680),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_586),
.B(n_479),
.Y(n_742)
);

AND2x6_ASAP7_75t_L g743 ( 
.A(n_584),
.B(n_515),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_584),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_591),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_588),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_592),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_562),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_665),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_568),
.B(n_364),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_R g751 ( 
.A(n_597),
.B(n_598),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_621),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_626),
.Y(n_753)
);

OA21x2_ASAP7_75t_L g754 ( 
.A1(n_675),
.A2(n_380),
.B(n_375),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_587),
.Y(n_755)
);

BUFx10_ASAP7_75t_L g756 ( 
.A(n_589),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_629),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_597),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_598),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_587),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_601),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_564),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_633),
.B(n_383),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_594),
.B(n_389),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_601),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_608),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_569),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_594),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_572),
.Y(n_769)
);

OA21x2_ASAP7_75t_L g770 ( 
.A1(n_677),
.A2(n_399),
.B(n_393),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_574),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_575),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_609),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_610),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_616),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_637),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_611),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_576),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_611),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_577),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_666),
.B(n_514),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_604),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_605),
.B(n_410),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_607),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_596),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_596),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_614),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_614),
.B(n_352),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_R g789 ( 
.A(n_615),
.B(n_423),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_746),
.B(n_685),
.Y(n_790)
);

AND2x6_ASAP7_75t_L g791 ( 
.A(n_764),
.B(n_515),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_R g792 ( 
.A(n_751),
.B(n_615),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_743),
.B(n_515),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_764),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_694),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_742),
.B(n_515),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_764),
.B(n_781),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_767),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_735),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_694),
.Y(n_800)
);

BUFx4f_ASAP7_75t_L g801 ( 
.A(n_696),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_696),
.B(n_617),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_778),
.B(n_600),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_767),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_686),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_698),
.B(n_515),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_780),
.B(n_600),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_764),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_696),
.B(n_619),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_696),
.B(n_619),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_697),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_782),
.B(n_632),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_752),
.Y(n_813)
);

OR2x6_ASAP7_75t_L g814 ( 
.A(n_704),
.B(n_628),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_767),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_698),
.A2(n_682),
.B1(n_652),
.B2(n_433),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_753),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_757),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_775),
.B(n_635),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_699),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_699),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_776),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_784),
.B(n_642),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_767),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_700),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_719),
.B(n_642),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_726),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_698),
.B(n_645),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_726),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_686),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_702),
.B(n_612),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_785),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_744),
.B(n_646),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_730),
.B(n_646),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_706),
.B(n_641),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_756),
.B(n_653),
.Y(n_836)
);

AND2x6_ASAP7_75t_L g837 ( 
.A(n_744),
.B(n_420),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_760),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_768),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_736),
.B(n_663),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_785),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_768),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_686),
.Y(n_843)
);

BUFx6f_ASAP7_75t_SL g844 ( 
.A(n_756),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_727),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_733),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_701),
.B(n_703),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_743),
.B(n_517),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_727),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_733),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_734),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_756),
.B(n_663),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_781),
.B(n_666),
.Y(n_853)
);

AO22x2_ASAP7_75t_L g854 ( 
.A1(n_788),
.A2(n_433),
.B1(n_467),
.B2(n_424),
.Y(n_854)
);

BUFx10_ASAP7_75t_L g855 ( 
.A(n_735),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_701),
.B(n_429),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_748),
.Y(n_857)
);

INVx4_ASAP7_75t_SL g858 ( 
.A(n_743),
.Y(n_858)
);

AO21x2_ASAP7_75t_L g859 ( 
.A1(n_783),
.A2(n_602),
.B(n_438),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_762),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_703),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_738),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_686),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_750),
.B(n_668),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_720),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_695),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_762),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_695),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_704),
.B(n_678),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_720),
.B(n_670),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_716),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_789),
.B(n_670),
.Y(n_872)
);

AND2x6_ASAP7_75t_L g873 ( 
.A(n_740),
.B(n_430),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_745),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_769),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_740),
.B(n_676),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_695),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_692),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_740),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_754),
.A2(n_556),
.B1(n_557),
.B2(n_467),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_741),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_755),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_721),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_755),
.Y(n_884)
);

AND2x6_ASAP7_75t_L g885 ( 
.A(n_755),
.B(n_786),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_695),
.Y(n_886)
);

AND2x6_ASAP7_75t_L g887 ( 
.A(n_786),
.B(n_447),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_786),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_771),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_771),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_716),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_777),
.B(n_679),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_743),
.Y(n_893)
);

INVxp33_ASAP7_75t_L g894 ( 
.A(n_738),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_772),
.Y(n_895)
);

OR2x6_ASAP7_75t_L g896 ( 
.A(n_711),
.B(n_634),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_772),
.Y(n_897)
);

CKINVDCx16_ASAP7_75t_R g898 ( 
.A(n_749),
.Y(n_898)
);

AO22x2_ASAP7_75t_L g899 ( 
.A1(n_714),
.A2(n_557),
.B1(n_556),
.B2(n_369),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_684),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_684),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_743),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_754),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_R g904 ( 
.A(n_745),
.B(n_679),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_754),
.A2(n_606),
.B1(n_570),
.B2(n_386),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_687),
.B(n_425),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_777),
.B(n_636),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_690),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_747),
.B(n_654),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_705),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_714),
.B(n_671),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_708),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_714),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_714),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_709),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_689),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_688),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_688),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_712),
.B(n_427),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_754),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_689),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_712),
.Y(n_922)
);

CKINVDCx16_ASAP7_75t_R g923 ( 
.A(n_739),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_SL g924 ( 
.A(n_758),
.B(n_321),
.C(n_318),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_715),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_715),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_722),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_722),
.B(n_431),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_725),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_710),
.Y(n_930)
);

OR2x6_ASAP7_75t_L g931 ( 
.A(n_717),
.B(n_659),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_913),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_801),
.B(n_770),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_825),
.B(n_710),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_825),
.A2(n_761),
.B1(n_765),
.B2(n_759),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_840),
.A2(n_834),
.B1(n_826),
.B2(n_809),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_889),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_802),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_903),
.B(n_710),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_826),
.B(n_759),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_903),
.B(n_710),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_SL g942 ( 
.A(n_883),
.B(n_765),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_880),
.B(n_770),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_834),
.B(n_766),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_L g945 ( 
.A(n_885),
.B(n_766),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_889),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_880),
.B(n_770),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_814),
.B(n_737),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_920),
.B(n_770),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_914),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_876),
.A2(n_763),
.B(n_387),
.C(n_401),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_840),
.B(n_846),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_920),
.B(n_725),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_797),
.B(n_459),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_828),
.Y(n_955)
);

AND2x6_ASAP7_75t_SL g956 ( 
.A(n_931),
.B(n_381),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_797),
.B(n_468),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_869),
.B(n_773),
.Y(n_958)
);

AND2x6_ASAP7_75t_L g959 ( 
.A(n_794),
.B(n_480),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_889),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_878),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_797),
.B(n_491),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_827),
.B(n_829),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_905),
.A2(n_570),
.B1(n_466),
.B2(n_496),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_827),
.B(n_492),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_907),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_914),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_850),
.B(n_774),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_914),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_838),
.B(n_503),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_909),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_839),
.B(n_842),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_794),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_808),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_905),
.A2(n_522),
.B1(n_559),
.B2(n_541),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_808),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_831),
.B(n_779),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_911),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_816),
.A2(n_899),
.B1(n_862),
.B2(n_796),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_879),
.B(n_787),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_862),
.B(n_787),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_861),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_894),
.A2(n_816),
.B(n_812),
.C(n_790),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_930),
.A2(n_672),
.B(n_673),
.C(n_671),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_819),
.B(n_691),
.Y(n_985)
);

INVxp67_ASAP7_75t_SL g986 ( 
.A(n_798),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_819),
.B(n_691),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_861),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_911),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_810),
.A2(n_453),
.B1(n_454),
.B2(n_446),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_865),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_865),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_833),
.B(n_693),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_882),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_795),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_921),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_851),
.B(n_573),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_882),
.B(n_457),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_878),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_881),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_853),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_792),
.B(n_312),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_884),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_884),
.B(n_473),
.Y(n_1004)
);

AND2x6_ASAP7_75t_SL g1005 ( 
.A(n_931),
.B(n_402),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_870),
.B(n_917),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_930),
.B(n_517),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_930),
.B(n_517),
.Y(n_1008)
);

BUFx12f_ASAP7_75t_L g1009 ( 
.A(n_799),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_888),
.B(n_517),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_803),
.B(n_517),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_853),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_807),
.B(n_517),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_883),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_813),
.B(n_672),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_798),
.Y(n_1016)
);

OAI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_835),
.A2(n_373),
.B1(n_388),
.B2(n_323),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_817),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_L g1019 ( 
.A(n_872),
.B(n_707),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_917),
.B(n_517),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_818),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_853),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_800),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_892),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_823),
.B(n_317),
.Y(n_1025)
);

BUFx2_ASAP7_75t_SL g1026 ( 
.A(n_874),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_822),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_798),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_864),
.B(n_320),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_864),
.B(n_713),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_922),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_885),
.B(n_832),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_876),
.B(n_713),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_885),
.B(n_517),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_847),
.A2(n_500),
.B(n_498),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_799),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_926),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_885),
.B(n_536),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_885),
.B(n_536),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_832),
.B(n_536),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_854),
.A2(n_332),
.B1(n_334),
.B2(n_320),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_927),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_814),
.B(n_404),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_872),
.B(n_836),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_929),
.B(n_502),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_841),
.B(n_536),
.Y(n_1046)
);

O2A1O1Ixp5_ASAP7_75t_L g1047 ( 
.A1(n_806),
.A2(n_796),
.B(n_902),
.C(n_893),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_899),
.A2(n_536),
.B1(n_414),
.B2(n_415),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_859),
.A2(n_854),
.B1(n_836),
.B2(n_852),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_SL g1050 ( 
.A1(n_871),
.A2(n_355),
.B1(n_397),
.B2(n_348),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_925),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_852),
.B(n_723),
.C(n_718),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_L g1053 ( 
.A(n_924),
.B(n_452),
.C(n_451),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_859),
.A2(n_506),
.B1(n_334),
.B2(n_337),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_841),
.B(n_536),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_854),
.A2(n_919),
.B1(n_928),
.B2(n_906),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_925),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_L g1058 ( 
.A(n_891),
.B(n_898),
.C(n_923),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_904),
.B(n_339),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_904),
.B(n_344),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_806),
.A2(n_432),
.B(n_435),
.C(n_428),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_908),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_800),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_910),
.B(n_344),
.Y(n_1064)
);

CKINVDCx14_ASAP7_75t_R g1065 ( 
.A(n_799),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_814),
.B(n_445),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_916),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_912),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_900),
.Y(n_1069)
);

OAI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_896),
.A2(n_931),
.B1(n_416),
.B2(n_436),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_915),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_896),
.B(n_855),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_896),
.B(n_724),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_890),
.B(n_349),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_900),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_901),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_837),
.A2(n_351),
.B1(n_354),
.B2(n_350),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_915),
.B(n_728),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_791),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_895),
.B(n_350),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_824),
.A2(n_354),
.B(n_351),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_855),
.B(n_728),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_901),
.B(n_359),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_918),
.B(n_359),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_918),
.B(n_510),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_950),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_974),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_SL g1088 ( 
.A(n_1050),
.B(n_325),
.C(n_322),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_1026),
.B(n_732),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_967),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_961),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_974),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_969),
.Y(n_1093)
);

INVx6_ASAP7_75t_L g1094 ( 
.A(n_982),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_936),
.A2(n_844),
.B1(n_837),
.B2(n_915),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1069),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_983),
.B(n_845),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1044),
.A2(n_1056),
.B1(n_952),
.B2(n_938),
.Y(n_1098)
);

NAND2xp33_ASAP7_75t_SL g1099 ( 
.A(n_975),
.B(n_844),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1075),
.Y(n_1100)
);

BUFx12f_ASAP7_75t_SL g1101 ( 
.A(n_948),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1076),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_974),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_SL g1104 ( 
.A(n_1070),
.B(n_326),
.C(n_325),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_982),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_964),
.A2(n_837),
.B1(n_848),
.B2(n_856),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_982),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_955),
.B(n_849),
.Y(n_1108)
);

OR2x6_ASAP7_75t_L g1109 ( 
.A(n_1009),
.B(n_462),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_966),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_989),
.Y(n_1111)
);

BUFx4f_ASAP7_75t_L g1112 ( 
.A(n_948),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1049),
.A2(n_844),
.B1(n_837),
.B2(n_856),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_999),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1051),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1014),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1065),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_995),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1023),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1006),
.B(n_893),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1057),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_1024),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1063),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_988),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_963),
.B(n_849),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_948),
.B(n_472),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_978),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_958),
.B(n_729),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_L g1129 ( 
.A(n_981),
.B(n_893),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_988),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_997),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1001),
.B(n_858),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_988),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_991),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1031),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_991),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_991),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1071),
.B(n_902),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1037),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_972),
.B(n_1042),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_994),
.B(n_857),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_932),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_994),
.B(n_860),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_992),
.Y(n_1144)
);

NOR3xp33_ASAP7_75t_SL g1145 ( 
.A(n_1017),
.B(n_329),
.C(n_326),
.Y(n_1145)
);

NOR3xp33_ASAP7_75t_SL g1146 ( 
.A(n_1053),
.B(n_330),
.C(n_329),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_937),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1012),
.B(n_858),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_971),
.B(n_855),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_977),
.B(n_729),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_996),
.B(n_731),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_973),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_976),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1022),
.A2(n_873),
.B1(n_887),
.B2(n_856),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_942),
.B(n_731),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1015),
.Y(n_1156)
);

OR2x6_ASAP7_75t_L g1157 ( 
.A(n_1036),
.B(n_474),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_992),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1067),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_997),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_992),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_946),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_979),
.B(n_860),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1015),
.Y(n_1164)
);

OR2x6_ASAP7_75t_L g1165 ( 
.A(n_1082),
.B(n_475),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1000),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_993),
.B(n_489),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_954),
.B(n_867),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_960),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_L g1170 ( 
.A(n_1071),
.B(n_856),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_1003),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_957),
.B(n_867),
.Y(n_1172)
);

NOR3xp33_ASAP7_75t_SL g1173 ( 
.A(n_935),
.B(n_336),
.C(n_330),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1043),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_1003),
.Y(n_1175)
);

BUFx12f_ASAP7_75t_L g1176 ( 
.A(n_956),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1003),
.Y(n_1177)
);

INVx5_ASAP7_75t_L g1178 ( 
.A(n_959),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_943),
.A2(n_504),
.B(n_511),
.C(n_501),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1018),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1048),
.A2(n_887),
.B1(n_873),
.B2(n_539),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1043),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1071),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1016),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_962),
.B(n_875),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_959),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1021),
.B(n_875),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_953),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_953),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1027),
.B(n_897),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_984),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1078),
.Y(n_1192)
);

AO22x1_ASAP7_75t_L g1193 ( 
.A1(n_985),
.A2(n_338),
.B1(n_340),
.B2(n_336),
.Y(n_1193)
);

NOR3xp33_ASAP7_75t_SL g1194 ( 
.A(n_1041),
.B(n_340),
.C(n_338),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_940),
.A2(n_944),
.B1(n_1033),
.B2(n_1030),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1043),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1062),
.B(n_897),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1068),
.B(n_805),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1016),
.Y(n_1199)
);

INVxp33_ASAP7_75t_L g1200 ( 
.A(n_1073),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1040),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1066),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1072),
.B(n_805),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1040),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_980),
.B(n_805),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_934),
.A2(n_887),
.B1(n_873),
.B2(n_540),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1083),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1079),
.B(n_1032),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1066),
.Y(n_1209)
);

NOR3xp33_ASAP7_75t_SL g1210 ( 
.A(n_987),
.B(n_353),
.C(n_342),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1010),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1046),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1207),
.B(n_1083),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1207),
.B(n_1084),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1120),
.A2(n_941),
.B(n_939),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1097),
.A2(n_1008),
.B(n_1007),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1132),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1192),
.B(n_1085),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1135),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1140),
.B(n_1085),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1120),
.A2(n_941),
.B(n_939),
.Y(n_1221)
);

CKINVDCx16_ASAP7_75t_R g1222 ( 
.A(n_1155),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1188),
.B(n_1189),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1114),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1203),
.B(n_1019),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1086),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1211),
.B(n_949),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1139),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1091),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1191),
.A2(n_1008),
.B(n_1007),
.Y(n_1230)
);

AOI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1163),
.A2(n_949),
.B(n_1208),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1116),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1191),
.A2(n_1047),
.B(n_1020),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1155),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1132),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1195),
.B(n_1098),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1179),
.A2(n_947),
.B(n_943),
.C(n_951),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1208),
.A2(n_1020),
.B(n_933),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1204),
.B(n_1212),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1200),
.B(n_968),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_SL g1241 ( 
.A1(n_1179),
.A2(n_947),
.B(n_1029),
.C(n_1034),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1095),
.A2(n_933),
.B1(n_1032),
.B2(n_1054),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1159),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1204),
.B(n_1080),
.Y(n_1244)
);

AOI221x1_ASAP7_75t_L g1245 ( 
.A1(n_1099),
.A2(n_1035),
.B1(n_1011),
.B2(n_1013),
.C(n_970),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1184),
.A2(n_1028),
.B(n_1079),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1086),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1114),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1184),
.A2(n_1028),
.B(n_1079),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1212),
.B(n_965),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1148),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1117),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1158),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1148),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1151),
.Y(n_1255)
);

NOR4xp25_ASAP7_75t_L g1256 ( 
.A(n_1167),
.B(n_1025),
.C(n_1061),
.D(n_1060),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1108),
.B(n_1045),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1201),
.B(n_1064),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1166),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1199),
.A2(n_1079),
.B(n_986),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1138),
.A2(n_945),
.B(n_998),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1180),
.B(n_1002),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1138),
.A2(n_1093),
.B(n_1090),
.Y(n_1263)
);

OAI21xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1106),
.A2(n_1038),
.B(n_1034),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1113),
.A2(n_1039),
.B(n_1038),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_L g1266 ( 
.A(n_1145),
.B(n_1052),
.C(n_990),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1168),
.A2(n_1185),
.A3(n_1172),
.B(n_1205),
.Y(n_1267)
);

AO32x2_ASAP7_75t_L g1268 ( 
.A1(n_1130),
.A2(n_863),
.A3(n_843),
.B1(n_959),
.B2(n_1039),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1090),
.A2(n_1055),
.B(n_868),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1127),
.B(n_1074),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1093),
.A2(n_868),
.B(n_866),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1206),
.A2(n_1004),
.B(n_815),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1206),
.A2(n_815),
.B(n_804),
.Y(n_1273)
);

OAI21xp33_ASAP7_75t_L g1274 ( 
.A1(n_1145),
.A2(n_1059),
.B(n_482),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1187),
.B(n_959),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1141),
.A2(n_868),
.B(n_866),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1158),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1125),
.A2(n_820),
.A3(n_821),
.B(n_811),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1096),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1239),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_1232),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1264),
.A2(n_1129),
.B(n_1181),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1223),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1217),
.B(n_1203),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1220),
.B(n_1122),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1217),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1276),
.A2(n_1198),
.B(n_1143),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1236),
.A2(n_1181),
.B(n_1106),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1213),
.B(n_1156),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1214),
.B(n_1164),
.Y(n_1290)
);

OA21x2_ASAP7_75t_L g1291 ( 
.A1(n_1245),
.A2(n_1197),
.B(n_1190),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1232),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_SL g1293 ( 
.A1(n_1265),
.A2(n_1154),
.B(n_1102),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1226),
.Y(n_1294)
);

BUFx8_ASAP7_75t_L g1295 ( 
.A(n_1229),
.Y(n_1295)
);

BUFx4_ASAP7_75t_R g1296 ( 
.A(n_1224),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1247),
.Y(n_1297)
);

AO32x2_ASAP7_75t_L g1298 ( 
.A1(n_1242),
.A2(n_1130),
.A3(n_1175),
.B1(n_1171),
.B2(n_1209),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_SL g1299 ( 
.A1(n_1231),
.A2(n_1261),
.B(n_1221),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1247),
.Y(n_1300)
);

INVx6_ASAP7_75t_L g1301 ( 
.A(n_1224),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1276),
.A2(n_1115),
.B(n_1100),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1274),
.A2(n_1150),
.B(n_1128),
.C(n_1104),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1237),
.A2(n_1121),
.A3(n_1162),
.B(n_1147),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1230),
.A2(n_1162),
.B(n_1147),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1218),
.B(n_1110),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1240),
.A2(n_1088),
.B1(n_1165),
.B2(n_1149),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1237),
.A2(n_1169),
.A3(n_1119),
.B(n_1123),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1266),
.A2(n_1104),
.B(n_1088),
.C(n_1173),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1255),
.B(n_1165),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1217),
.B(n_1177),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1248),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1230),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1235),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1235),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1269),
.A2(n_1169),
.B(n_1119),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1227),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1244),
.B(n_1194),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1257),
.A2(n_1152),
.B(n_1142),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1253),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1229),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1295),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1286),
.B(n_1263),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1286),
.B(n_1263),
.Y(n_1324)
);

BUFx12f_ASAP7_75t_L g1325 ( 
.A(n_1292),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1308),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1305),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1318),
.A2(n_1058),
.B1(n_1165),
.B2(n_1225),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1304),
.B(n_1267),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1288),
.A2(n_1256),
.B(n_1272),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1305),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_SL g1332 ( 
.A(n_1303),
.B(n_1210),
.C(n_1146),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1304),
.B(n_1267),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1282),
.A2(n_1215),
.B(n_1241),
.Y(n_1334)
);

NAND2x1_ASAP7_75t_L g1335 ( 
.A(n_1293),
.B(n_1183),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1289),
.A2(n_1279),
.B1(n_1228),
.B2(n_1259),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1305),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1305),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1280),
.B(n_1267),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1304),
.B(n_1267),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1285),
.A2(n_1222),
.B1(n_495),
.B2(n_505),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1292),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1307),
.A2(n_494),
.B1(n_535),
.B2(n_507),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1307),
.A2(n_1290),
.B1(n_1089),
.B2(n_1270),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1299),
.A2(n_1241),
.B(n_1273),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1308),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1308),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1295),
.A2(n_1234),
.B1(n_1089),
.B2(n_1176),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_L g1349 ( 
.A1(n_1309),
.A2(n_1193),
.B1(n_525),
.B2(n_391),
.C(n_545),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1283),
.B(n_1250),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1281),
.Y(n_1351)
);

BUFx10_ASAP7_75t_L g1352 ( 
.A(n_1306),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1304),
.B(n_1268),
.Y(n_1353)
);

INVx4_ASAP7_75t_L g1354 ( 
.A(n_1296),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_SL g1355 ( 
.A(n_1319),
.B(n_1210),
.C(n_1146),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1284),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1310),
.A2(n_1089),
.B1(n_1202),
.B2(n_1182),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1293),
.A2(n_1202),
.B1(n_1182),
.B2(n_1112),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1295),
.A2(n_1234),
.B1(n_537),
.B2(n_1112),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1321),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1308),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1317),
.A2(n_1219),
.B1(n_1262),
.B2(n_1258),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1304),
.B(n_1308),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1339),
.B(n_1313),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1334),
.A2(n_1317),
.A3(n_1298),
.B(n_1268),
.Y(n_1365)
);

AO22x1_ASAP7_75t_L g1366 ( 
.A1(n_1354),
.A2(n_1252),
.B1(n_353),
.B2(n_356),
.Y(n_1366)
);

INVx4_ASAP7_75t_L g1367 ( 
.A(n_1354),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1330),
.A2(n_1287),
.B(n_1316),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1363),
.B(n_1298),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1330),
.A2(n_1186),
.B(n_1178),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1354),
.A2(n_1349),
.B1(n_1344),
.B2(n_1332),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1345),
.A2(n_1316),
.B(n_1269),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1350),
.A2(n_1186),
.B(n_1178),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1355),
.A2(n_1126),
.B1(n_1284),
.B2(n_1157),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1363),
.B(n_1298),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1356),
.Y(n_1376)
);

AOI33xp33_ASAP7_75t_L g1377 ( 
.A1(n_1343),
.A2(n_1243),
.A3(n_673),
.B1(n_683),
.B2(n_1160),
.B3(n_1131),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1355),
.A2(n_1126),
.B1(n_1284),
.B2(n_1196),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1326),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1363),
.B(n_1298),
.Y(n_1380)
);

BUFx4f_ASAP7_75t_SL g1381 ( 
.A(n_1325),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1329),
.B(n_1291),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1349),
.A2(n_1174),
.B(n_1109),
.C(n_1275),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1341),
.A2(n_352),
.B1(n_516),
.B2(n_959),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1345),
.A2(n_1186),
.B(n_1178),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1329),
.B(n_1333),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1328),
.A2(n_516),
.B1(n_1101),
.B2(n_1311),
.Y(n_1387)
);

OAI321xp33_ASAP7_75t_L g1388 ( 
.A1(n_1362),
.A2(n_1077),
.A3(n_1109),
.B1(n_1153),
.B2(n_1297),
.C(n_1320),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1329),
.B(n_1298),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1333),
.B(n_1298),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1327),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1360),
.Y(n_1392)
);

AOI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1362),
.A2(n_460),
.B1(n_463),
.B2(n_458),
.C(n_455),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1359),
.A2(n_1312),
.B1(n_1301),
.B2(n_1248),
.Y(n_1394)
);

CKINVDCx14_ASAP7_75t_R g1395 ( 
.A(n_1351),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1342),
.Y(n_1396)
);

OAI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1357),
.A2(n_362),
.B1(n_365),
.B2(n_361),
.C(n_360),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1352),
.A2(n_1311),
.B1(n_1314),
.B2(n_1286),
.Y(n_1398)
);

OAI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1358),
.A2(n_365),
.B1(n_371),
.B2(n_361),
.C(n_360),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1352),
.A2(n_1311),
.B1(n_1315),
.B2(n_1314),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1322),
.A2(n_1186),
.B1(n_1087),
.B2(n_1314),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1340),
.B(n_1294),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1336),
.B(n_1294),
.Y(n_1403)
);

NOR2x1_ASAP7_75t_SL g1404 ( 
.A(n_1322),
.B(n_1287),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1335),
.A2(n_1170),
.B(n_1216),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1323),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1348),
.A2(n_1253),
.B1(n_1277),
.B2(n_1177),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1340),
.B(n_1300),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1348),
.A2(n_1315),
.B1(n_537),
.B2(n_1133),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1323),
.A2(n_1094),
.B1(n_465),
.B2(n_469),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1346),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1323),
.A2(n_1315),
.B1(n_1133),
.B2(n_1111),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1323),
.A2(n_1175),
.B1(n_1171),
.B2(n_1235),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1327),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1331),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1353),
.B(n_1291),
.Y(n_1416)
);

AND3x1_ASAP7_75t_L g1417 ( 
.A(n_1384),
.B(n_683),
.C(n_1005),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1391),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1379),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1371),
.B(n_1324),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1386),
.B(n_1369),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1386),
.B(n_1346),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1391),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1369),
.B(n_1347),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1375),
.B(n_1347),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1402),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1414),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1392),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1375),
.B(n_1347),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1367),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1380),
.B(n_1361),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1370),
.A2(n_1103),
.B(n_1092),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1376),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1406),
.B(n_1324),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1380),
.B(n_1361),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1389),
.B(n_1361),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1405),
.A2(n_1331),
.B(n_1287),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1402),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1408),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1408),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1382),
.B(n_1337),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1396),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1415),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1389),
.B(n_1337),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1364),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1406),
.B(n_1337),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1364),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1411),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1390),
.B(n_1338),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1366),
.B(n_510),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1338),
.Y(n_1451)
);

AO21x2_ASAP7_75t_L g1452 ( 
.A1(n_1372),
.A2(n_1271),
.B(n_1216),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1416),
.B(n_1268),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1404),
.B(n_1278),
.Y(n_1454)
);

OR2x6_ASAP7_75t_L g1455 ( 
.A(n_1367),
.B(n_1302),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1365),
.Y(n_1456)
);

NOR2x1_ASAP7_75t_L g1457 ( 
.A(n_1367),
.B(n_1302),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1365),
.Y(n_1458)
);

AO31x2_ASAP7_75t_L g1459 ( 
.A1(n_1385),
.A2(n_1260),
.A3(n_1249),
.B(n_1246),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1403),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1368),
.B(n_1302),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1365),
.B(n_1302),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1368),
.B(n_1278),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1372),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1383),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1398),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1400),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1376),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1376),
.Y(n_1469)
);

INVx3_ASAP7_75t_SL g1470 ( 
.A(n_1381),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1413),
.B(n_1278),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1394),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1399),
.A2(n_521),
.B1(n_523),
.B2(n_520),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1388),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1407),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1410),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1377),
.B(n_470),
.Y(n_1477)
);

NOR2x1_ASAP7_75t_SL g1478 ( 
.A(n_1401),
.B(n_1092),
.Y(n_1478)
);

BUFx2_ASAP7_75t_SL g1479 ( 
.A(n_1373),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1412),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1378),
.Y(n_1481)
);

OR2x6_ASAP7_75t_L g1482 ( 
.A(n_1374),
.B(n_1238),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1409),
.B(n_1233),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1393),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1397),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1387),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1379),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1391),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1392),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1406),
.B(n_1271),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1392),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1391),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1371),
.A2(n_478),
.B1(n_481),
.B2(n_471),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1386),
.B(n_10),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1391),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1392),
.Y(n_1496)
);

A2O1A1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1383),
.A2(n_519),
.B(n_528),
.C(n_513),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1379),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1395),
.B(n_513),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1379),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1379),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1379),
.Y(n_1502)
);

INVx8_ASAP7_75t_L g1503 ( 
.A(n_1376),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1386),
.B(n_13),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1484),
.A2(n_521),
.B1(n_523),
.B2(n_520),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1484),
.B(n_1493),
.C(n_1465),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1475),
.A2(n_527),
.B1(n_529),
.B2(n_526),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1419),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1470),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1474),
.A2(n_531),
.B1(n_532),
.B2(n_530),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1485),
.A2(n_547),
.B1(n_548),
.B2(n_546),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1421),
.B(n_14),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1497),
.B(n_558),
.C(n_552),
.Y(n_1513)
);

CKINVDCx14_ASAP7_75t_R g1514 ( 
.A(n_1442),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1485),
.A2(n_1417),
.B1(n_1476),
.B2(n_1473),
.C(n_1450),
.Y(n_1515)
);

NAND2xp33_ASAP7_75t_R g1516 ( 
.A(n_1475),
.B(n_15),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1428),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1460),
.B(n_484),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1486),
.A2(n_560),
.B1(n_486),
.B2(n_493),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1487),
.Y(n_1520)
);

AO21x2_ASAP7_75t_L g1521 ( 
.A1(n_1464),
.A2(n_1081),
.B(n_1118),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1468),
.B(n_16),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1481),
.A2(n_497),
.B1(n_499),
.B2(n_485),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1433),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1434),
.B(n_1105),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1441),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1498),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1472),
.A2(n_509),
.B1(n_508),
.B2(n_519),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1470),
.Y(n_1529)
);

AND2x6_ASAP7_75t_L g1530 ( 
.A(n_1430),
.B(n_1254),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1500),
.Y(n_1531)
);

AOI222xp33_ASAP7_75t_L g1532 ( 
.A1(n_1477),
.A2(n_555),
.B1(n_554),
.B2(n_553),
.C1(n_551),
.C2(n_550),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1466),
.A2(n_1467),
.B1(n_1420),
.B2(n_1480),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1434),
.B(n_1105),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1422),
.B(n_20),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1420),
.A2(n_544),
.B1(n_549),
.B2(n_543),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1503),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1501),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1433),
.Y(n_1540)
);

NAND4xp25_ASAP7_75t_L g1541 ( 
.A(n_1499),
.B(n_24),
.C(n_21),
.D(n_23),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1445),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1447),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1489),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1480),
.A2(n_1094),
.B1(n_1103),
.B2(n_1092),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1418),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1469),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1491),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1496),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1461),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1432),
.A2(n_1103),
.B(n_793),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1503),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1456),
.A2(n_1458),
.B(n_1462),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1480),
.B(n_1107),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1418),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1418),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1426),
.B(n_36),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_L g1558 ( 
.A(n_1432),
.B(n_1107),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1488),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1438),
.B(n_1439),
.Y(n_1560)
);

CKINVDCx12_ASAP7_75t_R g1561 ( 
.A(n_1494),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1495),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1440),
.B(n_36),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1434),
.B(n_1436),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1480),
.A2(n_1124),
.B1(n_1134),
.B2(n_1107),
.Y(n_1565)
);

INVx5_ASAP7_75t_L g1566 ( 
.A(n_1455),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1423),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1446),
.B(n_1124),
.Y(n_1568)
);

NAND3xp33_ASAP7_75t_SL g1569 ( 
.A(n_1504),
.B(n_40),
.C(n_41),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1482),
.A2(n_1251),
.B1(n_1254),
.B2(n_1136),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1446),
.B(n_1134),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1508),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1533),
.B(n_1430),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1546),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1564),
.B(n_1444),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1572),
.B(n_1526),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1526),
.B(n_1444),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1566),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1566),
.B(n_1455),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1520),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1546),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1553),
.B(n_1449),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1566),
.B(n_1524),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1449),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1527),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1517),
.B(n_1451),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1544),
.B(n_1425),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1548),
.B(n_1429),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1549),
.B(n_1429),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1524),
.B(n_1455),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1531),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1509),
.B(n_1430),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1529),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1550),
.B(n_1431),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1538),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1550),
.B(n_1431),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1539),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1560),
.B(n_1435),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1559),
.B(n_1435),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1562),
.B(n_1453),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1555),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1556),
.B(n_1462),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1558),
.B(n_1457),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1567),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1540),
.B(n_1454),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1547),
.B(n_1463),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1568),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1568),
.B(n_1571),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1525),
.B(n_1448),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1512),
.B(n_1463),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1561),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1563),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1533),
.B(n_1483),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1521),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1535),
.B(n_1427),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1506),
.A2(n_1479),
.B1(n_1483),
.B2(n_1471),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1557),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1522),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1534),
.B(n_1448),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1554),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1570),
.B(n_1443),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1518),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1537),
.B(n_1443),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1569),
.B(n_1492),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1552),
.B(n_1479),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1530),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1530),
.B(n_1490),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1514),
.B(n_1437),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1514),
.B(n_1437),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1583),
.B(n_1478),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1573),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1595),
.Y(n_1634)
);

OAI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1574),
.A2(n_1505),
.B1(n_1516),
.B2(n_1536),
.C(n_1523),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1610),
.B(n_1577),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1584),
.Y(n_1637)
);

OR2x2_ASAP7_75t_SL g1638 ( 
.A(n_1613),
.B(n_1513),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1610),
.B(n_1530),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1575),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1581),
.Y(n_1641)
);

OAI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1615),
.A2(n_1505),
.B1(n_1523),
.B2(n_1507),
.C(n_1541),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1626),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1582),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1624),
.B(n_1515),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1577),
.B(n_1459),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1576),
.B(n_1459),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1614),
.B(n_1532),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1576),
.B(n_1452),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1617),
.B(n_1452),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1586),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1592),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1597),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1626),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1612),
.B(n_1565),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1599),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1585),
.B(n_1545),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1630),
.B(n_1551),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1594),
.Y(n_1659)
);

NAND3xp33_ASAP7_75t_L g1660 ( 
.A(n_1618),
.B(n_1511),
.C(n_1528),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1622),
.B(n_1510),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1606),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1608),
.B(n_1519),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1608),
.B(n_46),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1606),
.Y(n_1665)
);

NOR2xp67_ASAP7_75t_L g1666 ( 
.A(n_1579),
.B(n_1584),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1578),
.B(n_50),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1584),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1605),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1604),
.Y(n_1670)
);

NAND2x1p5_ASAP7_75t_L g1671 ( 
.A(n_1579),
.B(n_1628),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1601),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1631),
.B(n_52),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1596),
.B(n_53),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1596),
.B(n_55),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1588),
.Y(n_1676)
);

INVx3_ASAP7_75t_SL g1677 ( 
.A(n_1595),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1633),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1643),
.B(n_1598),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1645),
.B(n_1593),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1636),
.B(n_1609),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1677),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1654),
.B(n_1620),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1641),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1634),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1639),
.B(n_1607),
.Y(n_1686)
);

NOR3xp33_ASAP7_75t_L g1687 ( 
.A(n_1635),
.B(n_1660),
.C(n_1642),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1659),
.B(n_1600),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1637),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1673),
.B(n_1651),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1655),
.B(n_1607),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1652),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1653),
.B(n_1602),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1648),
.B(n_1619),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1637),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1656),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1637),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1668),
.B(n_1591),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1644),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1657),
.B(n_1589),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1674),
.B(n_1602),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1666),
.B(n_1580),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1675),
.B(n_1669),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1662),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1676),
.B(n_1587),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1671),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1665),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1672),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1664),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1663),
.B(n_1590),
.Y(n_1710)
);

OAI211xp5_ASAP7_75t_L g1711 ( 
.A1(n_1661),
.A2(n_1627),
.B(n_1623),
.C(n_1616),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1638),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1658),
.B(n_1611),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1678),
.Y(n_1714)
);

NAND2x1p5_ASAP7_75t_L g1715 ( 
.A(n_1685),
.B(n_1667),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1682),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1691),
.B(n_1632),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1698),
.Y(n_1718)
);

AOI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1712),
.A2(n_1650),
.B(n_1640),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1684),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1687),
.A2(n_1647),
.B1(n_1646),
.B2(n_1629),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1686),
.B(n_1670),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1694),
.B(n_1649),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1692),
.Y(n_1724)
);

INVxp33_ASAP7_75t_L g1725 ( 
.A(n_1680),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1703),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1696),
.Y(n_1727)
);

AO22x2_ASAP7_75t_L g1728 ( 
.A1(n_1711),
.A2(n_1603),
.B1(n_1621),
.B2(n_1625),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1702),
.B(n_1706),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1690),
.A2(n_1144),
.B(n_1137),
.Y(n_1730)
);

OAI322xp33_ASAP7_75t_L g1731 ( 
.A1(n_1699),
.A2(n_57),
.A3(n_58),
.B1(n_63),
.B2(n_64),
.C1(n_65),
.C2(n_66),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1710),
.B(n_57),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1690),
.B(n_64),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1689),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1709),
.B(n_69),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1695),
.A2(n_77),
.B(n_78),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1713),
.B(n_1700),
.Y(n_1737)
);

OR2x6_ASAP7_75t_L g1738 ( 
.A(n_1697),
.B(n_1161),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1683),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1716),
.B(n_1701),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1725),
.A2(n_1679),
.B(n_1704),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1736),
.Y(n_1742)
);

NOR2x1_ASAP7_75t_L g1743 ( 
.A(n_1736),
.B(n_1707),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1729),
.B(n_1737),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1714),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1726),
.B(n_1708),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1735),
.B(n_1688),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1729),
.B(n_1681),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1733),
.B(n_1705),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1715),
.B(n_1693),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1732),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1717),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1720),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1738),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1724),
.Y(n_1755)
);

AOI211xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1731),
.A2(n_94),
.B(n_96),
.C(n_97),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1739),
.B(n_97),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1727),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1719),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.C(n_102),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1718),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1734),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1751),
.B(n_1722),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1742),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1745),
.Y(n_1764)
);

XNOR2x2_ASAP7_75t_L g1765 ( 
.A(n_1742),
.B(n_1728),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1744),
.B(n_1721),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1756),
.B(n_1730),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1743),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1748),
.B(n_1723),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1760),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1753),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1755),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1749),
.B(n_101),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1758),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1760),
.B(n_103),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1752),
.B(n_106),
.Y(n_1776)
);

NOR3xp33_ASAP7_75t_SL g1777 ( 
.A(n_1759),
.B(n_1740),
.C(n_1757),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1746),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1768),
.B(n_1741),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1776),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1763),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1770),
.Y(n_1782)
);

AND4x1_ASAP7_75t_L g1783 ( 
.A(n_1777),
.B(n_1747),
.C(n_1761),
.D(n_1750),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1766),
.B(n_1754),
.Y(n_1784)
);

AOI211xp5_ASAP7_75t_L g1785 ( 
.A1(n_1767),
.A2(n_111),
.B(n_112),
.C(n_113),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1769),
.B(n_116),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1770),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1762),
.Y(n_1788)
);

NOR2x1_ASAP7_75t_L g1789 ( 
.A(n_1775),
.B(n_119),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1765),
.Y(n_1790)
);

AOI221x1_ASAP7_75t_L g1791 ( 
.A1(n_1773),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.C(n_123),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1778),
.B(n_124),
.Y(n_1792)
);

OAI33xp33_ASAP7_75t_L g1793 ( 
.A1(n_1764),
.A2(n_126),
.A3(n_127),
.B1(n_128),
.B2(n_129),
.B3(n_130),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1778),
.B(n_126),
.Y(n_1794)
);

NOR4xp25_ASAP7_75t_L g1795 ( 
.A(n_1790),
.B(n_1771),
.C(n_1774),
.D(n_1772),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1781),
.Y(n_1796)
);

AOI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1779),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.C(n_147),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1784),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1789),
.Y(n_1799)
);

OAI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1791),
.A2(n_145),
.B(n_148),
.C(n_150),
.Y(n_1800)
);

NAND4xp25_ASAP7_75t_SL g1801 ( 
.A(n_1785),
.B(n_148),
.C(n_151),
.D(n_152),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1788),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.C(n_158),
.Y(n_1802)
);

NOR3xp33_ASAP7_75t_L g1803 ( 
.A(n_1780),
.B(n_153),
.C(n_159),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1783),
.A2(n_160),
.B1(n_811),
.B2(n_162),
.C(n_165),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1786),
.A2(n_887),
.B1(n_873),
.B2(n_791),
.Y(n_1805)
);

AOI211x1_ASAP7_75t_L g1806 ( 
.A1(n_1792),
.A2(n_167),
.B(n_170),
.C(n_171),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1782),
.A2(n_173),
.B1(n_174),
.B2(n_179),
.C(n_180),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1787),
.A2(n_791),
.B1(n_866),
.B2(n_877),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1793),
.A2(n_191),
.B1(n_197),
.B2(n_200),
.C(n_203),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_R g1810 ( 
.A(n_1801),
.B(n_1794),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1798),
.B(n_221),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_R g1812 ( 
.A(n_1799),
.B(n_222),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1796),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1795),
.B(n_224),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1804),
.A2(n_225),
.B1(n_227),
.B2(n_230),
.C(n_232),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1803),
.B(n_233),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1800),
.B(n_804),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_SL g1818 ( 
.A(n_1809),
.B(n_237),
.C(n_238),
.Y(n_1818)
);

NAND4xp75_ASAP7_75t_L g1819 ( 
.A(n_1814),
.B(n_1797),
.C(n_1802),
.D(n_1806),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1813),
.B(n_1805),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1812),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1816),
.B(n_1808),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1811),
.Y(n_1823)
);

NAND4xp75_ASAP7_75t_L g1824 ( 
.A(n_1817),
.B(n_1807),
.C(n_242),
.D(n_243),
.Y(n_1824)
);

INVx4_ASAP7_75t_L g1825 ( 
.A(n_1816),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1818),
.B(n_239),
.Y(n_1826)
);

NOR3xp33_ASAP7_75t_L g1827 ( 
.A(n_1825),
.B(n_1815),
.C(n_1810),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1821),
.A2(n_791),
.B1(n_245),
.B2(n_247),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1823),
.Y(n_1829)
);

NAND5xp2_ASAP7_75t_L g1830 ( 
.A(n_1822),
.B(n_244),
.C(n_254),
.D(n_257),
.E(n_259),
.Y(n_1830)
);

NAND3xp33_ASAP7_75t_SL g1831 ( 
.A(n_1826),
.B(n_260),
.C(n_261),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1829),
.B(n_1820),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1827),
.B(n_1819),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1831),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1832),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1833),
.B(n_1824),
.Y(n_1836)
);

XNOR2x1_ASAP7_75t_L g1837 ( 
.A(n_1836),
.B(n_1834),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1835),
.B(n_1828),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1837),
.Y(n_1839)
);

AND3x1_ASAP7_75t_L g1840 ( 
.A(n_1839),
.B(n_1838),
.C(n_1830),
.Y(n_1840)
);

OAI222xp33_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_264),
.B1(n_270),
.B2(n_280),
.C1(n_281),
.C2(n_282),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_830),
.B1(n_886),
.B2(n_877),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_284),
.B1(n_287),
.B2(n_288),
.C(n_291),
.Y(n_1843)
);

AOI211xp5_ASAP7_75t_L g1844 ( 
.A1(n_1843),
.A2(n_298),
.B(n_303),
.C(n_306),
.Y(n_1844)
);


endmodule