module fake_jpeg_8179_n_101 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx8_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_0),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_56),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_0),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_15),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_61),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_67),
.B1(n_20),
.B2(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_53),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_45),
.B1(n_39),
.B2(n_3),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_68),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_1),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_43),
.B1(n_3),
.B2(n_4),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_12),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_14),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx2_ASAP7_75t_SL g77 ( 
.A(n_74),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_75),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_79),
.B1(n_85),
.B2(n_75),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_22),
.A3(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_83),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_86),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_80),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_82),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_83),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_78),
.B1(n_81),
.B2(n_77),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_59),
.C(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

OAI21x1_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_26),
.B(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_30),
.Y(n_101)
);


endmodule