module fake_jpeg_1603_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_47),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_62),
.Y(n_91)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_63),
.Y(n_95)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_53),
.Y(n_130)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_1),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_69),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_2),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_76),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_17),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_3),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_80),
.Y(n_133)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_23),
.B(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_82),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_36),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_87),
.B(n_36),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_4),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_25),
.B(n_4),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_43),
.B1(n_33),
.B2(n_44),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_90),
.A2(n_92),
.B1(n_113),
.B2(n_114),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_43),
.B1(n_45),
.B2(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_54),
.B(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_101),
.B(n_115),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_58),
.A2(n_24),
.B1(n_35),
.B2(n_29),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_65),
.A2(n_28),
.B1(n_35),
.B2(n_45),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_40),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_34),
.B1(n_32),
.B2(n_36),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_68),
.B(n_26),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_47),
.B(n_34),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_47),
.B(n_32),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_129),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_57),
.A2(n_66),
.B1(n_59),
.B2(n_68),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_135),
.B1(n_113),
.B2(n_114),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_59),
.A2(n_36),
.B(n_7),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_131),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_26),
.C(n_11),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_71),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_82),
.C(n_81),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_6),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_66),
.A2(n_26),
.B1(n_12),
.B2(n_14),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_77),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_141),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_143),
.A2(n_158),
.B(n_170),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_144),
.Y(n_208)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

BUFx4f_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_165),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_84),
.B1(n_60),
.B2(n_73),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_160),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_6),
.B(n_12),
.C(n_14),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_143),
.B(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_6),
.B1(n_12),
.B2(n_130),
.Y(n_158)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_95),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_108),
.B(n_125),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_91),
.B(n_100),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_176),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_135),
.B1(n_109),
.B2(n_107),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_175),
.B1(n_181),
.B2(n_123),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_121),
.B1(n_98),
.B2(n_103),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_123),
.B1(n_110),
.B2(n_99),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_107),
.A2(n_109),
.B1(n_93),
.B2(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_103),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_178),
.Y(n_212)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_93),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_180),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_98),
.A2(n_99),
.B1(n_112),
.B2(n_110),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_191),
.C(n_192),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_187),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_155),
.B1(n_170),
.B2(n_140),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_194),
.A2(n_197),
.B1(n_205),
.B2(n_207),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_147),
.B(n_174),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_148),
.B1(n_150),
.B2(n_164),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_151),
.B1(n_162),
.B2(n_157),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_154),
.B1(n_146),
.B2(n_174),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_147),
.A2(n_174),
.B(n_176),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_168),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_215),
.B(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_142),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_169),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_172),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_184),
.B(n_145),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_198),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_202),
.B(n_188),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_198),
.B1(n_191),
.B2(n_204),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_230),
.B1(n_235),
.B2(n_209),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_167),
.B1(n_166),
.B2(n_179),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_232),
.Y(n_239)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_184),
.B(n_159),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_234),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_205),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_198),
.B1(n_207),
.B2(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_193),
.Y(n_253)
);

XNOR2x2_ASAP7_75t_SL g240 ( 
.A(n_227),
.B(n_212),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_221),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_250),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_206),
.C(n_213),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_244),
.C(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_206),
.C(n_190),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_211),
.A3(n_210),
.B1(n_183),
.B2(n_185),
.C1(n_186),
.C2(n_208),
.Y(n_247)
);

OAI322xp33_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_225),
.A3(n_235),
.B1(n_219),
.B2(n_214),
.C1(n_216),
.C2(n_220),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_202),
.C(n_185),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_221),
.B1(n_225),
.B2(n_223),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_250),
.B1(n_253),
.B2(n_211),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_258),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_SL g272 ( 
.A(n_257),
.B(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_245),
.B(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_225),
.B1(n_222),
.B2(n_236),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_261),
.A2(n_251),
.B1(n_237),
.B2(n_241),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_232),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_265),
.C(n_266),
.Y(n_267)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_239),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_230),
.C(n_193),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_252),
.C(n_238),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_274),
.B1(n_276),
.B2(n_255),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_254),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_273),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_238),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_266),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_259),
.B(n_264),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_281),
.Y(n_286)
);

AOI31xp67_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_257),
.A3(n_259),
.B(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_265),
.B1(n_249),
.B2(n_211),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_283),
.B1(n_267),
.B2(n_270),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_195),
.B1(n_267),
.B2(n_270),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_274),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_283),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_282),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_281),
.B1(n_280),
.B2(n_195),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_284),
.C(n_290),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_288),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_292),
.B(n_286),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_293),
.C(n_291),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_296),
.Y(n_299)
);


endmodule