module fake_jpeg_20922_n_52 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_52);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_26),
.Y(n_30)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_27),
.B1(n_31),
.B2(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.C(n_42),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_21),
.B1(n_4),
.B2(n_8),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_16),
.B(n_9),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_43),
.B(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_17),
.B1(n_12),
.B2(n_13),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_1),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_46),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_20),
.Y(n_52)
);


endmodule