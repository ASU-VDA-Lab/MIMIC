module fake_jpeg_25734_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_19),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_18),
.B1(n_28),
.B2(n_19),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_52),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_20),
.B1(n_28),
.B2(n_21),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_15),
.B1(n_17),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_50),
.B1(n_15),
.B2(n_17),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_24),
.B1(n_22),
.B2(n_26),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_56),
.Y(n_59)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_77),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_35),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_65),
.C(n_67),
.Y(n_87)
);

OAI211xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_37),
.B(n_35),
.C(n_34),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_68),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_36),
.C(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_27),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_73),
.B1(n_76),
.B2(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_17),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_27),
.B1(n_15),
.B2(n_3),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_78),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_30),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_43),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_30),
.B1(n_4),
.B2(n_5),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_54),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_68),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_93),
.C(n_60),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_47),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_56),
.C(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_61),
.B1(n_71),
.B2(n_75),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_89),
.B1(n_97),
.B2(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_99),
.Y(n_104)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_117),
.B1(n_84),
.B2(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_97),
.B1(n_87),
.B2(n_96),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_64),
.C(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_113),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_116),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_70),
.B1(n_74),
.B2(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_128),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_110),
.B1(n_104),
.B2(n_103),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_91),
.B(n_100),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_139),
.B(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_81),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_82),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_138),
.C(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_91),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_90),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_108),
.B(n_107),
.Y(n_153)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_99),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_79),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_140),
.A2(n_110),
.B1(n_92),
.B2(n_101),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_145),
.B1(n_148),
.B2(n_155),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_131),
.B1(n_139),
.B2(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_134),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_108),
.C(n_107),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_130),
.C(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_56),
.B1(n_53),
.B2(n_51),
.Y(n_155)
);

AOI221xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.C(n_7),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_4),
.B(n_5),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_127),
.C(n_132),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_142),
.C(n_148),
.Y(n_160)
);

OAI31xp33_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_124),
.A3(n_134),
.B(n_135),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_161),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_164),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_149),
.C(n_143),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_154),
.C(n_47),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_151),
.B1(n_152),
.B2(n_147),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_152),
.B1(n_154),
.B2(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_175),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_47),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_160),
.C(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_183),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_168),
.B(n_177),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_162),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_159),
.B1(n_45),
.B2(n_7),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_181),
.B1(n_182),
.B2(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_186),
.B(n_6),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_45),
.B1(n_9),
.B2(n_10),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_193),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_189),
.B(n_178),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_180),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_180),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g196 ( 
.A(n_195),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_197),
.B(n_190),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_185),
.B1(n_194),
.B2(n_9),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_11),
.Y(n_200)
);


endmodule