module fake_jpeg_17281_n_374 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_374);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_374;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_43),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_53),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_58),
.Y(n_114)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_20),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_62),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_63),
.B(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_29),
.B(n_1),
.Y(n_64)
);

BUFx12f_ASAP7_75t_SL g65 ( 
.A(n_20),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_37),
.B1(n_29),
.B2(n_20),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_15),
.B(n_1),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_16),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_68),
.A2(n_73),
.B1(n_74),
.B2(n_82),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_76),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_27),
.B1(n_24),
.B2(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_15),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_27),
.B1(n_24),
.B2(n_34),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_78),
.A2(n_88),
.B1(n_90),
.B2(n_94),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_26),
.Y(n_79)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_34),
.B1(n_37),
.B2(n_16),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_15),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_87),
.B(n_95),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_34),
.B1(n_36),
.B2(n_18),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_98),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_55),
.A2(n_23),
.B1(n_33),
.B2(n_32),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_99),
.B1(n_102),
.B2(n_111),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_36),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_38),
.A2(n_33),
.B1(n_32),
.B2(n_28),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_96),
.A2(n_97),
.B1(n_78),
.B2(n_85),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_39),
.A2(n_28),
.B1(n_25),
.B2(n_23),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_25),
.B1(n_21),
.B2(n_19),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_44),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_21),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_19),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_18),
.Y(n_106)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_52),
.A2(n_3),
.B(n_4),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_7),
.B(n_8),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_50),
.A2(n_16),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_65),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_147)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_123),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_71),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

CKINVDCx12_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_138),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_128),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_116),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_140),
.B1(n_152),
.B2(n_154),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_135),
.A2(n_102),
.B(n_96),
.Y(n_194)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_141),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_14),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_144),
.Y(n_170)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_10),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_149),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_72),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_148),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_14),
.B1(n_10),
.B2(n_12),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_81),
.A2(n_10),
.B1(n_14),
.B2(n_109),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_153),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_81),
.A2(n_14),
.B1(n_77),
.B2(n_101),
.Y(n_154)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_158),
.Y(n_205)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_91),
.B(n_117),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_159),
.B(n_114),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_160),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_117),
.B(n_115),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_161),
.B(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_162),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_93),
.A3(n_114),
.B1(n_89),
.B2(n_84),
.Y(n_165)
);

OR2x4_ASAP7_75t_L g166 ( 
.A(n_92),
.B(n_104),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_107),
.B(n_97),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_140),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_95),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_174),
.B(n_208),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_84),
.C(n_85),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_131),
.B1(n_136),
.B2(n_156),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_181),
.A2(n_183),
.B1(n_193),
.B2(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_136),
.A2(n_68),
.B1(n_101),
.B2(n_77),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_189),
.B(n_171),
.Y(n_245)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_98),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_133),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_196),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_146),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_101),
.B1(n_100),
.B2(n_80),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_210),
.B1(n_164),
.B2(n_141),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_113),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_124),
.B(n_130),
.C(n_137),
.Y(n_197)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_120),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_132),
.B(n_100),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_203),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_146),
.A2(n_100),
.B(n_135),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_202),
.A2(n_212),
.B(n_184),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_125),
.B(n_148),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_129),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_145),
.B(n_149),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_186),
.Y(n_230)
);

NAND2x1p5_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_134),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_213),
.A2(n_222),
.B(n_249),
.C(n_219),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_128),
.B1(n_167),
.B2(n_153),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_219),
.B1(n_231),
.B2(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_218),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_121),
.B1(n_153),
.B2(n_163),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_212),
.A2(n_121),
.B1(n_163),
.B2(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_185),
.Y(n_224)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_232),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_191),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_181),
.A2(n_190),
.B1(n_169),
.B2(n_192),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_233),
.A2(n_241),
.B1(n_246),
.B2(n_187),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_170),
.B(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_204),
.B1(n_172),
.B2(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_176),
.B(n_183),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_187),
.Y(n_265)
);

BUFx2_ASAP7_75t_SL g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_188),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_188),
.A2(n_172),
.B1(n_195),
.B2(n_202),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_188),
.A2(n_171),
.B1(n_178),
.B2(n_182),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_180),
.B1(n_179),
.B2(n_211),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_207),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_182),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_249),
.B(n_211),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_175),
.A2(n_184),
.B1(n_207),
.B2(n_200),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_179),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_175),
.B(n_180),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_198),
.C(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_254),
.B(n_280),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_255),
.A2(n_273),
.B(n_275),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_267),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_262),
.B(n_265),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_268),
.B1(n_276),
.B2(n_279),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_235),
.A2(n_198),
.B1(n_237),
.B2(n_226),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_277),
.C(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_214),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_227),
.B(n_223),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_223),
.A2(n_215),
.B1(n_227),
.B2(n_241),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_214),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_245),
.C(n_215),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_213),
.A2(n_233),
.B1(n_225),
.B2(n_231),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_281),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_242),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_221),
.C(n_234),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_286),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_262),
.A2(n_258),
.B(n_251),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_284),
.B(n_285),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_266),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_261),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_300),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_221),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_297),
.C(n_299),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_217),
.Y(n_295)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_221),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_258),
.A2(n_251),
.A3(n_271),
.B1(n_225),
.B2(n_279),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_309),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_256),
.Y(n_300)
);

OA22x2_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_216),
.B1(n_230),
.B2(n_246),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_273),
.B1(n_272),
.B2(n_252),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_220),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_273),
.B1(n_264),
.B2(n_252),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_269),
.B1(n_293),
.B2(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_255),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_307),
.Y(n_321)
);

A2O1A1O1Ixp25_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_221),
.B(n_236),
.C(n_275),
.D(n_276),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_269),
.B(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_313),
.A2(n_314),
.B1(n_318),
.B2(n_320),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_270),
.B1(n_277),
.B2(n_259),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_315),
.A2(n_327),
.B(n_325),
.C(n_310),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_324),
.B1(n_309),
.B2(n_291),
.Y(n_330)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_308),
.B1(n_292),
.B2(n_288),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_293),
.A2(n_304),
.B1(n_288),
.B2(n_305),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_323),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_301),
.A2(n_298),
.B1(n_295),
.B2(n_299),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_303),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_306),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_297),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_291),
.C(n_287),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_330),
.A2(n_332),
.B1(n_336),
.B2(n_337),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_302),
.C(n_287),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_331),
.B(n_341),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_334),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_329),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_324),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_335),
.A2(n_316),
.B1(n_343),
.B2(n_292),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_321),
.A2(n_312),
.B1(n_313),
.B2(n_320),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_336),
.A2(n_335),
.B1(n_318),
.B2(n_313),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_322),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_322),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_340),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_326),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_323),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_343),
.B(n_330),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_344),
.A2(n_329),
.B(n_315),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_345),
.Y(n_357)
);

NAND4xp25_ASAP7_75t_SL g348 ( 
.A(n_335),
.B(n_342),
.C(n_341),
.D(n_339),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_348),
.B(n_351),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_355),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_333),
.C(n_338),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_349),
.C(n_350),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_355),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_358),
.C(n_359),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_340),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_361),
.B(n_354),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_356),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_364),
.Y(n_368)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_360),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_SL g367 ( 
.A1(n_365),
.A2(n_348),
.B(n_346),
.C(n_352),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_359),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_366),
.B(n_367),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_363),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_369),
.A2(n_367),
.B(n_360),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_371),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_370),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_361),
.Y(n_374)
);


endmodule