module real_jpeg_16654_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_572;
wire n_412;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_1),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_1),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_2),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_2),
.A2(n_65),
.B1(n_155),
.B2(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_2),
.A2(n_155),
.B1(n_381),
.B2(n_495),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_2),
.A2(n_155),
.B1(n_504),
.B2(n_506),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_34),
.B1(n_65),
.B2(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_3),
.A2(n_68),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_3),
.A2(n_68),
.B1(n_249),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_3),
.A2(n_68),
.B1(n_433),
.B2(n_438),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_4),
.A2(n_177),
.B1(n_179),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_4),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_4),
.A2(n_181),
.B1(n_381),
.B2(n_383),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_5),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_5),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_6),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_6),
.A2(n_33),
.B1(n_249),
.B2(n_253),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_6),
.A2(n_33),
.B1(n_410),
.B2(n_413),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_6),
.A2(n_33),
.B1(n_482),
.B2(n_485),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_7),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_7),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_7),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_8),
.B(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_8),
.A2(n_84),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_8),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_8),
.A2(n_418),
.A3(n_421),
.B1(n_424),
.B2(n_429),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_8),
.B(n_69),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_8),
.A2(n_97),
.B1(n_520),
.B2(n_526),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_8),
.A2(n_327),
.B1(n_545),
.B2(n_549),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_9),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_9),
.A2(n_150),
.B1(n_303),
.B2(n_309),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_9),
.A2(n_150),
.B1(n_473),
.B2(n_477),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_9),
.A2(n_150),
.B1(n_521),
.B2(n_523),
.Y(n_520)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_104),
.B1(n_110),
.B2(n_111),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_10),
.A2(n_110),
.B1(n_220),
.B2(n_224),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_10),
.A2(n_110),
.B1(n_352),
.B2(n_356),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_10),
.A2(n_110),
.B1(n_580),
.B2(n_581),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_11),
.A2(n_120),
.B1(n_125),
.B2(n_129),
.Y(n_119)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_11),
.A2(n_129),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

AOI22x1_ASAP7_75t_SL g371 ( 
.A1(n_11),
.A2(n_129),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_12),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_13),
.A2(n_162),
.B1(n_167),
.B2(n_170),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_13),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_13),
.A2(n_170),
.B1(n_286),
.B2(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_13),
.A2(n_93),
.B1(n_170),
.B2(n_586),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_14),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_15),
.Y(n_109)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_15),
.Y(n_114)
);

BUFx4f_ASAP7_75t_L g321 ( 
.A(n_15),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_16),
.A2(n_232),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_16),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_16),
.A2(n_236),
.B1(n_258),
.B2(n_262),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_16),
.A2(n_236),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_16),
.A2(n_148),
.B1(n_236),
.B2(n_393),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_17),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_17),
.Y(n_154)
);

BUFx8_ASAP7_75t_L g582 ( 
.A(n_17),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_568),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_398),
.B(n_563),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_328),
.C(n_362),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_264),
.B(n_293),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_24),
.B(n_264),
.C(n_565),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_157),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_25),
.B(n_158),
.C(n_227),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_71),
.C(n_130),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_26),
.A2(n_130),
.B1(n_131),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_26),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_38),
.B1(n_64),
.B2(n_69),
.Y(n_26)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_27),
.Y(n_276)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_31),
.Y(n_275)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_31),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_32),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_32),
.Y(n_377)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g255 ( 
.A(n_38),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_38),
.A2(n_69),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_47),
.B(n_52),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_45),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_47),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_57),
.Y(n_287)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_60),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_60),
.Y(n_239)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_60),
.Y(n_291)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_60),
.Y(n_428)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_64),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_67),
.Y(n_588)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22x1_ASAP7_75t_L g254 ( 
.A1(n_70),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_70),
.A2(n_255),
.B1(n_272),
.B2(n_276),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_70),
.A2(n_255),
.B1(n_272),
.B2(n_302),
.Y(n_301)
);

OAI22x1_ASAP7_75t_SL g350 ( 
.A1(n_70),
.A2(n_255),
.B1(n_257),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_70),
.A2(n_255),
.B1(n_302),
.B2(n_544),
.Y(n_543)
);

OAI22x1_ASAP7_75t_SL g584 ( 
.A1(n_70),
.A2(n_255),
.B1(n_371),
.B2(n_585),
.Y(n_584)
);

XOR2x1_ASAP7_75t_L g265 ( 
.A(n_71),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_96),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_72),
.B(n_96),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_83),
.B1(n_87),
.B2(n_92),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_85),
.Y(n_282)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_85),
.Y(n_349)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AO21x2_ASAP7_75t_L g132 ( 
.A1(n_87),
.A2(n_133),
.B(n_141),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_89),
.Y(n_394)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_102),
.B1(n_115),
.B2(n_119),
.Y(n_96)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_97),
.A2(n_119),
.B1(n_161),
.B2(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_97),
.A2(n_173),
.B(n_176),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_97),
.A2(n_481),
.B1(n_488),
.B2(n_489),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_97),
.A2(n_115),
.B1(n_503),
.B2(n_520),
.Y(n_531)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_99),
.Y(n_325)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_101),
.Y(n_466)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_101),
.Y(n_522)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_103),
.A2(n_171),
.B1(n_314),
.B2(n_322),
.Y(n_313)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_109),
.Y(n_437)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_118),
.Y(n_488)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_124),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_146),
.B1(n_151),
.B2(n_152),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_132),
.A2(n_151),
.B1(n_152),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_132),
.A2(n_146),
.B1(n_151),
.B2(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_132),
.A2(n_151),
.B1(n_248),
.B2(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_132),
.A2(n_151),
.B1(n_348),
.B2(n_392),
.Y(n_391)
);

OAI22x1_ASAP7_75t_SL g578 ( 
.A1(n_132),
.A2(n_151),
.B1(n_392),
.B2(n_579),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_140),
.Y(n_252)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_144),
.Y(n_261)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_144),
.Y(n_420)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2x1_ASAP7_75t_R g326 ( 
.A(n_151),
.B(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_SL g253 ( 
.A(n_153),
.Y(n_253)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_156),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_227),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_182),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_159),
.A2(n_183),
.B(n_205),
.Y(n_345)
);

AOI22x1_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_165),
.Y(n_317)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_166),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_171),
.A2(n_314),
.B1(n_432),
.B2(n_440),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_171),
.A2(n_502),
.B1(n_509),
.B2(n_510),
.Y(n_501)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_205),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_195),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_206),
.B1(n_219),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_184),
.A2(n_206),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_184),
.A2(n_206),
.B1(n_469),
.B2(n_472),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_184),
.A2(n_206),
.B1(n_472),
.B2(n_494),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_184),
.A2(n_206),
.B1(n_409),
.B2(n_494),
.Y(n_553)
);

OA21x2_ASAP7_75t_L g589 ( 
.A1(n_184),
.A2(n_206),
.B(n_380),
.Y(n_589)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_185),
.A2(n_284),
.B1(n_285),
.B2(n_292),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_185),
.A2(n_196),
.B1(n_284),
.B2(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_185),
.A2(n_284),
.B1(n_285),
.B2(n_408),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_185),
.B(n_327),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_191),
.Y(n_487)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_204),
.Y(n_414)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_204),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_219),
.Y(n_205)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_206),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_212),
.B1(n_216),
.B2(n_218),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_210),
.Y(n_423)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_211),
.Y(n_457)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g461 ( 
.A(n_215),
.Y(n_461)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_217),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_226),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_226),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_226),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_246),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_228),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_240),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_229),
.A2(n_230),
.B1(n_240),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_235),
.Y(n_384)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_239),
.Y(n_471)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_244),
.Y(n_529)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_245),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_247),
.B(n_254),
.C(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx2_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_265),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_270),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_277),
.C(n_283),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_283),
.Y(n_298)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_291),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_294),
.B(n_296),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_297),
.B(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_299),
.B(n_300),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_312),
.C(n_326),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_301),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_308),
.Y(n_355)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_312),
.A2(n_313),
.B1(n_326),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_317),
.Y(n_439)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_321),
.Y(n_505)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_321),
.Y(n_508)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_321),
.Y(n_525)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_323),
.B(n_327),
.Y(n_518)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_327),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_327),
.B(n_455),
.Y(n_454)
);

OAI21xp33_ASAP7_75t_SL g469 ( 
.A1(n_327),
.A2(n_454),
.B(n_470),
.Y(n_469)
);

A2O1A1O1Ixp25_ASAP7_75t_L g563 ( 
.A1(n_328),
.A2(n_362),
.B(n_564),
.C(n_566),
.D(n_567),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_361),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_SL g566 ( 
.A(n_329),
.B(n_361),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_344),
.B1(n_359),
.B2(n_360),
.Y(n_332)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_360),
.C(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g343 ( 
.A(n_334),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_334),
.B(n_342),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_341),
.A2(n_342),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_341),
.A2(n_391),
.B(n_395),
.Y(n_574)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_344),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_350),
.C(n_365),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_351),
.Y(n_369)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_355),
.Y(n_358)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_396),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_363),
.B(n_396),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_364),
.B(n_571),
.C(n_572),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_386),
.Y(n_366)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_367),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_378),
.B(n_385),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_378),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_377),
.Y(n_551)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_385),
.A2(n_576),
.B1(n_591),
.B2(n_592),
.Y(n_575)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_385),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_386),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_388),
.B1(n_389),
.B2(n_395),
.Y(n_386)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_387),
.Y(n_395)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_443),
.B(n_562),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_400),
.B(n_402),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_407),
.C(n_415),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_403),
.A2(n_404),
.B1(n_558),
.B2(n_559),
.Y(n_557)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_407),
.A2(n_415),
.B1(n_416),
.B2(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_407),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_430),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_417),
.A2(n_430),
.B1(n_431),
.B2(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_417),
.Y(n_540)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_432),
.Y(n_489)
);

OAI32xp33_ASAP7_75t_L g448 ( 
.A1(n_433),
.A2(n_449),
.A3(n_451),
.B1(n_454),
.B2(n_458),
.Y(n_448)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx6_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx6_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_555),
.B(n_561),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_536),
.B(n_554),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_499),
.B(n_535),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_479),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_447),
.B(n_479),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_467),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_448),
.A2(n_467),
.B1(n_468),
.B2(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_448),
.Y(n_512)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_490),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_492),
.C(n_498),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_481),
.Y(n_510)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_492),
.B1(n_493),
.B2(n_498),
.Y(n_490)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_491),
.Y(n_498)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_513),
.B(n_534),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_511),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_501),
.B(n_511),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_514),
.A2(n_530),
.B(n_533),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_519),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_518),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx4_ASAP7_75t_SL g528 ( 
.A(n_529),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_532),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_538),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_537),
.B(n_538),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_541),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_539),
.B(n_542),
.C(n_553),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_542),
.A2(n_543),
.B1(n_552),
.B2(n_553),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_557),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_556),
.B(n_557),
.Y(n_561)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g568 ( 
.A(n_569),
.B(n_593),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_573),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_570),
.B(n_573),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_574),
.B(n_575),
.Y(n_573)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_576),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_577),
.A2(n_578),
.B1(n_583),
.B2(n_590),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

BUFx12f_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_583),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_589),
.Y(n_583)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);


endmodule