module real_jpeg_33158_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g142 ( 
.A(n_0),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_0),
.Y(n_330)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_0),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_1),
.A2(n_86),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_1),
.A2(n_90),
.B1(n_222),
.B2(n_225),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_1),
.A2(n_90),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_97),
.B1(n_98),
.B2(n_103),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_2),
.A2(n_97),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_2),
.A2(n_97),
.B1(n_225),
.B2(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_2),
.A2(n_97),
.B1(n_215),
.B2(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_3),
.B(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_3),
.A2(n_135),
.B(n_231),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_3),
.A2(n_113),
.A3(n_302),
.B1(n_307),
.B2(n_310),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_3),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_3),
.A2(n_311),
.B1(n_367),
.B2(n_372),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_3),
.B(n_73),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_3),
.A2(n_141),
.B1(n_450),
.B2(n_464),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_4),
.A2(n_162),
.B1(n_163),
.B2(n_166),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_4),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_4),
.A2(n_162),
.B1(n_183),
.B2(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_5),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_7),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_7),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_8),
.A2(n_203),
.B1(n_206),
.B2(n_210),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

AO22x1_ASAP7_75t_L g278 ( 
.A1(n_8),
.A2(n_210),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_8),
.A2(n_210),
.B1(n_332),
.B2(n_336),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_42),
.B1(n_46),
.B2(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_9),
.A2(n_50),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_9),
.A2(n_50),
.B1(n_186),
.B2(n_377),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_9),
.A2(n_50),
.B1(n_438),
.B2(n_441),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_10),
.Y(n_185)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_10),
.Y(n_195)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_12),
.A2(n_42),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_12),
.A2(n_64),
.B1(n_345),
.B2(n_348),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_12),
.A2(n_64),
.B1(n_404),
.B2(n_409),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_12),
.A2(n_64),
.B1(n_451),
.B2(n_453),
.Y(n_450)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_13),
.Y(n_177)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_15),
.A2(n_148),
.B1(n_149),
.B2(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_15),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_15),
.A2(n_148),
.B1(n_183),
.B2(n_186),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_16),
.A2(n_163),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_16),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_17),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_17),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_287),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_247),
.B(n_285),
.Y(n_19)
);

HB1xp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_22),
.B(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_169),
.C(n_217),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_24),
.B(n_495),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_117),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_70),
.B2(n_71),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_27),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_40),
.B1(n_51),
.B2(n_62),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_29),
.A2(n_63),
.B1(n_230),
.B2(n_234),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_29),
.A2(n_41),
.B1(n_234),
.B2(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_29),
.B(n_311),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_32),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_32),
.Y(n_371)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_45),
.Y(n_272)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_51),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_58),
.B2(n_60),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_58),
.Y(n_233)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_70),
.B(n_251),
.C(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_85),
.B1(n_96),
.B2(n_106),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g343 ( 
.A1(n_72),
.A2(n_106),
.B1(n_237),
.B2(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_72),
.A2(n_106),
.B1(n_344),
.B2(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_73),
.A2(n_236),
.B1(n_245),
.B2(n_246),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_73),
.A2(n_245),
.B1(n_278),
.B2(n_284),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AO21x2_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_107),
.B(n_113),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_80),
.B2(n_82),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_76),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_76),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_76),
.Y(n_209)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_81),
.Y(n_309)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_85),
.Y(n_284)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_89),
.Y(n_347)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_94),
.Y(n_280)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_96),
.Y(n_246)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_101),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_102),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_102),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_102),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g245 ( 
.A(n_106),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_138),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_118),
.B(n_138),
.Y(n_251)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.A3(n_124),
.B1(n_128),
.B2(n_134),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g484 ( 
.A1(n_119),
.A2(n_121),
.A3(n_124),
.B1(n_128),
.B2(n_134),
.Y(n_484)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_138),
.A2(n_139),
.B1(n_484),
.B2(n_485),
.Y(n_483)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_147),
.B1(n_157),
.B2(n_160),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_140),
.A2(n_319),
.B1(n_327),
.B2(n_331),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_140),
.A2(n_147),
.B1(n_331),
.B2(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_140),
.A2(n_436),
.B1(n_442),
.B2(n_443),
.Y(n_435)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_141),
.A2(n_161),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_141),
.A2(n_213),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_141),
.A2(n_418),
.B1(n_424),
.B2(n_427),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_141),
.A2(n_437),
.B1(n_450),
.B2(n_457),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_175),
.B1(n_178),
.B2(n_180),
.Y(n_174)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_146),
.Y(n_335)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_155),
.Y(n_452)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_156),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_156),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_157),
.Y(n_212)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_159),
.Y(n_261)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_166),
.Y(n_441)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx2_ASAP7_75t_SL g337 ( 
.A(n_167),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_168),
.Y(n_393)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_168),
.Y(n_456)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_170),
.B(n_218),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_211),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_171),
.B(n_211),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_182),
.B1(n_189),
.B2(n_202),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_172),
.A2(n_189),
.B1(n_202),
.B2(n_221),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_172),
.A2(n_182),
.B1(n_189),
.B2(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_172),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_172),
.A2(n_189),
.B1(n_376),
.B2(n_402),
.Y(n_430)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AO21x2_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_190),
.B(n_196),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_176),
.Y(n_395)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_185),
.Y(n_408)
);

BUFx6f_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_189),
.A2(n_221),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_189),
.Y(n_381)
);

NAND2xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_195),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_196),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_209),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_228),
.C(n_235),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_219),
.A2(n_220),
.B1(n_228),
.B2(n_229),
.Y(n_488)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_235),
.B(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_277),
.Y(n_268)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_491),
.B(n_496),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_480),
.B(n_490),
.Y(n_289)
);

OAI21x1_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_382),
.B(n_479),
.Y(n_290)
);

AOI211xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_340),
.B(n_360),
.C(n_361),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_292),
.A2(n_340),
.B(n_360),
.C(n_361),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_293),
.B(n_342),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_300),
.B1(n_338),
.B2(n_339),
.Y(n_293)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_294),
.B(n_338),
.C(n_341),
.Y(n_489)
);

OAI22x1_ASAP7_75t_L g401 ( 
.A1(n_295),
.A2(n_402),
.B1(n_410),
.B2(n_411),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_295),
.B(n_311),
.Y(n_461)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_296),
.A2(n_298),
.B1(n_375),
.B2(n_381),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_317),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_301),
.A2(n_317),
.B1(n_318),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_301),
.Y(n_363)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_311),
.B(n_397),
.Y(n_396)
);

OA21x2_ASAP7_75t_SL g411 ( 
.A1(n_311),
.A2(n_396),
.B(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_311),
.B(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_316),
.Y(n_380)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_319),
.Y(n_427)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_325),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_330),
.Y(n_445)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_351),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_343),
.B(n_352),
.C(n_359),
.Y(n_486)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_358),
.B2(n_359),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_356),
.Y(n_468)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_357),
.Y(n_460)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.C(n_374),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_362),
.B(n_476),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_364),
.A2(n_365),
.B1(n_374),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_381),
.Y(n_410)
);

AOI21x1_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_473),
.B(n_478),
.Y(n_382)
);

OAI21x1_ASAP7_75t_SL g383 ( 
.A1(n_384),
.A2(n_433),
.B(n_472),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_416),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_385),
.B(n_416),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_401),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_386),
.B(n_401),
.Y(n_446)
);

AO21x1_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_389),
.B(n_390),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_394),
.B(n_396),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx4f_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_408),
.Y(n_415)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_428),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_417),
.B(n_430),
.C(n_431),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_429),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_430),
.Y(n_432)
);

AOI21x1_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_447),
.B(n_471),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_446),
.Y(n_434)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_446),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_SL g443 ( 
.A(n_444),
.Y(n_443)
);

INVx8_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_462),
.B(n_470),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_461),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_449),
.B(n_461),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_458),
.Y(n_464)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_465),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_SL g478 ( 
.A(n_474),
.B(n_475),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_489),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_489),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_487),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_486),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_487),
.C(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_484),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_486),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_494),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_494),
.Y(n_497)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);


endmodule