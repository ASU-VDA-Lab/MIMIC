module real_jpeg_3231_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_29),
.B1(n_31),
.B2(n_57),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_33),
.B1(n_49),
.B2(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_7),
.B(n_24),
.C(n_38),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_7),
.B(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_7),
.B(n_22),
.C(n_29),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_7),
.B(n_50),
.C(n_60),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_7),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_7),
.B(n_53),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_7),
.B(n_59),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_104),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_103),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_15),
.B(n_90),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_67),
.B1(n_68),
.B2(n_89),
.Y(n_15)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_45),
.B(n_65),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_17),
.A2(n_65),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_34),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_18),
.A2(n_19),
.B1(n_34),
.B2(n_35),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_18),
.A2(n_19),
.B1(n_58),
.B2(n_94),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_18),
.A2(n_19),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_18),
.A2(n_58),
.B(n_114),
.C(n_175),
.Y(n_178)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_19),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_19),
.B(n_94),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_19),
.B(n_102),
.C(n_128),
.Y(n_127)
);

AO21x2_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_28),
.B(n_32),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_21)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

OA22x2_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_42),
.Y(n_43)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_24),
.B(n_143),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_28),
.Y(n_160)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_29),
.A2(n_31),
.B1(n_60),
.B2(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_29),
.B(n_154),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI211xp5_ASAP7_75t_SL g113 ( 
.A1(n_34),
.A2(n_58),
.B(n_66),
.C(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_34),
.A2(n_35),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

AO21x2_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_43),
.B(n_44),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_40),
.B(n_100),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_43),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_45),
.A2(n_70),
.B1(n_71),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_58),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_46),
.A2(n_58),
.B1(n_94),
.B2(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_46),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_50),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_50),
.B(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_73),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_58),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_58),
.B(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_58),
.A2(n_94),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_58),
.A2(n_94),
.B1(n_152),
.B2(n_153),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_58),
.A2(n_94),
.B1(n_140),
.B2(n_181),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_64),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_77),
.B1(n_87),
.B2(n_88),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_76),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_71),
.B1(n_97),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_86),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.C(n_96),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_93),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_136),
.C(n_140),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_94),
.B(n_102),
.C(n_159),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_101),
.A2(n_102),
.B1(n_128),
.B2(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_101),
.A2(n_102),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_101),
.A2(n_102),
.B1(n_141),
.B2(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_102),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_102),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_131),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_117),
.B(n_130),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_132),
.C(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_115),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_112),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_121),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_127),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_123),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_124),
.A2(n_125),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_147),
.B(n_183),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_144),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_177),
.B(n_182),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_171),
.B(n_176),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_161),
.B(n_170),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_155),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_179),
.Y(n_182)
);


endmodule