module fake_netlist_1_3714_n_903 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_903);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_903;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_857;
wire n_786;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_738;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_685;
wire n_362;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_522;
wire n_883;
wire n_573;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_721;
wire n_438;
wire n_656;
wire n_640;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_54), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_46), .Y(n_284) );
INVxp33_ASAP7_75t_L g285 ( .A(n_91), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_253), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_139), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_252), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_32), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_222), .Y(n_291) );
INVxp33_ASAP7_75t_L g292 ( .A(n_52), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_259), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_267), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_244), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_44), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_233), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_2), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_29), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_110), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_265), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_172), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_250), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g305 ( .A(n_256), .B(n_143), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_189), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_11), .Y(n_307) );
BUFx10_ASAP7_75t_L g308 ( .A(n_80), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g309 ( .A(n_166), .B(n_149), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_207), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_17), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_238), .Y(n_312) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_153), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_264), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_257), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_247), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_86), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_165), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_134), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_72), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_212), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_183), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_109), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_218), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_198), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_197), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_269), .B(n_18), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_9), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_211), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_255), .Y(n_330) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_229), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_98), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_60), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_232), .Y(n_334) );
BUFx10_ASAP7_75t_L g335 ( .A(n_245), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_181), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_145), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_276), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_66), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g340 ( .A(n_48), .B(n_159), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_161), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_262), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_71), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_95), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_261), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_278), .Y(n_346) );
INVx1_ASAP7_75t_SL g347 ( .A(n_135), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_186), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_4), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_40), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_10), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_140), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_73), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_129), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_133), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_56), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_11), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_92), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_242), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_105), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_138), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_273), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_147), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_42), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_275), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_270), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_204), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_251), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_179), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_74), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_93), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_228), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_63), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_272), .Y(n_374) );
INVxp67_ASAP7_75t_L g375 ( .A(n_243), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_37), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_13), .Y(n_377) );
CKINVDCx14_ASAP7_75t_R g378 ( .A(n_45), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_239), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_203), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_97), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_122), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_107), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_274), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_171), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_254), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_221), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_14), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_182), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_2), .Y(n_390) );
BUFx5_ASAP7_75t_L g391 ( .A(n_263), .Y(n_391) );
CKINVDCx14_ASAP7_75t_R g392 ( .A(n_156), .Y(n_392) );
CKINVDCx14_ASAP7_75t_R g393 ( .A(n_84), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_191), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_124), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_190), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_67), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_180), .Y(n_398) );
BUFx10_ASAP7_75t_L g399 ( .A(n_258), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_83), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_27), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_141), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_271), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_268), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_28), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_215), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_293), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_291), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_328), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_297), .B(n_0), .Y(n_410) );
OA21x2_ASAP7_75t_L g411 ( .A1(n_288), .A2(n_20), .B(n_19), .Y(n_411) );
OA21x2_ASAP7_75t_L g412 ( .A1(n_289), .A2(n_294), .B(n_290), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_298), .B(n_0), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_391), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_391), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_307), .A2(n_4), .B1(n_1), .B2(n_3), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_296), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_299), .Y(n_418) );
NAND2xp33_ASAP7_75t_L g419 ( .A(n_391), .B(n_21), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_283), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_293), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_315), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_384), .B(n_1), .Y(n_423) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_293), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_311), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_349), .B(n_3), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_322), .B(n_5), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_414), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_408), .B(n_285), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_415), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_422), .B(n_292), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_425), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_417), .B(n_308), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_417), .B(n_378), .Y(n_434) );
INVx4_ASAP7_75t_SL g435 ( .A(n_410), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_426), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_427), .Y(n_437) );
AND2x6_ASAP7_75t_L g438 ( .A(n_410), .B(n_300), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_418), .B(n_295), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_412), .A2(n_388), .B1(n_357), .B2(n_377), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_412), .Y(n_441) );
XOR2xp5_ASAP7_75t_L g442 ( .A(n_420), .B(n_284), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_413), .A2(n_390), .B1(n_393), .B2(n_392), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_423), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_437), .B(n_409), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_444), .A2(n_419), .B1(n_304), .B2(n_312), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_428), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_434), .B(n_286), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_430), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_429), .B(n_303), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_442), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_431), .B(n_310), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_432), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_436), .A2(n_318), .B1(n_337), .B2(n_302), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_438), .A2(n_385), .B1(n_398), .B2(n_395), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_438), .B(n_314), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_441), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_438), .B(n_316), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_435), .B(n_319), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_438), .B(n_321), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_439), .B(n_325), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_433), .B(n_308), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_435), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_443), .B(n_345), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_440), .B(n_301), .Y(n_465) );
INVx4_ASAP7_75t_L g466 ( .A(n_435), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_445), .A2(n_416), .B1(n_351), .B2(n_313), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_466), .B(n_352), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_457), .A2(n_411), .B(n_403), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_453), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_465), .B(n_327), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_448), .A2(n_411), .B(n_405), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_465), .B(n_368), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_464), .A2(n_375), .B(n_317), .C(n_323), .Y(n_474) );
OR2x6_ASAP7_75t_SL g475 ( .A(n_451), .B(n_355), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_454), .B(n_335), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_446), .A2(n_331), .B(n_324), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_456), .A2(n_326), .B(n_320), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_446), .B(n_330), .C(n_329), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_455), .A2(n_332), .B1(n_334), .B2(n_333), .Y(n_480) );
NOR2x1_ASAP7_75t_L g481 ( .A(n_466), .B(n_459), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_450), .B(n_367), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_462), .A2(n_372), .B1(n_386), .B2(n_369), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_458), .A2(n_341), .B(n_336), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_452), .B(n_387), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_460), .A2(n_348), .B(n_342), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g487 ( .A(n_463), .B(n_287), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_461), .A2(n_354), .B1(n_356), .B2(n_350), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_462), .B(n_397), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_447), .A2(n_359), .B(n_360), .C(n_358), .Y(n_490) );
BUFx5_ASAP7_75t_L g491 ( .A(n_476), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_487), .B(n_305), .Y(n_492) );
AO31x2_ASAP7_75t_L g493 ( .A1(n_469), .A2(n_362), .A3(n_363), .B(n_361), .Y(n_493) );
O2A1O1Ixp5_ASAP7_75t_L g494 ( .A1(n_472), .A2(n_339), .B(n_343), .C(n_338), .Y(n_494) );
AOI21x1_ASAP7_75t_L g495 ( .A1(n_471), .A2(n_340), .B(n_309), .Y(n_495) );
NAND2xp33_ASAP7_75t_L g496 ( .A(n_470), .B(n_449), .Y(n_496) );
AO31x2_ASAP7_75t_L g497 ( .A1(n_488), .A2(n_366), .A3(n_370), .B(n_365), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_489), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_479), .A2(n_344), .B1(n_353), .B2(n_347), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_474), .A2(n_373), .B(n_374), .C(n_371), .Y(n_500) );
O2A1O1Ixp5_ASAP7_75t_L g501 ( .A1(n_477), .A2(n_484), .B(n_486), .C(n_478), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_481), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_475), .Y(n_503) );
OAI21x1_ASAP7_75t_L g504 ( .A1(n_473), .A2(n_381), .B(n_380), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_467), .B(n_383), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_482), .A2(n_394), .B(n_389), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_480), .B(n_396), .Y(n_507) );
OAI21x1_ASAP7_75t_L g508 ( .A1(n_468), .A2(n_401), .B(n_400), .Y(n_508) );
AO31x2_ASAP7_75t_L g509 ( .A1(n_485), .A2(n_402), .A3(n_404), .B(n_391), .Y(n_509) );
AO31x2_ASAP7_75t_L g510 ( .A1(n_490), .A2(n_391), .A3(n_421), .B(n_407), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_479), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_483), .A2(n_382), .B1(n_406), .B2(n_346), .Y(n_512) );
NOR2xp67_ASAP7_75t_SL g513 ( .A(n_476), .B(n_379), .Y(n_513) );
AO32x2_ASAP7_75t_L g514 ( .A1(n_480), .A2(n_424), .A3(n_421), .B1(n_407), .B2(n_399), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_469), .A2(n_364), .B(n_306), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_476), .B(n_335), .Y(n_516) );
AO31x2_ASAP7_75t_L g517 ( .A1(n_469), .A2(n_421), .A3(n_424), .B(n_407), .Y(n_517) );
OAI21x1_ASAP7_75t_L g518 ( .A1(n_469), .A2(n_364), .B(n_306), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_470), .Y(n_519) );
AOI221x1_ASAP7_75t_L g520 ( .A1(n_469), .A2(n_424), .B1(n_376), .B2(n_364), .C(n_306), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_519), .Y(n_521) );
BUFx3_ASAP7_75t_L g522 ( .A(n_503), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_493), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_501), .A2(n_399), .B(n_5), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_498), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_491), .A2(n_376), .B1(n_8), .B2(n_6), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_491), .B(n_6), .Y(n_527) );
OAI21x1_ASAP7_75t_L g528 ( .A1(n_518), .A2(n_376), .B(n_23), .Y(n_528) );
BUFx2_ASAP7_75t_SL g529 ( .A(n_491), .Y(n_529) );
INVx4_ASAP7_75t_L g530 ( .A(n_492), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_497), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_506), .A2(n_9), .B(n_7), .C(n_8), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_505), .B(n_7), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_515), .A2(n_24), .B(n_22), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_494), .A2(n_26), .B(n_25), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_516), .B(n_10), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_496), .A2(n_31), .B(n_30), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_507), .B(n_12), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_504), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_520), .A2(n_34), .B(n_33), .Y(n_540) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_495), .A2(n_36), .B(n_35), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_511), .A2(n_39), .B(n_38), .Y(n_542) );
AO31x2_ASAP7_75t_L g543 ( .A1(n_500), .A2(n_14), .A3(n_12), .B(n_13), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_508), .Y(n_544) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_517), .A2(n_502), .B(n_510), .Y(n_545) );
BUFx12f_ASAP7_75t_L g546 ( .A(n_513), .Y(n_546) );
AO31x2_ASAP7_75t_L g547 ( .A1(n_517), .A2(n_43), .A3(n_47), .B(n_41), .Y(n_547) );
NOR2x1_ASAP7_75t_SL g548 ( .A(n_512), .B(n_15), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_499), .A2(n_17), .B(n_15), .C(n_16), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_497), .B(n_16), .Y(n_550) );
INVx6_ASAP7_75t_L g551 ( .A(n_514), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_510), .Y(n_552) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_509), .A2(n_50), .B(n_49), .Y(n_553) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_509), .A2(n_53), .B(n_51), .Y(n_554) );
INVx6_ASAP7_75t_L g555 ( .A(n_514), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_519), .Y(n_556) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_518), .A2(n_57), .B(n_55), .Y(n_557) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_519), .Y(n_558) );
BUFx2_ASAP7_75t_L g559 ( .A(n_519), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_491), .B(n_18), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_501), .A2(n_58), .B(n_59), .Y(n_561) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_518), .A2(n_61), .B(n_62), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_491), .B(n_64), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_515), .A2(n_65), .B(n_68), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_556), .B(n_69), .Y(n_565) );
OA21x2_ASAP7_75t_L g566 ( .A1(n_524), .A2(n_70), .B(n_75), .Y(n_566) );
BUFx2_ASAP7_75t_L g567 ( .A(n_546), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_544), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_558), .Y(n_569) );
OA21x2_ASAP7_75t_L g570 ( .A1(n_552), .A2(n_76), .B(n_77), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_556), .B(n_78), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_559), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_539), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_529), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_525), .B(n_79), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_558), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_545), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_550), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_522), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_531), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_545), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_538), .Y(n_583) );
OA21x2_ASAP7_75t_L g584 ( .A1(n_561), .A2(n_81), .B(n_82), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_543), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_548), .B(n_85), .Y(n_586) );
BUFx4f_ASAP7_75t_SL g587 ( .A(n_530), .Y(n_587) );
NOR2xp33_ASAP7_75t_SL g588 ( .A(n_527), .B(n_87), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_536), .B(n_88), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_551), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_523), .B(n_89), .Y(n_591) );
AO21x2_ASAP7_75t_L g592 ( .A1(n_540), .A2(n_90), .B(n_94), .Y(n_592) );
AO21x2_ASAP7_75t_L g593 ( .A1(n_528), .A2(n_96), .B(n_99), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_543), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_543), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_560), .Y(n_596) );
INVx2_ASAP7_75t_SL g597 ( .A(n_563), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_533), .B(n_100), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_532), .B(n_101), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_551), .Y(n_600) );
BUFx2_ASAP7_75t_L g601 ( .A(n_555), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_555), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_549), .B(n_526), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_541), .B(n_102), .Y(n_604) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_557), .A2(n_103), .B(n_104), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_547), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_547), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_553), .B(n_106), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_553), .B(n_108), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_554), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_562), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_554), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_564), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_535), .Y(n_614) );
AND2x4_ASAP7_75t_SL g615 ( .A(n_537), .B(n_542), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_534), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_558), .Y(n_617) );
BUFx12f_ASAP7_75t_L g618 ( .A(n_546), .Y(n_618) );
AO22x1_ASAP7_75t_L g619 ( .A1(n_527), .A2(n_111), .B1(n_112), .B2(n_113), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_556), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_544), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_544), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_556), .B(n_114), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_521), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_556), .B(n_115), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_544), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_556), .B(n_116), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_521), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_556), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_556), .B(n_117), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_544), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_521), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_556), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_556), .B(n_118), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_544), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_578), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_628), .B(n_119), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_620), .B(n_120), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_620), .B(n_121), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_629), .B(n_123), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_629), .B(n_125), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_569), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_633), .B(n_126), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_578), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_624), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_633), .B(n_127), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_583), .B(n_128), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_632), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_572), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_581), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_573), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_582), .Y(n_652) );
BUFx3_ASAP7_75t_L g653 ( .A(n_569), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_582), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_573), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_577), .B(n_130), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_574), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_577), .B(n_131), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_623), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_574), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_568), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_623), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_575), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_575), .B(n_282), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_568), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_621), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_617), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_565), .A2(n_132), .B1(n_136), .B2(n_137), .Y(n_668) );
INVx3_ASAP7_75t_L g669 ( .A(n_617), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_579), .B(n_142), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_596), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_603), .A2(n_144), .B1(n_146), .B2(n_148), .C(n_150), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_585), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_594), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_621), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_576), .B(n_151), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_595), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_580), .B(n_281), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_571), .B(n_152), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_625), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_627), .B(n_154), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_597), .B(n_155), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_630), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_634), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_586), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_590), .Y(n_686) );
BUFx2_ASAP7_75t_L g687 ( .A(n_587), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_622), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g689 ( .A(n_587), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_598), .B(n_157), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_590), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_622), .Y(n_692) );
INVx4_ASAP7_75t_L g693 ( .A(n_618), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_602), .B(n_158), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_626), .Y(n_695) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_626), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_607), .B(n_160), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_600), .Y(n_698) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_631), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_589), .B(n_162), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_599), .B(n_567), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_601), .B(n_280), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_631), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_600), .B(n_163), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_635), .B(n_279), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_635), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_588), .B(n_164), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_588), .B(n_606), .Y(n_708) );
BUFx3_ASAP7_75t_L g709 ( .A(n_591), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_608), .B(n_167), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_591), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_611), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_616), .B(n_604), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_619), .B(n_168), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_611), .Y(n_715) );
INVx2_ASAP7_75t_SL g716 ( .A(n_570), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_593), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_605), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_593), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_570), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_566), .A2(n_169), .B1(n_170), .B2(n_173), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_566), .Y(n_722) );
BUFx3_ASAP7_75t_L g723 ( .A(n_615), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_609), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_613), .B(n_174), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_655), .B(n_612), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_663), .B(n_616), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_671), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_645), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_648), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_650), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_680), .B(n_610), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_649), .Y(n_733) );
INVxp67_ASAP7_75t_L g734 ( .A(n_655), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_683), .B(n_610), .Y(n_735) );
AND2x2_ASAP7_75t_SL g736 ( .A(n_659), .B(n_584), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_636), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_684), .B(n_592), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_651), .B(n_592), .Y(n_739) );
AND2x4_ASAP7_75t_L g740 ( .A(n_659), .B(n_615), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_686), .B(n_614), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_674), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_711), .B(n_614), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_685), .B(n_584), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_691), .B(n_175), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_701), .B(n_176), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_698), .B(n_177), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_713), .B(n_178), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_677), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_636), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_667), .B(n_184), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_665), .B(n_185), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_713), .B(n_187), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_673), .B(n_709), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_666), .B(n_188), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_662), .B(n_192), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_673), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_675), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_639), .B(n_193), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_640), .B(n_194), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_688), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_644), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_641), .B(n_195), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_692), .Y(n_764) );
INVx4_ASAP7_75t_L g765 ( .A(n_687), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_652), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_643), .B(n_196), .Y(n_767) );
INVx3_ASAP7_75t_L g768 ( .A(n_723), .Y(n_768) );
INVx3_ASAP7_75t_L g769 ( .A(n_723), .Y(n_769) );
INVx2_ASAP7_75t_SL g770 ( .A(n_689), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_646), .B(n_199), .Y(n_771) );
OR2x2_ASAP7_75t_L g772 ( .A(n_654), .B(n_200), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_709), .A2(n_201), .B1(n_202), .B2(n_205), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_654), .B(n_206), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_696), .B(n_208), .Y(n_775) );
BUFx2_ASAP7_75t_L g776 ( .A(n_642), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_657), .Y(n_777) );
OR2x2_ASAP7_75t_L g778 ( .A(n_696), .B(n_209), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_657), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_653), .B(n_210), .Y(n_780) );
NOR2xp67_ASAP7_75t_L g781 ( .A(n_714), .B(n_213), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_669), .B(n_214), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_660), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_669), .B(n_216), .Y(n_784) );
OR2x2_ASAP7_75t_L g785 ( .A(n_699), .B(n_217), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_660), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_647), .B(n_219), .Y(n_787) );
BUFx3_ASAP7_75t_L g788 ( .A(n_689), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_638), .B(n_220), .Y(n_789) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_699), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_661), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_734), .B(n_661), .Y(n_792) );
NOR2x1_ASAP7_75t_L g793 ( .A(n_765), .B(n_693), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_731), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_765), .B(n_693), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_728), .B(n_724), .Y(n_796) );
NAND2xp33_ASAP7_75t_L g797 ( .A(n_768), .B(n_668), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_740), .A2(n_672), .B1(n_708), .B2(n_668), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_781), .A2(n_672), .B1(n_707), .B2(n_681), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_733), .B(n_695), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_770), .B(n_678), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_729), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_737), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_737), .B(n_695), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_730), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_742), .B(n_703), .Y(n_806) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_776), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_727), .B(n_703), .Y(n_808) );
OR2x2_ASAP7_75t_L g809 ( .A(n_790), .B(n_706), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_749), .B(n_757), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_732), .B(n_706), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_735), .B(n_704), .Y(n_812) );
AND2x4_ASAP7_75t_L g813 ( .A(n_740), .B(n_712), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_758), .B(n_697), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_761), .B(n_697), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_726), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_788), .B(n_664), .Y(n_817) );
NAND4xp25_ASAP7_75t_L g818 ( .A(n_781), .B(n_721), .C(n_670), .D(n_682), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_790), .Y(n_819) );
INVx2_ASAP7_75t_SL g820 ( .A(n_788), .Y(n_820) );
NOR2x1_ASAP7_75t_L g821 ( .A(n_768), .B(n_702), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_754), .B(n_712), .Y(n_822) );
AND2x2_ASAP7_75t_SL g823 ( .A(n_769), .B(n_679), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_754), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_764), .B(n_725), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_769), .B(n_710), .Y(n_826) );
NAND2x1_ASAP7_75t_L g827 ( .A(n_766), .B(n_718), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_744), .B(n_717), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_777), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g830 ( .A(n_736), .B(n_694), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_791), .B(n_670), .Y(n_831) );
AOI32xp33_ASAP7_75t_L g832 ( .A1(n_793), .A2(n_746), .A3(n_789), .B1(n_760), .B2(n_759), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_810), .Y(n_833) );
AND2x4_ASAP7_75t_L g834 ( .A(n_807), .B(n_738), .Y(n_834) );
INVx2_ASAP7_75t_SL g835 ( .A(n_820), .Y(n_835) );
AND3x2_ASAP7_75t_L g836 ( .A(n_795), .B(n_780), .C(n_767), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_794), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g838 ( .A(n_823), .B(n_736), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_797), .A2(n_748), .B1(n_753), .B2(n_739), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_824), .B(n_743), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_816), .B(n_743), .Y(n_841) );
OR2x2_ASAP7_75t_L g842 ( .A(n_819), .B(n_750), .Y(n_842) );
OR2x2_ASAP7_75t_L g843 ( .A(n_822), .B(n_762), .Y(n_843) );
INVxp67_ASAP7_75t_L g844 ( .A(n_801), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_811), .B(n_741), .Y(n_845) );
NOR2xp67_ASAP7_75t_L g846 ( .A(n_799), .B(n_721), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_808), .B(n_741), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_802), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_812), .B(n_779), .Y(n_849) );
NOR2x1_ASAP7_75t_L g850 ( .A(n_821), .B(n_775), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_813), .B(n_783), .Y(n_851) );
A2O1A1Ixp33_ASAP7_75t_L g852 ( .A1(n_799), .A2(n_787), .B(n_748), .C(n_753), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_809), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g854 ( .A1(n_833), .A2(n_805), .B1(n_796), .B2(n_830), .C(n_817), .Y(n_854) );
AOI32xp33_ASAP7_75t_L g855 ( .A1(n_838), .A2(n_798), .A3(n_826), .B1(n_813), .B2(n_763), .Y(n_855) );
OAI21xp5_ASAP7_75t_SL g856 ( .A1(n_836), .A2(n_818), .B(n_773), .Y(n_856) );
NOR3xp33_ASAP7_75t_L g857 ( .A(n_852), .B(n_818), .C(n_745), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_837), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_849), .B(n_803), .Y(n_859) );
NAND2xp5_ASAP7_75t_SL g860 ( .A(n_832), .B(n_846), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_848), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_834), .B(n_828), .Y(n_862) );
O2A1O1Ixp33_ASAP7_75t_L g863 ( .A1(n_844), .A2(n_814), .B(n_815), .C(n_831), .Y(n_863) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_841), .A2(n_825), .B1(n_829), .B2(n_806), .C(n_800), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_840), .B(n_792), .Y(n_865) );
AOI21xp33_ASAP7_75t_L g866 ( .A1(n_835), .A2(n_745), .B(n_682), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_853), .B(n_804), .Y(n_867) );
O2A1O1Ixp33_ASAP7_75t_SL g868 ( .A1(n_860), .A2(n_839), .B(n_847), .C(n_845), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_856), .A2(n_834), .B1(n_850), .B2(n_851), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_863), .A2(n_855), .B1(n_864), .B2(n_854), .C(n_857), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_858), .Y(n_871) );
OAI221xp5_ASAP7_75t_SL g872 ( .A1(n_865), .A2(n_843), .B1(n_842), .B2(n_773), .C(n_771), .Y(n_872) );
NAND3xp33_ASAP7_75t_L g873 ( .A(n_866), .B(n_827), .C(n_747), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_862), .B(n_786), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_861), .A2(n_751), .B1(n_756), .B2(n_782), .Y(n_875) );
OAI211xp5_ASAP7_75t_L g876 ( .A1(n_866), .A2(n_690), .B(n_676), .C(n_700), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_867), .A2(n_784), .B1(n_656), .B2(n_658), .Y(n_877) );
OAI21xp33_ASAP7_75t_SL g878 ( .A1(n_859), .A2(n_785), .B(n_778), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_860), .A2(n_774), .B(n_772), .Y(n_879) );
AOI221xp5_ASAP7_75t_L g880 ( .A1(n_860), .A2(n_637), .B1(n_719), .B2(n_716), .C(n_718), .Y(n_880) );
OR2x2_ASAP7_75t_L g881 ( .A(n_865), .B(n_715), .Y(n_881) );
OAI21xp33_ASAP7_75t_L g882 ( .A1(n_860), .A2(n_755), .B(n_752), .Y(n_882) );
NOR3xp33_ASAP7_75t_L g883 ( .A(n_870), .B(n_868), .C(n_872), .Y(n_883) );
NAND4xp25_ASAP7_75t_L g884 ( .A(n_869), .B(n_880), .C(n_876), .D(n_879), .Y(n_884) );
A2O1A1Ixp33_ASAP7_75t_L g885 ( .A1(n_878), .A2(n_873), .B(n_882), .C(n_871), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_881), .A2(n_874), .B1(n_875), .B2(n_877), .C(n_722), .Y(n_886) );
NOR3xp33_ASAP7_75t_L g887 ( .A(n_883), .B(n_705), .C(n_720), .Y(n_887) );
NOR2x1_ASAP7_75t_L g888 ( .A(n_884), .B(n_715), .Y(n_888) );
NAND4xp25_ASAP7_75t_L g889 ( .A(n_885), .B(n_223), .C(n_224), .D(n_225), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_888), .Y(n_890) );
XOR2x2_ASAP7_75t_L g891 ( .A(n_887), .B(n_886), .Y(n_891) );
XOR2x2_ASAP7_75t_L g892 ( .A(n_889), .B(n_226), .Y(n_892) );
INVx3_ASAP7_75t_L g893 ( .A(n_890), .Y(n_893) );
XNOR2xp5_ASAP7_75t_L g894 ( .A(n_892), .B(n_227), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g895 ( .A1(n_893), .A2(n_891), .B1(n_230), .B2(n_231), .Y(n_895) );
XNOR2x1_ASAP7_75t_L g896 ( .A(n_894), .B(n_277), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_896), .A2(n_234), .B(n_235), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_895), .Y(n_898) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_898), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_897), .A2(n_236), .B(n_237), .Y(n_900) );
OAI21xp5_ASAP7_75t_L g901 ( .A1(n_899), .A2(n_240), .B(n_241), .Y(n_901) );
AOI21xp5_ASAP7_75t_L g902 ( .A1(n_901), .A2(n_900), .B(n_246), .Y(n_902) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_902), .A2(n_248), .B(n_249), .Y(n_903) );
endmodule