module fake_jpeg_3229_n_675 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_675);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_675;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_0),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_60),
.B(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_61),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_20),
.B(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_62),
.B(n_63),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_65),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_66),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_67),
.B(n_74),
.Y(n_200)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_69),
.Y(n_205)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_72),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_26),
.B(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_80),
.B(n_89),
.Y(n_148)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_85),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_33),
.B(n_15),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_86),
.B(n_116),
.Y(n_209)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_38),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_90),
.Y(n_216)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_91),
.Y(n_225)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

CKINVDCx9p33_ASAP7_75t_R g173 ( 
.A(n_96),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_97),
.Y(n_220)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_101),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g188 ( 
.A(n_102),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_38),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_107),
.Y(n_157)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_38),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_55),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_112),
.B(n_114),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_39),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_15),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_15),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_118),
.B(n_28),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_54),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_120),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_39),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_27),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_122),
.B(n_129),
.Y(n_189)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_43),
.B(n_49),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_29),
.Y(n_140)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_30),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_30),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_130),
.B(n_58),
.Y(n_193)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_43),
.Y(n_131)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_47),
.Y(n_132)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_72),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_134),
.A2(n_133),
.B1(n_156),
.B2(n_199),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_140),
.B(n_125),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_52),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_144),
.B(n_145),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_47),
.Y(n_145)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_146),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_147),
.B(n_150),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_152),
.B(n_2),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_153),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_73),
.A2(n_58),
.B(n_28),
.C(n_29),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_160),
.B(n_164),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_70),
.B(n_49),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_109),
.A2(n_30),
.B1(n_51),
.B2(n_50),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_169),
.A2(n_195),
.B1(n_212),
.B2(n_228),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_75),
.B(n_31),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_171),
.B(n_6),
.Y(n_277)
);

BUFx8_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_174),
.Y(n_291)
);

BUFx24_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

INVx6_ASAP7_75t_SL g182 ( 
.A(n_68),
.Y(n_182)
);

CKINVDCx12_ASAP7_75t_R g239 ( 
.A(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_111),
.A2(n_51),
.B1(n_50),
.B2(n_31),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_194),
.A2(n_218),
.B1(n_10),
.B2(n_13),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_61),
.A2(n_40),
.B1(n_35),
.B2(n_34),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_76),
.B(n_40),
.C(n_35),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_196),
.B(n_6),
.C(n_8),
.Y(n_278)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_88),
.B(n_34),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_207),
.B(n_221),
.Y(n_252)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_208),
.Y(n_288)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_66),
.A2(n_48),
.B1(n_42),
.B2(n_3),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_91),
.Y(n_213)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_95),
.Y(n_217)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_69),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_101),
.Y(n_219)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_99),
.B(n_14),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_110),
.B(n_1),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_222),
.B(n_223),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_82),
.B(n_1),
.Y(n_223)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_79),
.Y(n_226)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_84),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_94),
.Y(n_229)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

INVx3_ASAP7_75t_SL g346 ( 
.A(n_231),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_189),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_234),
.B(n_238),
.C(n_244),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_235),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_236),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_237),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_240),
.B(n_241),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_128),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_92),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_243),
.B(n_253),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_164),
.B(n_113),
.Y(n_244)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_246),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_138),
.B(n_4),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_247),
.B(n_249),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_143),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_248),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_173),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_250),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_191),
.A2(n_103),
.B1(n_85),
.B2(n_78),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_251),
.A2(n_267),
.B1(n_305),
.B2(n_311),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_159),
.B(n_108),
.Y(n_253)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_151),
.Y(n_254)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_254),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_162),
.B(n_4),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_255),
.B(n_257),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_187),
.Y(n_256)
);

INVx6_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_170),
.B(n_102),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

INVx8_ASAP7_75t_L g361 ( 
.A(n_261),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_262),
.B(n_264),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_183),
.B(n_97),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_167),
.Y(n_266)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_191),
.A2(n_106),
.B1(n_6),
.B2(n_8),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_197),
.B(n_5),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_268),
.B(n_276),
.Y(n_349)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_136),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_271),
.Y(n_343)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_151),
.Y(n_273)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_136),
.Y(n_274)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_274),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_186),
.B(n_5),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_277),
.B(n_280),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_299),
.Y(n_315)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_214),
.Y(n_279)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_145),
.B(n_9),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_205),
.Y(n_282)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_148),
.B(n_9),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_283),
.B(n_284),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_160),
.B(n_9),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_188),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_285),
.A2(n_142),
.B1(n_141),
.B2(n_185),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_157),
.B(n_10),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_286),
.B(n_294),
.Y(n_367)
);

CKINVDCx12_ASAP7_75t_R g290 ( 
.A(n_151),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_290),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_292),
.A2(n_300),
.B1(n_188),
.B2(n_224),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_211),
.Y(n_293)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_171),
.Y(n_294)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_141),
.Y(n_295)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_180),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_297),
.B(n_298),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_153),
.B(n_211),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_192),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_134),
.A2(n_220),
.B1(n_185),
.B2(n_158),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_154),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_301),
.Y(n_332)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_178),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_307),
.Y(n_334)
);

OR2x4_ASAP7_75t_L g303 ( 
.A(n_144),
.B(n_177),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_303),
.A2(n_227),
.B(n_146),
.Y(n_359)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_215),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_304),
.Y(n_373)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_154),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_306),
.Y(n_338)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_202),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_214),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_203),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_309),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_137),
.B(n_161),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_149),
.Y(n_314)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_155),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_139),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_312),
.A2(n_174),
.B1(n_287),
.B2(n_236),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_R g389 ( 
.A(n_314),
.B(n_359),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_317),
.A2(n_323),
.B1(n_331),
.B2(n_340),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_190),
.C(n_165),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_319),
.B(n_321),
.C(n_355),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_270),
.B(n_168),
.C(n_166),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_259),
.B(n_175),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_326),
.B(n_328),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_198),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_296),
.A2(n_158),
.B1(n_220),
.B2(n_224),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g335 ( 
.A(n_303),
.B(n_133),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_335),
.B(n_306),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_292),
.A2(n_206),
.B1(n_215),
.B2(n_163),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_244),
.A2(n_206),
.B1(n_163),
.B2(n_156),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_341),
.A2(n_342),
.B1(n_293),
.B2(n_237),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_275),
.A2(n_201),
.B1(n_225),
.B2(n_216),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_278),
.B(n_179),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_368),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_287),
.A2(n_142),
.B1(n_139),
.B2(n_184),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_354),
.A2(n_372),
.B1(n_291),
.B2(n_269),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_281),
.B(n_184),
.C(n_201),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_252),
.A2(n_227),
.B1(n_208),
.B2(n_177),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_357),
.A2(n_362),
.B1(n_335),
.B2(n_317),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_298),
.A2(n_251),
.B(n_267),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_362),
.A2(n_254),
.B(n_273),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_245),
.B(n_311),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_289),
.B(n_233),
.C(n_266),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_248),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_272),
.B(n_265),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_269),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_258),
.A2(n_265),
.B1(n_260),
.B2(n_263),
.Y(n_372)
);

OA22x2_ASAP7_75t_L g375 ( 
.A1(n_333),
.A2(n_285),
.B1(n_305),
.B2(n_304),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_SL g455 ( 
.A1(n_375),
.A2(n_391),
.B(n_232),
.C(n_351),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_305),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_376),
.A2(n_315),
.B(n_341),
.Y(n_438)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_371),
.Y(n_377)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_377),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_378),
.A2(n_402),
.B1(n_410),
.B2(n_416),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_R g379 ( 
.A(n_350),
.B(n_326),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_387),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_349),
.B(n_316),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_380),
.B(n_381),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_356),
.B(n_308),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_242),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_383),
.Y(n_439)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_385),
.Y(n_460)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_336),
.B(n_258),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_353),
.B(n_260),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_388),
.B(n_392),
.Y(n_447)
);

OAI22x1_ASAP7_75t_SL g391 ( 
.A1(n_335),
.A2(n_271),
.B1(n_274),
.B2(n_279),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_368),
.B(n_299),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_393),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_324),
.B(n_299),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_395),
.B(n_404),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_396),
.B(n_347),
.Y(n_461)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_313),
.Y(n_397)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_397),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_334),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_407),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_401),
.A2(n_418),
.B(n_357),
.Y(n_434)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_403),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_374),
.B(n_231),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_406),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_301),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_322),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_409),
.Y(n_433)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx13_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_320),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_412),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_295),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_330),
.B(n_246),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_414),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_318),
.B(n_250),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_314),
.B(n_256),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_419),
.Y(n_451)
);

INVx13_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_315),
.A2(n_261),
.B1(n_282),
.B2(n_235),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_417),
.A2(n_331),
.B1(n_340),
.B2(n_346),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_328),
.A2(n_239),
.B(n_230),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_321),
.B(n_230),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_420),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_334),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_421),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_422),
.A2(n_421),
.B1(n_399),
.B2(n_420),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_366),
.B(n_334),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_347),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_430),
.A2(n_431),
.B1(n_452),
.B2(n_435),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_394),
.A2(n_400),
.B1(n_376),
.B2(n_377),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_400),
.A2(n_315),
.B1(n_319),
.B2(n_323),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_435),
.A2(n_459),
.B1(n_464),
.B2(n_396),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_438),
.A2(n_453),
.B(n_375),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_378),
.A2(n_342),
.B1(n_373),
.B2(n_363),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_441),
.A2(n_450),
.B1(n_462),
.B2(n_411),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_355),
.C(n_320),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_417),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_376),
.A2(n_373),
.B1(n_363),
.B2(n_338),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_394),
.A2(n_351),
.B1(n_338),
.B2(n_332),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_389),
.A2(n_332),
.B(n_366),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_454),
.B(n_395),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_455),
.A2(n_343),
.B1(n_291),
.B2(n_339),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_401),
.A2(n_327),
.B(n_352),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_457),
.A2(n_463),
.B(n_382),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_458),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_405),
.A2(n_346),
.B1(n_358),
.B2(n_364),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_449),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_390),
.A2(n_346),
.B1(n_343),
.B2(n_364),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_398),
.A2(n_327),
.B(n_352),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_390),
.A2(n_358),
.B1(n_361),
.B2(n_337),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_381),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_465),
.B(n_476),
.Y(n_535)
);

CKINVDCx10_ASAP7_75t_R g466 ( 
.A(n_463),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_466),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_436),
.B(n_388),
.Y(n_467)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_467),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_468),
.A2(n_495),
.B1(n_430),
.B2(n_462),
.Y(n_524)
);

INVx6_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_469),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_470),
.B(n_475),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_SL g508 ( 
.A(n_471),
.B(n_478),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_425),
.B(n_380),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_472),
.B(n_483),
.Y(n_513)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_473),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_427),
.A2(n_415),
.B1(n_375),
.B2(n_392),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_479),
.B1(n_431),
.B2(n_438),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_419),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_379),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_437),
.Y(n_477)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_477),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_453),
.A2(n_382),
.B(n_418),
.Y(n_478)
);

NOR3xp33_ASAP7_75t_SL g480 ( 
.A(n_443),
.B(n_398),
.C(n_391),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_480),
.B(n_499),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_481),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_482),
.B(n_491),
.C(n_452),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_439),
.B(n_329),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_484),
.A2(n_490),
.B(n_455),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_425),
.B(n_329),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_485),
.B(n_486),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_348),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_433),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_487),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_489),
.B(n_454),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_434),
.A2(n_375),
.B(n_406),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_397),
.Y(n_491)
);

INVx13_ASAP7_75t_L g492 ( 
.A(n_457),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_492),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_433),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_493),
.Y(n_534)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_494),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_427),
.A2(n_384),
.B1(n_409),
.B2(n_408),
.Y(n_495)
);

INVx13_ASAP7_75t_L g496 ( 
.A(n_455),
.Y(n_496)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_496),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_436),
.B(n_386),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_428),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_498),
.A2(n_432),
.B(n_424),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_426),
.B(n_403),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_437),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_502),
.Y(n_506)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_504),
.A2(n_511),
.B1(n_519),
.B2(n_524),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_451),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_505),
.B(n_514),
.C(n_517),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_472),
.B(n_460),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_512),
.B(n_518),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_491),
.B(n_447),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_516),
.A2(n_471),
.B(n_484),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_460),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_479),
.A2(n_428),
.B1(n_441),
.B2(n_450),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_477),
.B(n_456),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_520),
.B(n_528),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_482),
.B(n_447),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_531),
.C(n_538),
.Y(n_553)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_522),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_499),
.B(n_456),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_481),
.B(n_468),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_470),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_490),
.A2(n_488),
.B1(n_500),
.B2(n_467),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_536),
.A2(n_455),
.B1(n_492),
.B2(n_496),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_469),
.B(n_443),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_537),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_459),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_541),
.B(n_544),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_505),
.B(n_500),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_522),
.B(n_497),
.Y(n_545)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_545),
.Y(n_575)
);

BUFx24_ASAP7_75t_SL g546 ( 
.A(n_535),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_546),
.B(n_510),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_513),
.B(n_448),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_547),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_548),
.A2(n_559),
.B(n_508),
.Y(n_576)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_506),
.Y(n_549)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_549),
.Y(n_577)
);

BUFx2_ASAP7_75t_SL g550 ( 
.A(n_526),
.Y(n_550)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_550),
.Y(n_573)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_523),
.Y(n_554)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_554),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_503),
.A2(n_487),
.B1(n_493),
.B2(n_495),
.Y(n_555)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_555),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_517),
.B(n_474),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_556),
.B(n_570),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_502),
.C(n_494),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_557),
.B(n_561),
.C(n_562),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_536),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_558),
.B(n_567),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_509),
.A2(n_466),
.B(n_492),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_473),
.C(n_445),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_514),
.B(n_445),
.C(n_444),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_563),
.A2(n_539),
.B1(n_525),
.B2(n_527),
.Y(n_587)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_523),
.Y(n_564)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_564),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_513),
.B(n_530),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_565),
.B(n_566),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_515),
.B(n_446),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_509),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_504),
.A2(n_475),
.B1(n_496),
.B2(n_480),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_568),
.A2(n_569),
.B1(n_516),
.B2(n_534),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_519),
.A2(n_455),
.B1(n_446),
.B2(n_440),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_532),
.B(n_464),
.Y(n_570)
);

XNOR2x1_ASAP7_75t_L g571 ( 
.A(n_544),
.B(n_538),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_571),
.B(n_585),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_572),
.A2(n_548),
.B1(n_567),
.B2(n_559),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_581),
.B(n_562),
.Y(n_612)
);

NOR3xp33_ASAP7_75t_L g584 ( 
.A(n_542),
.B(n_545),
.C(n_543),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_584),
.B(n_586),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_SL g585 ( 
.A(n_553),
.B(n_503),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_560),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_587),
.A2(n_593),
.B1(n_563),
.B2(n_569),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_552),
.A2(n_534),
.B1(n_527),
.B2(n_507),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_588),
.A2(n_529),
.B1(n_568),
.B2(n_533),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_551),
.B(n_525),
.C(n_526),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_589),
.Y(n_607)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_570),
.Y(n_590)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_590),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_558),
.A2(n_507),
.B1(n_511),
.B2(n_539),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_SL g594 ( 
.A(n_553),
.B(n_515),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_594),
.B(n_551),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_588),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_596),
.B(n_597),
.Y(n_621)
);

CKINVDCx14_ASAP7_75t_R g597 ( 
.A(n_582),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_589),
.B(n_540),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_600),
.B(n_603),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_602),
.B(n_609),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_SL g603 ( 
.A(n_575),
.B(n_577),
.C(n_583),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_573),
.Y(n_604)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_604),
.Y(n_620)
);

INVx13_ASAP7_75t_L g605 ( 
.A(n_573),
.Y(n_605)
);

INVx11_ASAP7_75t_L g619 ( 
.A(n_605),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_606),
.A2(n_574),
.B(n_576),
.Y(n_626)
);

BUFx24_ASAP7_75t_SL g608 ( 
.A(n_592),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_608),
.B(n_599),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_580),
.B(n_557),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_580),
.B(n_556),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_610),
.B(n_595),
.Y(n_618)
);

INVxp33_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_611),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_612),
.B(n_616),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_614),
.A2(n_615),
.B1(n_593),
.B2(n_572),
.Y(n_622)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_578),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_618),
.B(n_624),
.Y(n_635)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_622),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_607),
.B(n_609),
.C(n_610),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_602),
.B(n_595),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_625),
.B(n_630),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_626),
.A2(n_627),
.B1(n_529),
.B2(n_533),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_606),
.A2(n_613),
.B1(n_611),
.B2(n_598),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_613),
.B(n_594),
.C(n_579),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_601),
.B(n_579),
.C(n_590),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_631),
.B(n_618),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_632),
.B(n_440),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_603),
.A2(n_587),
.B(n_541),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_633),
.A2(n_339),
.B(n_385),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_628),
.A2(n_591),
.B1(n_561),
.B2(n_585),
.Y(n_634)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_634),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_627),
.A2(n_571),
.B1(n_601),
.B2(n_605),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_638),
.B(n_640),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_639),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_626),
.A2(n_621),
.B(n_623),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_SL g648 ( 
.A1(n_641),
.A2(n_620),
.B(n_619),
.Y(n_648)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_629),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_642),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_643),
.A2(n_644),
.B(n_647),
.Y(n_655)
);

NOR2x1_ASAP7_75t_L g644 ( 
.A(n_630),
.B(n_622),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_645),
.B(n_646),
.Y(n_649)
);

INVx11_ASAP7_75t_L g646 ( 
.A(n_619),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_633),
.A2(n_393),
.B(n_385),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_648),
.A2(n_650),
.B(n_647),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_635),
.A2(n_624),
.B(n_617),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_SL g653 ( 
.A(n_636),
.B(n_617),
.Y(n_653)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_653),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_644),
.Y(n_656)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_656),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_651),
.B(n_637),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_658),
.B(n_659),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_654),
.B(n_641),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_660),
.A2(n_661),
.B(n_662),
.Y(n_665)
);

AOI322xp5_ASAP7_75t_L g661 ( 
.A1(n_657),
.A2(n_646),
.A3(n_640),
.B1(n_638),
.B2(n_645),
.C1(n_631),
.C2(n_625),
.Y(n_661)
);

AOI211xp5_ASAP7_75t_L g662 ( 
.A1(n_652),
.A2(n_393),
.B(n_385),
.C(n_410),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_664),
.B(n_649),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_666),
.B(n_667),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_661),
.A2(n_655),
.B(n_657),
.Y(n_667)
);

NOR3xp33_ASAP7_75t_SL g670 ( 
.A(n_668),
.B(n_663),
.C(n_665),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_670),
.B(n_250),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_671),
.B(n_669),
.C(n_365),
.Y(n_672)
);

AO21x1_ASAP7_75t_L g673 ( 
.A1(n_672),
.A2(n_365),
.B(n_416),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_SL g674 ( 
.A1(n_673),
.A2(n_348),
.B1(n_232),
.B2(n_288),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_674),
.B(n_288),
.C(n_173),
.Y(n_675)
);


endmodule