module fake_aes_7679_n_26 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
AOI22xp5_ASAP7_75t_L g14 ( .A1(n_8), .A2(n_10), .B1(n_2), .B2(n_12), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_9), .B(n_1), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_11), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
A2O1A1Ixp33_ASAP7_75t_L g19 ( .A1(n_15), .A2(n_0), .B(n_2), .C(n_3), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_18), .B(n_13), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_16), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_22), .B(n_19), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_14), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_15), .B1(n_3), .B2(n_0), .Y(n_25) );
OAI31xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_4), .A3(n_5), .B(n_6), .Y(n_26) );
endmodule