module fake_netlist_1_409_n_42 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_2), .B(n_8), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_7), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_6), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_12), .B(n_0), .Y(n_20) );
NOR3xp33_ASAP7_75t_SL g21 ( .A(n_18), .B(n_0), .C(n_1), .Y(n_21) );
BUFx2_ASAP7_75t_L g22 ( .A(n_12), .Y(n_22) );
CKINVDCx11_ASAP7_75t_R g23 ( .A(n_17), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_11), .Y(n_24) );
NAND2xp33_ASAP7_75t_R g25 ( .A(n_22), .B(n_18), .Y(n_25) );
INVx3_ASAP7_75t_L g26 ( .A(n_19), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_20), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_22), .A2(n_16), .B1(n_3), .B2(n_4), .Y(n_28) );
OAI332xp33_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_24), .A3(n_19), .B1(n_23), .B2(n_21), .B3(n_1), .C1(n_7), .C2(n_4), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_26), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_26), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_27), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_33), .B(n_29), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
NAND4xp75_ASAP7_75t_L g36 ( .A(n_34), .B(n_33), .C(n_24), .D(n_32), .Y(n_36) );
OAI211xp5_ASAP7_75t_SL g37 ( .A1(n_35), .A2(n_28), .B(n_31), .C(n_30), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_35), .B(n_33), .Y(n_38) );
OR3x2_ASAP7_75t_L g39 ( .A(n_36), .B(n_3), .C(n_9), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
AOI22xp33_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_37), .B1(n_40), .B2(n_34), .Y(n_41) );
BUFx2_ASAP7_75t_L g42 ( .A(n_41), .Y(n_42) );
endmodule