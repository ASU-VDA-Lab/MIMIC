module fake_jpeg_27569_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_38),
.Y(n_51)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g39 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_2),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_26),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_44),
.B(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_32),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_22),
.B1(n_30),
.B2(n_25),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_57),
.B1(n_38),
.B2(n_31),
.Y(n_86)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_16),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_30),
.B1(n_25),
.B2(n_29),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_35),
.B1(n_38),
.B2(n_36),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_30),
.B1(n_25),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_41),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_29),
.B1(n_27),
.B2(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_57),
.B1(n_45),
.B2(n_42),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_28),
.B1(n_20),
.B2(n_24),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_67),
.B(n_75),
.Y(n_98)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_65),
.B(n_68),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_72),
.Y(n_93)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_76),
.B(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_37),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_21),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_33),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_38),
.B1(n_36),
.B2(n_31),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_86),
.B1(n_82),
.B2(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_32),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_66),
.B1(n_77),
.B2(n_68),
.Y(n_134)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_109),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_97),
.B(n_107),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_43),
.B(n_44),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_103),
.B(n_98),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_69),
.A2(n_43),
.B(n_47),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_110),
.B(n_78),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_60),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_45),
.B(n_58),
.C(n_49),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_58),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_58),
.B1(n_45),
.B2(n_42),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_120),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_64),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_115),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_64),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_124),
.B(n_125),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_131),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_71),
.C(n_67),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_19),
.C(n_50),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_132),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_65),
.B(n_74),
.C(n_73),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_137),
.B(n_89),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_100),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_112),
.B1(n_107),
.B2(n_94),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_81),
.B1(n_66),
.B2(n_63),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_92),
.A2(n_77),
.B1(n_17),
.B2(n_24),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_100),
.B1(n_95),
.B2(n_105),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_33),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_91),
.B(n_21),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_156),
.B(n_159),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_152),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_160),
.B1(n_126),
.B2(n_19),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_3),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_87),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_154),
.B(n_155),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_89),
.B(n_87),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_106),
.B(n_105),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_108),
.B1(n_19),
.B2(n_33),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_4),
.C(n_5),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_19),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_123),
.A3(n_122),
.B1(n_135),
.B2(n_128),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_143),
.A3(n_154),
.B1(n_161),
.B2(n_144),
.C1(n_146),
.C2(n_15),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_176),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_159),
.B1(n_152),
.B2(n_146),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_3),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_4),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_4),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_9),
.B(n_10),
.Y(n_202)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_162),
.C(n_139),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_179),
.A2(n_171),
.B1(n_168),
.B2(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_142),
.C(n_151),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_201),
.C(n_185),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_140),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_166),
.A2(n_144),
.B1(n_143),
.B2(n_147),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_195),
.Y(n_210)
);

AOI321xp33_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_15),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_183),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_5),
.C(n_6),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_183),
.B(n_10),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_215),
.C(n_201),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_173),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_192),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_182),
.C(n_167),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_196),
.C(n_188),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_217),
.B(n_222),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_224),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_221),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_193),
.B1(n_177),
.B2(n_190),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_215),
.B1(n_202),
.B2(n_210),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_203),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_218),
.A2(n_204),
.B1(n_208),
.B2(n_212),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_229),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_195),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_14),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_210),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_233),
.A2(n_200),
.B(n_11),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_222),
.B1(n_216),
.B2(n_225),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_234),
.A2(n_238),
.B1(n_226),
.B2(n_230),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_220),
.C(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_228),
.C(n_11),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_237),
.B(n_9),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_239),
.B(n_12),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_246),
.B(n_11),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_12),
.Y(n_250)
);


endmodule