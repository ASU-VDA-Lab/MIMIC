module fake_jpeg_18461_n_188 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_0),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_30),
.B(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_13),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_44),
.Y(n_46)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_29),
.C(n_18),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_52),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_18),
.B1(n_14),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_17),
.B1(n_25),
.B2(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_54),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_24),
.B1(n_28),
.B2(n_23),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_72),
.B1(n_27),
.B2(n_22),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_65),
.Y(n_84)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_21),
.Y(n_82)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_15),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_26),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_23),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_26),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_34),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_25),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_6),
.C(n_7),
.Y(n_97)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_97),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_88),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_69),
.B1(n_62),
.B2(n_58),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_19),
.B1(n_25),
.B2(n_3),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_95),
.B1(n_82),
.B2(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_1),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_96),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_25),
.B(n_2),
.C(n_5),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_98),
.B(n_8),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_25),
.B1(n_2),
.B2(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_70),
.B1(n_59),
.B2(n_73),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_47),
.B(n_7),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_7),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_48),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_61),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_11),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_115),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_98),
.B(n_86),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_68),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_76),
.A3(n_97),
.B1(n_92),
.B2(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_117),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_58),
.B1(n_64),
.B2(n_50),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_78),
.B1(n_57),
.B2(n_81),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_49),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_119),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_103),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_95),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_104),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_112),
.A2(n_96),
.B1(n_50),
.B2(n_75),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_136),
.B1(n_138),
.B2(n_107),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_47),
.C(n_49),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_130),
.C(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_137),
.A2(n_119),
.B1(n_111),
.B2(n_105),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_93),
.B1(n_57),
.B2(n_74),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_142),
.B1(n_143),
.B2(n_150),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_147),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_119),
.B1(n_101),
.B2(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_119),
.B(n_118),
.Y(n_147)
);

OAI22x1_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_117),
.B1(n_110),
.B2(n_108),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_131),
.B1(n_107),
.B2(n_120),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_151),
.A2(n_139),
.B1(n_137),
.B2(n_126),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_156),
.B1(n_159),
.B2(n_150),
.Y(n_164)
);

AO32x1_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_133),
.A3(n_122),
.B1(n_124),
.B2(n_128),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_122),
.B(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_143),
.C(n_144),
.Y(n_162)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_163),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_166),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_145),
.B(n_142),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_157),
.B(n_158),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_140),
.C(n_152),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_148),
.C(n_135),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_148),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_161),
.B1(n_162),
.B2(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_160),
.B(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_173),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_180),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_167),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_170),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_178),
.A2(n_171),
.B(n_175),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_183),
.B(n_178),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_185),
.B(n_169),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_173),
.Y(n_188)
);


endmodule