module fake_aes_10596_n_659 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_659);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_659;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_617;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_597;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_3), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_55), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_31), .Y(n_77) );
NOR2xp67_ASAP7_75t_L g78 ( .A(n_33), .B(n_72), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_67), .Y(n_79) );
INVx1_ASAP7_75t_SL g80 ( .A(n_62), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_20), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_39), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_27), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_69), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_24), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_12), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_35), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_47), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_32), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_18), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_10), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
BUFx8_ASAP7_75t_SL g93 ( .A(n_65), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_68), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_42), .Y(n_95) );
CKINVDCx14_ASAP7_75t_R g96 ( .A(n_23), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_37), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_25), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_74), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_16), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_34), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_21), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_5), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_48), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_14), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_1), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_60), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_36), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_61), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_52), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_17), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_2), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_64), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_57), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_7), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_5), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_12), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_94), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_118), .B(n_0), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_118), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_94), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_81), .B(n_4), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_117), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_100), .Y(n_128) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_117), .A2(n_43), .B(n_71), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_108), .B(n_6), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_100), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
INVx5_ASAP7_75t_L g134 ( .A(n_93), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
AOI22xp5_ASAP7_75t_SL g136 ( .A1(n_115), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_86), .B(n_8), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_116), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_76), .Y(n_140) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_79), .A2(n_44), .B(n_70), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
INVx5_ASAP7_75t_L g143 ( .A(n_96), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_106), .B(n_9), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_106), .B(n_9), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_82), .B(n_11), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_83), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_89), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_90), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_99), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_75), .B(n_13), .Y(n_152) );
OA21x2_ASAP7_75t_L g153 ( .A1(n_102), .A2(n_45), .B(n_66), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_104), .B(n_13), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_109), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_112), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_98), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_91), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_92), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_103), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
INVxp67_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
INVx4_ASAP7_75t_SL g164 ( .A(n_122), .Y(n_164) );
NAND3xp33_ASAP7_75t_L g165 ( .A(n_124), .B(n_105), .C(n_107), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_158), .B(n_77), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_152), .A2(n_110), .B1(n_120), .B2(n_77), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_158), .B(n_95), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_158), .B(n_78), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_158), .B(n_143), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_134), .Y(n_174) );
NAND2xp33_ASAP7_75t_L g175 ( .A(n_143), .B(n_84), .Y(n_175) );
OR2x6_ASAP7_75t_L g176 ( .A(n_122), .B(n_115), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_128), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_158), .B(n_95), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_158), .B(n_111), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_126), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_134), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_151), .B(n_111), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_137), .B(n_84), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_128), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_152), .B(n_80), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
INVx1_ASAP7_75t_SL g190 ( .A(n_134), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_160), .B(n_14), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_151), .B(n_114), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_143), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_161), .B(n_114), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_133), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_133), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_124), .B(n_88), .Y(n_198) );
BUFx8_ASAP7_75t_SL g199 ( .A(n_148), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_128), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_130), .B(n_101), .Y(n_201) );
INVx4_ASAP7_75t_SL g202 ( .A(n_128), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_130), .B(n_119), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_148), .B(n_88), .Y(n_204) );
INVx5_ASAP7_75t_L g205 ( .A(n_140), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_138), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_134), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_129), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_138), .Y(n_210) );
OR2x2_ASAP7_75t_L g211 ( .A(n_160), .B(n_161), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_148), .B(n_101), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_135), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_147), .Y(n_215) );
BUFx4f_ASAP7_75t_L g216 ( .A(n_139), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_123), .A2(n_119), .B1(n_15), .B2(n_22), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_143), .B(n_49), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_123), .A2(n_15), .B1(n_19), .B2(n_26), .Y(n_219) );
NOR2xp67_ASAP7_75t_L g220 ( .A(n_217), .B(n_148), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_185), .A2(n_129), .B(n_141), .Y(n_221) );
NOR3xp33_ASAP7_75t_L g222 ( .A(n_195), .B(n_145), .C(n_144), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_183), .B(n_139), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_187), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_216), .B(n_135), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_209), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_180), .B(n_147), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_215), .B(n_143), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_163), .B(n_147), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_180), .B(n_143), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_176), .B(n_131), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_201), .A2(n_146), .B1(n_154), .B2(n_149), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_191), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_184), .A2(n_149), .B1(n_138), .B2(n_159), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_SL g235 ( .A1(n_168), .A2(n_149), .B(n_159), .C(n_127), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_196), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_184), .B(n_159), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_211), .B(n_142), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_204), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_192), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_207), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_216), .B(n_142), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_187), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_208), .B(n_135), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_204), .B(n_125), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_197), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_208), .B(n_135), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_168), .A2(n_121), .B1(n_135), .B2(n_127), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_166), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_208), .B(n_135), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_181), .B(n_179), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_193), .A2(n_136), .B1(n_125), .B2(n_121), .Y(n_252) );
INVx4_ASAP7_75t_L g253 ( .A(n_164), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_188), .A2(n_121), .B1(n_156), .B2(n_155), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_206), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_210), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_170), .B(n_157), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_213), .B(n_157), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_213), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_188), .A2(n_157), .B1(n_156), .B2(n_155), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_188), .A2(n_157), .B1(n_156), .B2(n_155), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_169), .B(n_157), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_203), .B(n_157), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_188), .A2(n_156), .B1(n_155), .B2(n_150), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_165), .A2(n_156), .B1(n_155), .B2(n_150), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_165), .A2(n_153), .B(n_141), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_164), .Y(n_267) );
NOR2x2_ASAP7_75t_L g268 ( .A(n_176), .B(n_153), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_172), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_172), .B(n_155), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_167), .B(n_156), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_176), .B(n_150), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_198), .A2(n_150), .B1(n_140), .B2(n_132), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_199), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_178), .B(n_150), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_203), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_219), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_219), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_214), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_214), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_259), .A2(n_217), .B(n_150), .C(n_140), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_239), .B(n_198), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_229), .B(n_227), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_221), .A2(n_173), .B(n_175), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_277), .A2(n_198), .B1(n_140), .B2(n_132), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_274), .Y(n_287) );
INVxp67_ASAP7_75t_SL g288 ( .A(n_276), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_229), .B(n_198), .Y(n_289) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_278), .B(n_153), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_252), .A2(n_182), .B(n_190), .C(n_189), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_231), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_262), .A2(n_182), .B(n_190), .C(n_218), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_253), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_240), .A2(n_174), .B1(n_140), .B2(n_132), .Y(n_296) );
BUFx4f_ASAP7_75t_L g297 ( .A(n_231), .Y(n_297) );
INVx5_ASAP7_75t_L g298 ( .A(n_253), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_237), .B(n_140), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_238), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_226), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_231), .B(n_132), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_272), .B(n_132), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_237), .A2(n_212), .B(n_162), .C(n_171), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_251), .A2(n_186), .B(n_177), .C(n_200), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_234), .A2(n_194), .B1(n_153), .B2(n_141), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_241), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_224), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_241), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_251), .A2(n_205), .B(n_141), .C(n_202), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_220), .A2(n_205), .B1(n_194), .B2(n_202), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_222), .B(n_205), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_244), .A2(n_28), .B(n_29), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_223), .B(n_30), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_249), .Y(n_315) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_232), .A2(n_38), .B1(n_40), .B2(n_41), .C(n_46), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_233), .Y(n_317) );
O2A1O1Ixp5_ASAP7_75t_L g318 ( .A1(n_266), .A2(n_73), .B(n_51), .C(n_53), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_226), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_243), .B(n_50), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_262), .A2(n_245), .B(n_258), .C(n_235), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_244), .A2(n_54), .B(n_56), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_243), .B(n_269), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_236), .Y(n_324) );
BUFx2_ASAP7_75t_SL g325 ( .A(n_246), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_267), .B(n_63), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_242), .B(n_58), .Y(n_327) );
NOR2xp33_ASAP7_75t_SL g328 ( .A(n_297), .B(n_255), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_317), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_287), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_281), .A2(n_256), .B(n_257), .C(n_235), .Y(n_331) );
AO31x2_ASAP7_75t_L g332 ( .A1(n_310), .A2(n_257), .A3(n_271), .B(n_275), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_324), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_300), .A2(n_248), .B1(n_273), .B2(n_230), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_297), .Y(n_335) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_283), .A2(n_270), .B(n_225), .C(n_228), .Y(n_336) );
AOI221x1_ASAP7_75t_L g337 ( .A1(n_306), .A2(n_268), .B1(n_273), .B2(n_254), .C(n_264), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_298), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_325), .A2(n_270), .B1(n_225), .B2(n_261), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_292), .B(n_247), .Y(n_341) );
AO21x1_ASAP7_75t_L g342 ( .A1(n_321), .A2(n_247), .B(n_250), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_284), .A2(n_250), .B(n_279), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g345 ( .A1(n_291), .A2(n_260), .B(n_248), .C(n_265), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_314), .A2(n_280), .B(n_265), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_313), .A2(n_59), .B(n_318), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_323), .B(n_288), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_288), .A2(n_285), .B1(n_307), .B2(n_309), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_298), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_282), .A2(n_295), .B1(n_308), .B2(n_289), .Y(n_351) );
INVx3_ASAP7_75t_SL g352 ( .A(n_298), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_318), .A2(n_293), .B(n_322), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_290), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_327), .A2(n_286), .B1(n_295), .B2(n_308), .Y(n_355) );
AOI21x1_ASAP7_75t_L g356 ( .A1(n_320), .A2(n_299), .B(n_296), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_L g357 ( .A1(n_355), .A2(n_312), .B(n_302), .C(n_316), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_343), .A2(n_286), .B1(n_311), .B2(n_304), .C(n_305), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_344), .A2(n_290), .B(n_303), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_329), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_348), .B(n_294), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_349), .A2(n_294), .B(n_326), .C(n_319), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_335), .B(n_301), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_331), .A2(n_301), .B(n_319), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_348), .B(n_301), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_333), .B(n_301), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_353), .A2(n_319), .B(n_347), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_354), .B(n_319), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_328), .B(n_341), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_346), .A2(n_331), .B(n_342), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_336), .B(n_334), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_354), .A2(n_341), .B1(n_350), .B2(n_352), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_332), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_352), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_345), .A2(n_337), .B(n_351), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_345), .A2(n_340), .B(n_339), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_332), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_332), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_332), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_361), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_374), .A2(n_350), .B1(n_339), .B2(n_338), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_361), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_358), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_364), .B(n_356), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_364), .B(n_330), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_376), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_358), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_379), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_369), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_376), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_369), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_376), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_376), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_376), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_379), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_370), .B(n_380), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_362), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_368), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_362), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_381), .B(n_382), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_370), .B(n_380), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_367), .Y(n_407) );
OR2x6_ASAP7_75t_L g408 ( .A(n_378), .B(n_360), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_368), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_366), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_381), .B(n_382), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_365), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_372), .A2(n_373), .B(n_357), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_371), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_359), .A2(n_363), .B1(n_377), .B2(n_375), .C(n_381), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_412), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_391), .B(n_382), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_388), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_391), .B(n_375), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_407), .B(n_377), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_389), .B(n_366), .Y(n_422) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_411), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_388), .A2(n_404), .B1(n_401), .B2(n_415), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_389), .B(n_405), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_392), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_392), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_388), .B(n_394), .Y(n_429) );
NAND2x1_ASAP7_75t_L g430 ( .A(n_399), .B(n_402), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_411), .B(n_405), .Y(n_431) );
INVx5_ASAP7_75t_SL g432 ( .A(n_388), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_402), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_389), .B(n_383), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_407), .B(n_383), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_398), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_411), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_411), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_385), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_385), .B(n_386), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_387), .Y(n_443) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_386), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_403), .B(n_409), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_387), .B(n_413), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_400), .B(n_406), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_400), .B(n_406), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_400), .B(n_406), .Y(n_449) );
OAI21xp33_ASAP7_75t_L g450 ( .A1(n_414), .A2(n_408), .B(n_416), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_390), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_400), .B(n_406), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_410), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_403), .B(n_409), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_397), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_410), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_408), .B(n_397), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_396), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_408), .B(n_397), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_408), .B(n_397), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_393), .Y(n_461) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_395), .A2(n_413), .B(n_410), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_384), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_408), .Y(n_464) );
INVxp33_ASAP7_75t_L g465 ( .A(n_395), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_417), .B(n_454), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_434), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_454), .B(n_426), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_427), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_431), .B(n_426), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_431), .B(n_443), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_431), .B(n_443), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_431), .B(n_439), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_439), .B(n_440), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_439), .B(n_440), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_440), .B(n_424), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_424), .B(n_449), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_421), .B(n_437), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_430), .B(n_434), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_424), .B(n_449), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_424), .B(n_447), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_433), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_464), .B(n_460), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_432), .B(n_429), .Y(n_485) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_450), .B(n_419), .C(n_463), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_447), .B(n_428), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_428), .B(n_446), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_433), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_428), .B(n_446), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_453), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_435), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_435), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_432), .B(n_425), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_441), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_451), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_441), .B(n_437), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_453), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_434), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_425), .B(n_442), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_421), .B(n_448), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_436), .Y(n_502) );
NOR2x1_ASAP7_75t_L g503 ( .A(n_430), .B(n_451), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_436), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_456), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_446), .B(n_418), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_464), .B(n_460), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_455), .B(n_438), .Y(n_508) );
NOR2xp67_ASAP7_75t_L g509 ( .A(n_438), .B(n_456), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_446), .B(n_418), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_442), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_452), .B(n_445), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_420), .B(n_457), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_420), .B(n_457), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_445), .B(n_432), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_422), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_459), .B(n_422), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_459), .B(n_444), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_432), .B(n_458), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_464), .B(n_455), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_462), .B(n_461), .Y(n_521) );
NAND2x1_ASAP7_75t_SL g522 ( .A(n_509), .B(n_503), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_495), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_517), .B(n_465), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_495), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_469), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_517), .B(n_462), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_467), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_468), .B(n_432), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_505), .Y(n_530) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_503), .B(n_462), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_509), .B(n_423), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_469), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_471), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_513), .B(n_462), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_501), .B(n_461), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_501), .B(n_461), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_466), .B(n_450), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_511), .B(n_423), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_479), .B(n_423), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_511), .B(n_423), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_470), .B(n_423), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_513), .B(n_423), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_514), .B(n_510), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_505), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_471), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_486), .A2(n_494), .B1(n_472), .B2(n_473), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_514), .B(n_510), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_506), .B(n_472), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_470), .B(n_487), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_480), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_483), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_505), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_483), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
NOR2x1_ASAP7_75t_L g556 ( .A(n_485), .B(n_499), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_489), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_506), .B(n_473), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_480), .B(n_508), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_487), .B(n_474), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_474), .B(n_488), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_492), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_479), .B(n_512), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_512), .B(n_500), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
NOR2x1_ASAP7_75t_L g566 ( .A(n_519), .B(n_515), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_520), .A2(n_496), .B1(n_518), .B2(n_478), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_520), .A2(n_484), .B(n_507), .C(n_497), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_518), .A2(n_482), .B1(n_481), .B2(n_478), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_516), .B(n_504), .Y(n_570) );
INVx1_ASAP7_75t_SL g571 ( .A(n_528), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_563), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_560), .B(n_481), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_564), .B(n_516), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_538), .B(n_504), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_570), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_523), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_538), .B(n_502), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_525), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_526), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_533), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_530), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_534), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_535), .B(n_502), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_560), .B(n_482), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_549), .B(n_490), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_546), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_552), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_527), .B(n_490), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_554), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_527), .B(n_488), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_555), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_557), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_562), .Y(n_595) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_547), .A2(n_507), .B(n_484), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_544), .B(n_493), .Y(n_597) );
NOR2xp33_ASAP7_75t_SL g598 ( .A(n_568), .B(n_480), .Y(n_598) );
AOI21xp33_ASAP7_75t_SL g599 ( .A1(n_559), .A2(n_508), .B(n_507), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_544), .B(n_493), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_536), .B(n_475), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_549), .B(n_477), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_558), .B(n_477), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_530), .Y(n_604) );
AO22x1_ASAP7_75t_L g605 ( .A1(n_571), .A2(n_556), .B1(n_551), .B2(n_566), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_583), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_582), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_582), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_572), .B(n_548), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_588), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_588), .Y(n_611) );
OAI22xp33_ASAP7_75t_SL g612 ( .A1(n_598), .A2(n_559), .B1(n_551), .B2(n_532), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_575), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_585), .B(n_537), .Y(n_614) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_581), .Y(n_615) );
AND2x4_ASAP7_75t_L g616 ( .A(n_573), .B(n_568), .Y(n_616) );
AOI21xp5_ASAP7_75t_SL g617 ( .A1(n_596), .A2(n_532), .B(n_522), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_578), .B(n_548), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_577), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_599), .A2(n_547), .B(n_551), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_576), .A2(n_567), .B1(n_569), .B2(n_524), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_574), .A2(n_524), .B1(n_565), .B2(n_558), .C(n_543), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_585), .B(n_561), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_579), .B(n_550), .Y(n_624) );
BUFx2_ASAP7_75t_L g625 ( .A(n_601), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_605), .A2(n_600), .B(n_597), .Y(n_626) );
AOI211xp5_ASAP7_75t_SL g627 ( .A1(n_612), .A2(n_529), .B(n_484), .C(n_507), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_620), .A2(n_580), .B1(n_591), .B2(n_595), .C(n_594), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_613), .A2(n_531), .B(n_593), .Y(n_629) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_616), .A2(n_484), .B1(n_586), .B2(n_573), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_625), .A2(n_590), .B1(n_601), .B2(n_592), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_617), .A2(n_586), .B(n_584), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_618), .B(n_590), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g634 ( .A(n_622), .B(n_621), .C(n_623), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_616), .A2(n_542), .B1(n_543), .B2(n_589), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_619), .A2(n_540), .B(n_541), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_622), .B(n_587), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_615), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_627), .A2(n_609), .B(n_624), .C(n_614), .Y(n_639) );
NAND4xp25_ASAP7_75t_SL g640 ( .A(n_632), .B(n_624), .C(n_587), .D(n_603), .Y(n_640) );
NAND4xp75_ASAP7_75t_L g641 ( .A(n_637), .B(n_611), .C(n_610), .D(n_608), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_634), .A2(n_607), .B(n_606), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_638), .A2(n_603), .B1(n_602), .B2(n_561), .Y(n_643) );
AOI211xp5_ASAP7_75t_L g644 ( .A1(n_628), .A2(n_602), .B(n_539), .C(n_604), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_631), .A2(n_604), .B1(n_583), .B2(n_553), .C(n_545), .Y(n_645) );
NAND5xp2_ASAP7_75t_L g646 ( .A(n_639), .B(n_630), .C(n_626), .D(n_629), .E(n_635), .Y(n_646) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_640), .B(n_633), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_642), .B(n_636), .C(n_553), .Y(n_648) );
OAI321xp33_ASAP7_75t_L g649 ( .A1(n_644), .A2(n_508), .A3(n_545), .B1(n_521), .B2(n_498), .C(n_491), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_648), .B(n_643), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_647), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_651), .B(n_646), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_650), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_653), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_652), .B1(n_645), .B2(n_649), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_655), .A2(n_652), .B(n_641), .Y(n_656) );
OAI21xp33_ASAP7_75t_SL g657 ( .A1(n_656), .A2(n_521), .B(n_491), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_657), .B(n_498), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_658), .A2(n_475), .B1(n_476), .B2(n_652), .Y(n_659) );
endmodule