module fake_ariane_461_n_54 (n_8, n_3, n_2, n_11, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_10, n_54);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;
input n_10;

output n_54;

wire n_24;
wire n_22;
wire n_43;
wire n_49;
wire n_13;
wire n_20;
wire n_27;
wire n_48;
wire n_29;
wire n_17;
wire n_41;
wire n_50;
wire n_38;
wire n_47;
wire n_18;
wire n_32;
wire n_28;
wire n_37;
wire n_51;
wire n_45;
wire n_34;
wire n_26;
wire n_46;
wire n_14;
wire n_52;
wire n_36;
wire n_33;
wire n_44;
wire n_19;
wire n_30;
wire n_39;
wire n_40;
wire n_31;
wire n_42;
wire n_16;
wire n_12;
wire n_15;
wire n_53;
wire n_21;
wire n_23;
wire n_35;
wire n_25;

INVx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_11),
.A2(n_2),
.B1(n_8),
.B2(n_0),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_3),
.B(n_6),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_3),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_12),
.B(n_18),
.C(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_21),
.Y(n_31)
);

OAI21x1_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_15),
.B(n_20),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_13),
.B(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_28),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_32),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_27),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_40),
.B(n_41),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_35),
.Y(n_46)
);

AOI31xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_26),
.A3(n_45),
.B(n_37),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_43),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

AOI222xp33_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_21),
.B1(n_39),
.B2(n_36),
.C1(n_13),
.C2(n_43),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_47),
.B1(n_36),
.B2(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_21),
.B1(n_13),
.B2(n_38),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_51),
.B(n_13),
.Y(n_54)
);


endmodule