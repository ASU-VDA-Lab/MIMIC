module fake_ariane_2423_n_569 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_92, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_49, n_20, n_17, n_50, n_62, n_51, n_76, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_72, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_14, n_88, n_68, n_78, n_39, n_59, n_63, n_16, n_5, n_35, n_54, n_25, n_569);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_92;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_49;
input n_20;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_72;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_14;
input n_88;
input n_68;
input n_78;
input n_39;
input n_59;
input n_63;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_569;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_124;
wire n_119;
wire n_386;
wire n_307;
wire n_516;
wire n_332;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_205;
wire n_341;
wire n_109;
wire n_245;
wire n_421;
wire n_96;
wire n_549;
wire n_522;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_528;
wire n_387;
wire n_406;
wire n_117;
wire n_139;
wire n_524;
wire n_130;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_95;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_152;
wire n_405;
wire n_557;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_115;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_247;
wire n_567;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_108;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_511;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_104;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_565;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_448;
wire n_249;
wire n_534;
wire n_123;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_102;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_125;
wire n_407;
wire n_254;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_99;
wire n_544;
wire n_216;
wire n_540;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_509;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_98;
wire n_375;
wire n_113;
wire n_114;
wire n_324;
wire n_337;
wire n_437;
wire n_111;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_105;
wire n_494;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_118;
wire n_121;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_97;
wire n_408;
wire n_322;
wire n_251;
wire n_506;
wire n_558;
wire n_116;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_127;
wire n_531;

INVx1_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_30),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_6),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_9),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_20),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_39),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_5),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_34),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_37),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_62),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_70),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_74),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_24),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_L g123 ( 
.A(n_7),
.B(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_42),
.Y(n_130)
);

BUFx8_ASAP7_75t_SL g131 ( 
.A(n_31),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_22),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_17),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_75),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_50),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_21),
.Y(n_137)
);

NOR2xp67_ASAP7_75t_L g138 ( 
.A(n_16),
.B(n_8),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_73),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_2),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_36),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_15),
.B(n_35),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_47),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_38),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_3),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_66),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_49),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_19),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_11),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_18),
.Y(n_155)
);

BUFx8_ASAP7_75t_SL g156 ( 
.A(n_23),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_53),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_13),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_56),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_L g161 ( 
.A(n_10),
.B(n_33),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_67),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_1),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_11),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_2),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_71),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_28),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_57),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_46),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_4),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_55),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_44),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_86),
.Y(n_177)
);

BUFx2_ASAP7_75t_SL g178 ( 
.A(n_83),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_25),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_14),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_15),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_5),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_45),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_99),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_95),
.A2(n_0),
.B(n_4),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_112),
.B(n_0),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_103),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_98),
.B(n_80),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_97),
.B(n_6),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_8),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_100),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_102),
.A2(n_12),
.B(n_13),
.Y(n_198)
);

OAI21x1_ASAP7_75t_L g199 ( 
.A1(n_98),
.A2(n_32),
.B(n_43),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_14),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_99),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_64),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g206 ( 
.A1(n_108),
.A2(n_77),
.B(n_82),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_109),
.B(n_114),
.Y(n_213)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_99),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_109),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_112),
.B(n_153),
.Y(n_216)
);

AOI22x1_ASAP7_75t_SL g217 ( 
.A1(n_103),
.A2(n_154),
.B1(n_173),
.B2(n_140),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_114),
.B(n_135),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_112),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

CKINVDCx6p67_ASAP7_75t_R g222 ( 
.A(n_100),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_127),
.A2(n_150),
.B(n_183),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_110),
.A2(n_111),
.B1(n_173),
.B2(n_181),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_131),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_133),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_142),
.B(n_152),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_110),
.A2(n_111),
.B1(n_140),
.B2(n_181),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_147),
.B(n_184),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_155),
.A2(n_170),
.B(n_169),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_157),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g237 ( 
.A1(n_159),
.A2(n_160),
.B(n_165),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_168),
.A2(n_179),
.B(n_176),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_131),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_154),
.B(n_182),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_167),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_96),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_180),
.B(n_134),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g248 ( 
.A(n_178),
.B(n_156),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_101),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_104),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_107),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_123),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_113),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_115),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_118),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_156),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_119),
.B(n_120),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_121),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_130),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_256),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_191),
.Y(n_274)
);

OR2x6_ASAP7_75t_L g275 ( 
.A(n_189),
.B(n_214),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_242),
.B(n_136),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_226),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_226),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_192),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_137),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_233),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_162),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_192),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_177),
.C(n_139),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_205),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_225),
.Y(n_298)
);

CKINVDCx6p67_ASAP7_75t_R g299 ( 
.A(n_248),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_192),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_227),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_223),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_214),
.B(n_148),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_216),
.B(n_151),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_227),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_223),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_213),
.A2(n_218),
.B1(n_231),
.B2(n_239),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_255),
.B(n_171),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_225),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_203),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_205),
.Y(n_312)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_138),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_258),
.B(n_172),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

OAI221xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_231),
.B1(n_193),
.B2(n_195),
.C(n_200),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_231),
.B(n_235),
.C(n_205),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_263),
.B(n_287),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_297),
.A2(n_218),
.B1(n_213),
.B2(n_198),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_275),
.A2(n_248),
.B1(n_214),
.B2(n_220),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

NOR3xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_232),
.C(n_224),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_214),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_257),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_208),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_265),
.B(n_251),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_251),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_275),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_298),
.Y(n_334)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_305),
.B(n_259),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_259),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_301),
.A2(n_213),
.B1(n_218),
.B2(n_198),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_275),
.A2(n_196),
.B1(n_208),
.B2(n_241),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_253),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_264),
.B(n_253),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_271),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_306),
.B(n_248),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_293),
.A2(n_244),
.B1(n_220),
.B2(n_279),
.Y(n_344)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_271),
.Y(n_346)
);

OAI221xp5_ASAP7_75t_L g347 ( 
.A1(n_311),
.A2(n_252),
.B1(n_212),
.B2(n_219),
.C(n_236),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_313),
.B(n_185),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_185),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_253),
.Y(n_350)
);

O2A1O1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_278),
.A2(n_236),
.B(n_211),
.C(n_229),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_234),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_314),
.B(n_254),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_260),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_248),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_292),
.B(n_234),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_292),
.B(n_235),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_292),
.B(n_286),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_303),
.B(n_197),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_284),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_306),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_329),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_222),
.Y(n_365)
);

CKINVDCx10_ASAP7_75t_R g366 ( 
.A(n_323),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_317),
.A2(n_299),
.B1(n_161),
.B2(n_236),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_318),
.A2(n_303),
.B(n_206),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_327),
.A2(n_300),
.B(n_286),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_354),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_343),
.B(n_201),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_333),
.B(n_222),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_324),
.B(n_201),
.Y(n_375)
);

OAI21xp33_ASAP7_75t_L g376 ( 
.A1(n_331),
.A2(n_252),
.B(n_204),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_353),
.A2(n_206),
.B(n_199),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_261),
.Y(n_380)
);

AOI22x1_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_273),
.B1(n_260),
.B2(n_266),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_333),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_246),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_299),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_322),
.A2(n_204),
.B1(n_209),
.B2(n_221),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_339),
.B(n_348),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_272),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_221),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_355),
.A2(n_199),
.B(n_237),
.Y(n_391)
);

O2A1O1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_347),
.A2(n_336),
.B(n_351),
.C(n_344),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_332),
.A2(n_198),
.B1(n_188),
.B2(n_229),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_358),
.A2(n_238),
.B(n_294),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_349),
.B(n_246),
.Y(n_395)
);

BUFx12f_ASAP7_75t_L g396 ( 
.A(n_335),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_228),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_269),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_321),
.A2(n_188),
.B1(n_228),
.B2(n_290),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_243),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_321),
.A2(n_188),
.B1(n_295),
.B2(n_290),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_359),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_338),
.B(n_190),
.Y(n_405)
);

NAND2x1p5_ASAP7_75t_L g406 ( 
.A(n_338),
.B(n_207),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_318),
.A2(n_238),
.B(n_268),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_320),
.B(n_190),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_318),
.A2(n_270),
.B(n_277),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_329),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_320),
.B(n_202),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_320),
.A2(n_296),
.B(n_295),
.C(n_289),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_333),
.B(n_207),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_320),
.B(n_217),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_320),
.B(n_202),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_328),
.A2(n_266),
.B(n_267),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_329),
.B(n_207),
.Y(n_418)
);

NAND2x1p5_ASAP7_75t_L g419 ( 
.A(n_329),
.B(n_280),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_288),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_366),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_382),
.B(n_194),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_191),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_288),
.C(n_285),
.Y(n_424)
);

A2O1A1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_387),
.A2(n_283),
.B(n_281),
.C(n_280),
.Y(n_425)
);

AOI21x1_ASAP7_75t_SL g426 ( 
.A1(n_390),
.A2(n_192),
.B(n_262),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

BUFx12f_ASAP7_75t_L g428 ( 
.A(n_388),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_363),
.B(n_194),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_405),
.A2(n_281),
.B1(n_187),
.B2(n_186),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_191),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_385),
.A2(n_262),
.B(n_191),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g434 ( 
.A1(n_368),
.A2(n_394),
.B(n_391),
.Y(n_434)
);

OR2x6_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_186),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_377),
.A2(n_187),
.B(n_192),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_366),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_364),
.B(n_194),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_407),
.A2(n_194),
.B(n_217),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_409),
.A2(n_412),
.B(n_417),
.Y(n_440)
);

A2O1A1Ixp33_ASAP7_75t_L g441 ( 
.A1(n_392),
.A2(n_415),
.B(n_376),
.C(n_383),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_400),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_414),
.B(n_410),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_365),
.B(n_395),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_367),
.A2(n_406),
.B1(n_375),
.B2(n_384),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_413),
.B(n_389),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_386),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_419),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_380),
.A2(n_401),
.B1(n_378),
.B2(n_374),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_399),
.B(n_371),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_403),
.A2(n_381),
.B(n_369),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_398),
.B(n_372),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_404),
.B(n_397),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_379),
.A2(n_397),
.B(n_368),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_379),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_368),
.A2(n_394),
.B(n_391),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_364),
.B(n_408),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_362),
.B(n_320),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_362),
.B(n_408),
.Y(n_459)
);

AO32x2_ASAP7_75t_L g460 ( 
.A1(n_393),
.A2(n_401),
.A3(n_403),
.B1(n_367),
.B2(n_344),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_370),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_362),
.B(n_320),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_368),
.A2(n_394),
.B(n_391),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_373),
.Y(n_466)
);

INVx3_ASAP7_75t_SL g467 ( 
.A(n_388),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_364),
.B(n_408),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_362),
.B(n_343),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_368),
.A2(n_394),
.B(n_391),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_368),
.A2(n_394),
.B(n_391),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_362),
.B(n_320),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_362),
.B(n_343),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_368),
.A2(n_394),
.B(n_391),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_364),
.B(n_408),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_396),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_373),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_458),
.A2(n_464),
.B(n_472),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_459),
.A2(n_430),
.B1(n_439),
.B2(n_475),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_445),
.B(n_441),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_444),
.B(n_457),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_451),
.A2(n_436),
.B(n_426),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_443),
.Y(n_483)
);

BUFx2_ASAP7_75t_R g484 ( 
.A(n_467),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_476),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_476),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_434),
.A2(n_456),
.B(n_474),
.Y(n_487)
);

NAND3xp33_ASAP7_75t_SL g488 ( 
.A(n_468),
.B(n_445),
.C(n_442),
.Y(n_488)
);

OAI22xp33_ASAP7_75t_L g489 ( 
.A1(n_446),
.A2(n_448),
.B1(n_477),
.B2(n_466),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_465),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

AOI222xp33_ASAP7_75t_L g493 ( 
.A1(n_439),
.A2(n_430),
.B1(n_427),
.B2(n_437),
.C1(n_421),
.C2(n_447),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_473),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_471),
.B(n_454),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g496 ( 
.A1(n_435),
.A2(n_420),
.B1(n_450),
.B2(n_424),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

HB1xp67_ASAP7_75t_SL g498 ( 
.A(n_455),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

BUFx4_ASAP7_75t_SL g500 ( 
.A(n_435),
.Y(n_500)
);

CKINVDCx11_ASAP7_75t_R g501 ( 
.A(n_461),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_462),
.Y(n_502)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_424),
.A2(n_449),
.B(n_425),
.C(n_460),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_453),
.Y(n_504)
);

OAI222xp33_ASAP7_75t_L g505 ( 
.A1(n_452),
.A2(n_438),
.B1(n_422),
.B2(n_460),
.C1(n_431),
.C2(n_423),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_460),
.A2(n_440),
.B1(n_429),
.B2(n_433),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

AO31x2_ASAP7_75t_L g508 ( 
.A1(n_503),
.A2(n_506),
.A3(n_494),
.B(n_480),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_500),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_488),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_502),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_481),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_484),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_481),
.B(n_483),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_479),
.B(n_493),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_503),
.A2(n_505),
.B(n_496),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_483),
.B(n_489),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_504),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_495),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_498),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_499),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_491),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_507),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_501),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_487),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_482),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_508),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_523),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_510),
.B(n_518),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_517),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_525),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_519),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_518),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_527),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_518),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_526),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_533),
.B(n_509),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_529),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_521),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_541),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_537),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_542),
.B(n_532),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_541),
.B(n_530),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_529),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_532),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_510),
.B1(n_520),
.B2(n_530),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_545),
.B(n_538),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_544),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_545),
.A2(n_540),
.B1(n_538),
.B2(n_539),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_550),
.Y(n_553)
);

AOI211xp5_ASAP7_75t_L g554 ( 
.A1(n_552),
.A2(n_543),
.B(n_546),
.C(n_547),
.Y(n_554)
);

AOI21x1_ASAP7_75t_L g555 ( 
.A1(n_553),
.A2(n_551),
.B(n_534),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_514),
.Y(n_556)
);

NOR4xp25_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_509),
.C(n_522),
.D(n_549),
.Y(n_557)
);

NOR3x1_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_490),
.C(n_546),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_558),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_558),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_559),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_561),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_562),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_563),
.A2(n_560),
.B1(n_512),
.B2(n_485),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_564),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_554),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_486),
.B(n_492),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_486),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_501),
.B1(n_497),
.B2(n_492),
.Y(n_569)
);


endmodule