module fake_jpeg_24726_n_74 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_69;
wire n_40;
wire n_71;
wire n_35;
wire n_48;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_70;
wire n_66;

INVx11_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_9),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_37),
.B1(n_33),
.B2(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_46),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_1),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_37),
.C(n_38),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_39),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_41),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_42),
.C(n_4),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_47),
.B1(n_20),
.B2(n_5),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_3),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_22),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_62),
.B1(n_29),
.B2(n_10),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_65),
.Y(n_66)
);

AO221x1_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.C(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_17),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_65),
.Y(n_71)
);

AOI322xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_18),
.A3(n_19),
.B1(n_23),
.B2(n_24),
.C1(n_25),
.C2(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_27),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);


endmodule