module fake_netlist_5_1096_n_1723 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1723);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1723;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_52),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_40),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_17),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_43),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_12),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_15),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_9),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_16),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_1),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_3),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_77),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_10),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_1),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_27),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_99),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_49),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_21),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_95),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_39),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_136),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_23),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_16),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_23),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_22),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_62),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_102),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_87),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_40),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_80),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_19),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_42),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_22),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_34),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_2),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_18),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_60),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_4),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_83),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_88),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_5),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_124),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_0),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_70),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_79),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_90),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_36),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_82),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_53),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_71),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_10),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_74),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_73),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_85),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_138),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_118),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_50),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_122),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_107),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_120),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_45),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_42),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_17),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_29),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_129),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_116),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_8),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_6),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_114),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_54),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_109),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_8),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_111),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_119),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_39),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_51),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_44),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_91),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_100),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_47),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_68),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_24),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_66),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_3),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_46),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_55),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_86),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_45),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_34),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_106),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_47),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_20),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_49),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_56),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_21),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_94),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_140),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_92),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_97),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_30),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_28),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_61),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_67),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_105),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_103),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_15),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_108),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_26),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_75),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_151),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_115),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_137),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_117),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_2),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_153),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_24),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_69),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_27),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_104),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_142),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_93),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_11),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_96),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_41),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_64),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_4),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_84),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_33),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_72),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_229),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_191),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_155),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_185),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_185),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_185),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_185),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_185),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_195),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_234),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_195),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_161),
.B(n_5),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_195),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_195),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_267),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_193),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_195),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_199),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_283),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_241),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_199),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_178),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_299),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_297),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_205),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_207),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_208),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_233),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_213),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_214),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_199),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_161),
.B(n_6),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_216),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_217),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_278),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_163),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_233),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_178),
.B(n_7),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_219),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_163),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_276),
.B(n_9),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_199),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_223),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_276),
.B(n_12),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_227),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_199),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_278),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_176),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_176),
.B(n_13),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_228),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_240),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_248),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_251),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_253),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_164),
.B(n_13),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_256),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_258),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_261),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_197),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_262),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_197),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_266),
.B(n_212),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_166),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_260),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_220),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_220),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_260),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_268),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_166),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_170),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_268),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_294),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_170),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_311),
.B(n_212),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_172),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_226),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_316),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_226),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_172),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_319),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_323),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_383),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_351),
.Y(n_411)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_327),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_354),
.B(n_235),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_341),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_352),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_354),
.B(n_235),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_372),
.A2(n_175),
.B1(n_190),
.B2(n_238),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_369),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_371),
.A2(n_158),
.B(n_156),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_371),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_374),
.B(n_244),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_377),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_377),
.B(n_244),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_378),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_378),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_382),
.B(n_249),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_359),
.B(n_249),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

CKINVDCx8_ASAP7_75t_R g442 ( 
.A(n_324),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_321),
.B(n_293),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_342),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_365),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_331),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_331),
.B(n_294),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_328),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_332),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_309),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g452 ( 
.A(n_333),
.B(n_293),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_444),
.A2(n_288),
.B1(n_183),
.B2(n_173),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_442),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_451),
.B(n_329),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

NOR2x1p5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_308),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_448),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_446),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_398),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_451),
.B(n_329),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_442),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_451),
.B(n_345),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_384),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_324),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_325),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_442),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_413),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_394),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_390),
.B(n_179),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_413),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_430),
.Y(n_480)
);

BUFx4f_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_430),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_446),
.A2(n_236),
.B1(n_198),
.B2(n_162),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_430),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_387),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_390),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_335),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_449),
.B(n_345),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_417),
.A2(n_201),
.B1(n_187),
.B2(n_282),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_430),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_410),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_411),
.B(n_340),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_395),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_449),
.B(n_357),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_448),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_395),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_390),
.B(n_157),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_387),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_388),
.B(n_343),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_388),
.B(n_349),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_417),
.B(n_293),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_449),
.B(n_357),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_438),
.B(n_350),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_450),
.B(n_355),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_450),
.B(n_361),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_412),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_450),
.B(n_362),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_442),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_408),
.B(n_373),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_386),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_417),
.A2(n_422),
.B1(n_443),
.B2(n_440),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_386),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_402),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g527 ( 
.A(n_448),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_417),
.A2(n_284),
.B1(n_292),
.B2(n_304),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_401),
.B(n_363),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_438),
.B(n_347),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_398),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_403),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_386),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_410),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_411),
.B(n_364),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_403),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_403),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_411),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_389),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_385),
.Y(n_540)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_447),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_438),
.B(n_338),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_411),
.B(n_366),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_398),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_447),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_401),
.B(n_368),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_411),
.B(n_370),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_398),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_406),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_389),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_406),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_406),
.Y(n_553)
);

NAND2x1p5_ASAP7_75t_L g554 ( 
.A(n_443),
.B(n_160),
.Y(n_554)
);

BUFx8_ASAP7_75t_SL g555 ( 
.A(n_410),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_411),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_423),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_407),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_389),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_398),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_391),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_407),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_391),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_423),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_423),
.B(n_334),
.Y(n_566)
);

INVx4_ASAP7_75t_SL g567 ( 
.A(n_412),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_407),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_390),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_411),
.B(n_245),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_400),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_400),
.B(n_159),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_400),
.B(n_336),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_398),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_398),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_412),
.A2(n_344),
.B1(n_367),
.B2(n_337),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_400),
.B(n_339),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_411),
.B(n_353),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_422),
.B(n_293),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_422),
.B(n_360),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_443),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_412),
.B(n_379),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_398),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_422),
.B(n_278),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_440),
.B(n_165),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_443),
.B(n_293),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_411),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_391),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_412),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_412),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_443),
.A2(n_196),
.B1(n_307),
.B2(n_218),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_397),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_443),
.B(n_272),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_397),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_452),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_407),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_412),
.B(n_169),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_452),
.B(n_440),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_397),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_452),
.B(n_174),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_499),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_578),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_475),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_577),
.B(n_441),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_530),
.Y(n_606)
);

AOI221xp5_ASAP7_75t_L g607 ( 
.A1(n_558),
.A2(n_264),
.B1(n_300),
.B2(n_296),
.C(n_181),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_540),
.B(n_452),
.Y(n_608)
);

AND2x6_ASAP7_75t_SL g609 ( 
.A(n_489),
.B(n_177),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_481),
.B(n_254),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_464),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_524),
.B(n_452),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_480),
.A2(n_452),
.B1(n_440),
.B2(n_445),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_480),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_470),
.B(n_380),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_507),
.B(n_452),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_509),
.B(n_452),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_529),
.B(n_452),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_460),
.B(n_174),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_570),
.B(n_445),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_460),
.B(n_182),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_475),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_547),
.B(n_452),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_570),
.B(n_452),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_501),
.B(n_182),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_476),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_488),
.B(n_452),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_527),
.B(n_441),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_457),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_476),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_541),
.B(n_441),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_598),
.A2(n_385),
.B(n_432),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_473),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_461),
.B(n_441),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_482),
.A2(n_485),
.B1(n_517),
.B2(n_494),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_457),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_457),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_501),
.B(n_441),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_492),
.B(n_441),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_479),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_572),
.B(n_184),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_488),
.B(n_477),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_477),
.B(n_440),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_573),
.B(n_168),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_542),
.B(n_184),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_477),
.B(n_594),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_477),
.B(n_440),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_542),
.B(n_186),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_530),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_490),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_581),
.B(n_310),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_479),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_506),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_523),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_581),
.B(n_318),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_514),
.B(n_445),
.Y(n_658)
);

NAND2x1_ASAP7_75t_L g659 ( 
.A(n_514),
.B(n_392),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_523),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_525),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_514),
.B(n_445),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_500),
.B(n_186),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_583),
.B(n_230),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_514),
.B(n_399),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_545),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_512),
.B(n_230),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_585),
.B(n_231),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g669 ( 
.A1(n_565),
.A2(n_167),
.B1(n_300),
.B2(n_296),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_482),
.A2(n_385),
.B(n_432),
.C(n_435),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_514),
.B(n_399),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_574),
.B(n_188),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_533),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_574),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_515),
.B(n_231),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_514),
.B(n_399),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_586),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_585),
.B(n_265),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_485),
.B(n_404),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_494),
.B(n_404),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_517),
.B(n_404),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_513),
.B(n_265),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_499),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_522),
.B(n_405),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_522),
.B(n_405),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_513),
.B(n_275),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_518),
.B(n_192),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_533),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_573),
.B(n_168),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_497),
.A2(n_432),
.B(n_435),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_490),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_545),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_481),
.B(n_254),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_518),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_504),
.B(n_405),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_453),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_516),
.B(n_519),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_487),
.B(n_194),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_504),
.B(n_416),
.Y(n_699)
);

NOR2xp67_ASAP7_75t_L g700 ( 
.A(n_455),
.B(n_427),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_539),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_466),
.B(n_275),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_504),
.B(n_416),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_539),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_504),
.B(n_416),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_469),
.B(n_279),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_473),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_481),
.B(n_279),
.Y(n_708)
);

BUFx6f_ASAP7_75t_SL g709 ( 
.A(n_555),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_472),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_483),
.A2(n_254),
.B1(n_221),
.B2(n_224),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_487),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_518),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_551),
.B(n_419),
.Y(n_714)
);

AOI221xp5_ASAP7_75t_L g715 ( 
.A1(n_566),
.A2(n_181),
.B1(n_180),
.B2(n_171),
.C(n_306),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_551),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_458),
.B(n_505),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_560),
.Y(n_718)
);

NOR2x1p5_ASAP7_75t_L g719 ( 
.A(n_520),
.B(n_171),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_491),
.Y(n_720)
);

BUFx6f_ASAP7_75t_SL g721 ( 
.A(n_586),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_560),
.B(n_419),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_562),
.B(n_419),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_505),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_493),
.B(n_242),
.C(n_204),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_592),
.A2(n_320),
.B1(n_232),
.B2(n_225),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_562),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_564),
.B(n_421),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_491),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_456),
.B(n_280),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_564),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_491),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_599),
.A2(n_246),
.B(n_270),
.C(n_273),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_498),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_579),
.A2(n_301),
.B1(n_274),
.B2(n_281),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_596),
.B(n_254),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_590),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_463),
.A2(n_290),
.B1(n_305),
.B2(n_280),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_SL g739 ( 
.A(n_521),
.B(n_286),
.Y(n_739)
);

BUFx5_ASAP7_75t_L g740 ( 
.A(n_596),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_589),
.B(n_421),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_498),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_589),
.B(n_421),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_586),
.A2(n_290),
.B1(n_286),
.B2(n_287),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_593),
.B(n_424),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_593),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_596),
.B(n_287),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_595),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_595),
.B(n_424),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_596),
.B(n_289),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_600),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_582),
.B(n_289),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_469),
.B(n_233),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_498),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_502),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_582),
.B(n_295),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_600),
.B(n_424),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_502),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_571),
.B(n_392),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_502),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_465),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_495),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_473),
.B(n_392),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_503),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_465),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_473),
.B(n_392),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_590),
.B(n_291),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_473),
.B(n_392),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_554),
.B(n_295),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_473),
.B(n_392),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_467),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_582),
.B(n_254),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_602),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_603),
.B(n_534),
.Y(n_774)
);

AOI21x1_ASAP7_75t_L g775 ( 
.A1(n_659),
.A2(n_543),
.B(n_535),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_648),
.A2(n_548),
.B(n_590),
.Y(n_776)
);

NOR3xp33_ASAP7_75t_L g777 ( 
.A(n_615),
.B(n_601),
.C(n_305),
.Y(n_777)
);

INVx5_ASAP7_75t_L g778 ( 
.A(n_687),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_603),
.B(n_554),
.Y(n_779)
);

OAI21xp33_ASAP7_75t_L g780 ( 
.A1(n_739),
.A2(n_454),
.B(n_528),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_632),
.B(n_582),
.Y(n_781)
);

AO21x1_ASAP7_75t_L g782 ( 
.A1(n_735),
.A2(n_554),
.B(n_435),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_643),
.A2(n_591),
.B(n_538),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_644),
.A2(n_649),
.B(n_658),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_715),
.A2(n_586),
.B1(n_511),
.B2(n_580),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_662),
.A2(n_614),
.B(n_636),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_712),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_615),
.B(n_591),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_602),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_632),
.B(n_591),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_697),
.A2(n_459),
.B(n_584),
.C(n_575),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_614),
.A2(n_556),
.B(n_588),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_636),
.A2(n_556),
.B(n_588),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_627),
.A2(n_586),
.B1(n_511),
.B2(n_580),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_762),
.B(n_666),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_762),
.B(n_303),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_602),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_665),
.A2(n_569),
.B(n_588),
.Y(n_798)
);

NOR2x1_ASAP7_75t_R g799 ( 
.A(n_611),
.B(n_180),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_717),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_671),
.A2(n_569),
.B(n_588),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_635),
.B(n_511),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_724),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_607),
.B(n_303),
.C(n_257),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_635),
.B(n_511),
.Y(n_805)
);

BUFx4f_ASAP7_75t_L g806 ( 
.A(n_698),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_697),
.A2(n_459),
.B(n_584),
.C(n_575),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_676),
.A2(n_556),
.B(n_538),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_690),
.A2(n_597),
.B(n_503),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_628),
.B(n_511),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_694),
.A2(n_556),
.B(n_538),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_628),
.B(n_511),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_694),
.A2(n_569),
.B(n_538),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_713),
.A2(n_569),
.B(n_575),
.Y(n_814)
);

CKINVDCx10_ASAP7_75t_R g815 ( 
.A(n_709),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_612),
.A2(n_486),
.B1(n_584),
.B2(n_575),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_620),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_713),
.A2(n_561),
.B(n_531),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_639),
.B(n_511),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_740),
.B(n_567),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_737),
.A2(n_531),
.B(n_549),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_710),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_639),
.B(n_606),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_666),
.B(n_263),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_709),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_656),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_737),
.A2(n_531),
.B(n_549),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_606),
.B(n_580),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_692),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_759),
.A2(n_531),
.B(n_549),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_740),
.B(n_567),
.Y(n_831)
);

AOI21x1_ASAP7_75t_L g832 ( 
.A1(n_736),
.A2(n_484),
.B(n_478),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_651),
.B(n_580),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_696),
.B(n_189),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_660),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_651),
.A2(n_580),
.B1(n_587),
.B2(n_567),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_736),
.A2(n_484),
.B(n_478),
.Y(n_837)
);

OAI21xp33_ASAP7_75t_L g838 ( 
.A1(n_663),
.A2(n_269),
.B(n_263),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_653),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_608),
.A2(n_467),
.B(n_468),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_613),
.A2(n_633),
.B(n_624),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_657),
.Y(n_842)
);

BUFx4f_ASAP7_75t_L g843 ( 
.A(n_698),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_613),
.A2(n_550),
.B(n_468),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_692),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_602),
.B(n_486),
.Y(n_846)
);

OAI321xp33_ASAP7_75t_L g847 ( 
.A1(n_669),
.A2(n_433),
.A3(n_436),
.B1(n_437),
.B2(n_439),
.C(n_429),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_696),
.B(n_200),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_640),
.B(n_580),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_740),
.B(n_567),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_640),
.B(n_580),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_661),
.B(n_587),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_670),
.A2(n_536),
.B(n_471),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_630),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_677),
.B(n_427),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_772),
.A2(n_536),
.B(n_471),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_772),
.A2(n_537),
.B(n_474),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_673),
.B(n_587),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_695),
.A2(n_537),
.B(n_474),
.Y(n_859)
);

INVx8_ASAP7_75t_L g860 ( 
.A(n_677),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_655),
.Y(n_861)
);

INVx11_ASAP7_75t_L g862 ( 
.A(n_687),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_630),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_688),
.B(n_587),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_616),
.A2(n_597),
.B(n_546),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_699),
.A2(n_553),
.B(n_526),
.Y(n_866)
);

NOR3xp33_ASAP7_75t_L g867 ( 
.A(n_675),
.B(n_667),
.C(n_663),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_701),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_704),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_703),
.A2(n_553),
.B(n_526),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_716),
.B(n_718),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_727),
.B(n_587),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_731),
.B(n_746),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_674),
.B(n_202),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_677),
.B(n_427),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_700),
.B(n_567),
.Y(n_876)
);

AOI21xp33_ASAP7_75t_L g877 ( 
.A1(n_675),
.A2(n_252),
.B(n_203),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_667),
.A2(n_544),
.B(n_486),
.C(n_584),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_664),
.A2(n_532),
.B(n_550),
.C(n_552),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_753),
.B(n_655),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_642),
.B(n_206),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_748),
.B(n_587),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_706),
.B(n_269),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_705),
.A2(n_532),
.B(n_552),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_679),
.A2(n_597),
.B(n_503),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_617),
.A2(n_508),
.B(n_568),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_763),
.A2(n_486),
.B(n_496),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_751),
.B(n_587),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_604),
.B(n_496),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_680),
.A2(n_546),
.B(n_568),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_672),
.B(n_429),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_618),
.A2(n_557),
.B(n_568),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_622),
.B(n_496),
.Y(n_893)
);

AO21x1_ASAP7_75t_L g894 ( 
.A1(n_623),
.A2(n_563),
.B(n_559),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_L g895 ( 
.A(n_669),
.B(n_222),
.C(n_211),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_706),
.B(n_646),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_740),
.B(n_576),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_626),
.B(n_496),
.Y(n_898)
);

AO21x1_ASAP7_75t_L g899 ( 
.A1(n_610),
.A2(n_563),
.B(n_559),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_668),
.B(n_209),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_631),
.B(n_544),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_641),
.B(n_544),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_681),
.A2(n_546),
.B(n_563),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_634),
.A2(n_561),
.B(n_544),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_634),
.A2(n_561),
.B(n_549),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_654),
.B(n_561),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_629),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_630),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_678),
.B(n_215),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_740),
.B(n_605),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_689),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_769),
.B(n_508),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_707),
.A2(n_576),
.B(n_462),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_769),
.B(n_508),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_707),
.A2(n_576),
.B(n_462),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_630),
.A2(n_683),
.B1(n_685),
.B2(n_684),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_744),
.A2(n_510),
.B(n_559),
.C(n_557),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_610),
.A2(n_557),
.B(n_510),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_761),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_683),
.B(n_510),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_683),
.B(n_576),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_SL g922 ( 
.A(n_721),
.B(n_271),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_637),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_766),
.A2(n_576),
.B(n_462),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_683),
.B(n_393),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_687),
.Y(n_926)
);

NAND2x1p5_ASAP7_75t_L g927 ( 
.A(n_693),
.B(n_462),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_768),
.A2(n_462),
.B(n_409),
.Y(n_928)
);

NOR2x1_ASAP7_75t_L g929 ( 
.A(n_719),
.B(n_393),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_682),
.A2(n_439),
.B(n_437),
.C(n_436),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_771),
.B(n_393),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_638),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_730),
.B(n_237),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_693),
.A2(n_414),
.B(n_393),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_770),
.A2(n_414),
.B(n_393),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_647),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_645),
.A2(n_414),
.B(n_393),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_765),
.B(n_396),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_686),
.B(n_271),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_652),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_721),
.Y(n_941)
);

AO21x1_ASAP7_75t_L g942 ( 
.A1(n_714),
.A2(n_429),
.B(n_437),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_650),
.B(n_702),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_619),
.A2(n_439),
.B(n_433),
.C(n_436),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_722),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_726),
.B(n_433),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_691),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_720),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_698),
.B(n_277),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_621),
.B(n_243),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_625),
.B(n_247),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_723),
.A2(n_409),
.B(n_415),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_728),
.A2(n_757),
.B(n_745),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_729),
.B(n_462),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_741),
.B(n_425),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_672),
.B(n_306),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_732),
.A2(n_425),
.B(n_414),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_743),
.B(n_425),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_738),
.B(n_254),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_672),
.B(n_725),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_867),
.A2(n_733),
.B(n_756),
.C(n_752),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_774),
.B(n_609),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_877),
.A2(n_896),
.B(n_911),
.C(n_823),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_795),
.B(n_708),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_945),
.B(n_749),
.Y(n_965)
);

O2A1O1Ixp5_ASAP7_75t_L g966 ( 
.A1(n_942),
.A2(n_747),
.B(n_750),
.C(n_760),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_787),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_800),
.B(n_734),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_SL g969 ( 
.A1(n_788),
.A2(n_754),
.B(n_764),
.C(n_758),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_860),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_786),
.A2(n_711),
.B1(n_755),
.B2(n_742),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_786),
.B(n_767),
.Y(n_972)
);

NAND2xp33_ASAP7_75t_SL g973 ( 
.A(n_936),
.B(n_711),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_779),
.B(n_250),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_880),
.B(n_943),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_780),
.A2(n_255),
.B(n_259),
.C(n_302),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_SL g977 ( 
.A(n_838),
.B(n_277),
.C(n_285),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_826),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_860),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_845),
.B(n_285),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_871),
.A2(n_302),
.B1(n_431),
.B2(n_428),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_918),
.A2(n_425),
.B(n_396),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_829),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_861),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_803),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_804),
.A2(n_431),
.B(n_428),
.C(n_414),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_773),
.B(n_789),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_960),
.A2(n_767),
.B1(n_687),
.B2(n_254),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_796),
.B(n_767),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_950),
.A2(n_431),
.B(n_428),
.C(n_396),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_SL g991 ( 
.A(n_900),
.B(n_14),
.C(n_20),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_951),
.A2(n_431),
.B(n_428),
.C(n_396),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_910),
.A2(n_767),
.B(n_687),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_860),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_842),
.B(n_767),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_789),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_784),
.A2(n_396),
.B(n_425),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_824),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_891),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_784),
.A2(n_396),
.B(n_425),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_839),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_822),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_817),
.B(n_254),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_781),
.A2(n_414),
.B(n_420),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_940),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_777),
.A2(n_434),
.B1(n_426),
.B2(n_418),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_891),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_933),
.A2(n_420),
.B(n_415),
.C(n_409),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_868),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_835),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_883),
.B(n_434),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_869),
.B(n_873),
.Y(n_1012)
);

AO32x1_ASAP7_75t_L g1013 ( 
.A1(n_916),
.A2(n_409),
.A3(n_415),
.B1(n_420),
.B2(n_28),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_881),
.A2(n_420),
.B(n_415),
.C(n_434),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_919),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_789),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_940),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_785),
.A2(n_434),
.B1(n_426),
.B2(n_418),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_909),
.A2(n_434),
.B(n_426),
.C(n_418),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_790),
.B(n_434),
.Y(n_1020)
);

AO31x2_ASAP7_75t_L g1021 ( 
.A1(n_894),
.A2(n_14),
.A3(n_25),
.B(n_26),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_849),
.A2(n_434),
.B1(n_426),
.B2(n_418),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_949),
.B(n_434),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_956),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_773),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_R g1026 ( 
.A(n_825),
.B(n_63),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_941),
.B(n_65),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_907),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_841),
.A2(n_434),
.B(n_426),
.C(n_418),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_L g1030 ( 
.A(n_895),
.B(n_434),
.C(n_426),
.Y(n_1030)
);

NOR2xp67_ASAP7_75t_SL g1031 ( 
.A(n_778),
.B(n_426),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_806),
.B(n_426),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_851),
.A2(n_426),
.B1(n_418),
.B2(n_30),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_778),
.A2(n_418),
.B1(n_29),
.B2(n_31),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_897),
.A2(n_418),
.B(n_59),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_923),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_947),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_946),
.A2(n_25),
.B(n_31),
.C(n_32),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_939),
.B(n_834),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_799),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_947),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_953),
.B(n_418),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_953),
.A2(n_76),
.B(n_152),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_848),
.B(n_32),
.Y(n_1044)
);

OAI211xp5_ASAP7_75t_SL g1045 ( 
.A1(n_874),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_912),
.B(n_35),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_SL g1047 ( 
.A1(n_791),
.A2(n_81),
.B(n_147),
.C(n_139),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_941),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_929),
.A2(n_78),
.B1(n_134),
.B2(n_131),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_855),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_807),
.A2(n_959),
.B(n_930),
.C(n_847),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_878),
.A2(n_833),
.B(n_828),
.C(n_944),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_932),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_948),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_782),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_914),
.B(n_38),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_841),
.A2(n_43),
.B(n_44),
.C(n_46),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_863),
.B(n_48),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_815),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_SL g1060 ( 
.A1(n_809),
.A2(n_892),
.B(n_865),
.C(n_886),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_776),
.A2(n_110),
.B(n_57),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_810),
.A2(n_48),
.B(n_58),
.C(n_98),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_776),
.A2(n_121),
.B(n_126),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_806),
.B(n_128),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_921),
.A2(n_154),
.B(n_793),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_793),
.A2(n_920),
.B(n_805),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_931),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_855),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_843),
.A2(n_812),
.B1(n_922),
.B2(n_875),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_797),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_802),
.A2(n_831),
.B(n_820),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_843),
.B(n_778),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_778),
.A2(n_819),
.B1(n_875),
.B2(n_794),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_876),
.B(n_926),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_854),
.B(n_908),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_917),
.A2(n_816),
.B(n_889),
.C(n_906),
.Y(n_1076)
);

BUFx8_ASAP7_75t_L g1077 ( 
.A(n_926),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_876),
.B(n_926),
.Y(n_1078)
);

AO21x1_ASAP7_75t_L g1079 ( 
.A1(n_853),
.A2(n_859),
.B(n_866),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_783),
.A2(n_879),
.B(n_844),
.C(n_859),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_850),
.A2(n_783),
.B(n_808),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_908),
.B(n_925),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_SL g1083 ( 
.A(n_852),
.B(n_864),
.C(n_872),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_L g1084 ( 
.A(n_858),
.B(n_888),
.C(n_882),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_893),
.B(n_898),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_844),
.B(n_958),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_901),
.B(n_902),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_846),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_836),
.A2(n_899),
.B1(n_955),
.B2(n_938),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_798),
.A2(n_801),
.B(n_792),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_846),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_935),
.B(n_840),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_840),
.B(n_934),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_866),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_954),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_937),
.A2(n_957),
.B(n_853),
.C(n_856),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_856),
.A2(n_857),
.B(n_870),
.C(n_884),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_954),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_862),
.A2(n_927),
.B1(n_903),
.B2(n_890),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_870),
.B(n_884),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_R g1101 ( 
.A(n_832),
.B(n_837),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_952),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1039),
.B(n_903),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_967),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_964),
.A2(n_857),
.B(n_830),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_982),
.A2(n_887),
.B(n_775),
.Y(n_1106)
);

CKINVDCx6p67_ASAP7_75t_R g1107 ( 
.A(n_985),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_1002),
.Y(n_1108)
);

AOI221x1_ASAP7_75t_L g1109 ( 
.A1(n_1045),
.A2(n_952),
.B1(n_890),
.B2(n_885),
.C(n_928),
.Y(n_1109)
);

NOR2x1_ASAP7_75t_SL g1110 ( 
.A(n_1072),
.B(n_927),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1012),
.B(n_885),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_1001),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_984),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_1048),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1060),
.A2(n_1066),
.B(n_1086),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1086),
.A2(n_792),
.B(n_915),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_965),
.A2(n_827),
.B1(n_818),
.B2(n_821),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_961),
.A2(n_904),
.B(n_905),
.C(n_924),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_962),
.A2(n_814),
.B(n_913),
.C(n_811),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_SL g1120 ( 
.A1(n_1062),
.A2(n_813),
.B(n_1057),
.C(n_1032),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1090),
.A2(n_972),
.B(n_1081),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1024),
.A2(n_973),
.B1(n_998),
.B2(n_1044),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_963),
.A2(n_975),
.B(n_974),
.C(n_1038),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_976),
.A2(n_991),
.B(n_1034),
.C(n_1056),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1079),
.A2(n_1029),
.A3(n_1080),
.B(n_1019),
.Y(n_1125)
);

AND2x6_ASAP7_75t_L g1126 ( 
.A(n_1064),
.B(n_1098),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_984),
.B(n_983),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1024),
.A2(n_1007),
.B1(n_999),
.B2(n_1010),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1034),
.A2(n_1046),
.B(n_1033),
.C(n_977),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1033),
.A2(n_965),
.B(n_1058),
.C(n_1047),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_1074),
.A2(n_1078),
.B(n_972),
.C(n_1003),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_1059),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1096),
.A2(n_1085),
.B(n_1099),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1026),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_968),
.B(n_1009),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_983),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_L g1137 ( 
.A(n_970),
.B(n_979),
.Y(n_1137)
);

OA21x2_ASAP7_75t_L g1138 ( 
.A1(n_1042),
.A2(n_966),
.B(n_1094),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1069),
.A2(n_989),
.B1(n_1015),
.B2(n_995),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1099),
.A2(n_1092),
.B(n_1076),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1097),
.A2(n_1071),
.B(n_997),
.Y(n_1141)
);

OA21x2_ASAP7_75t_L g1142 ( 
.A1(n_1065),
.A2(n_1020),
.B(n_1100),
.Y(n_1142)
);

O2A1O1Ixp5_ASAP7_75t_SL g1143 ( 
.A1(n_1102),
.A2(n_981),
.B(n_1073),
.C(n_971),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1073),
.A2(n_969),
.B(n_1011),
.C(n_1067),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1087),
.B(n_1028),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1036),
.B(n_1053),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_SL g1147 ( 
.A1(n_1051),
.A2(n_992),
.B(n_990),
.C(n_1014),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_970),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1082),
.B(n_1023),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1000),
.A2(n_1004),
.B(n_1052),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1082),
.B(n_1037),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_980),
.B(n_1068),
.Y(n_1152)
);

OA21x2_ASAP7_75t_L g1153 ( 
.A1(n_1089),
.A2(n_1008),
.B(n_1093),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1030),
.A2(n_1043),
.B(n_1083),
.C(n_993),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_994),
.B(n_970),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1005),
.B(n_1017),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1054),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_971),
.A2(n_1063),
.B(n_1061),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_1077),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1050),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_988),
.A2(n_1055),
.B(n_1084),
.C(n_1027),
.Y(n_1161)
);

NOR2x1_ASAP7_75t_L g1162 ( 
.A(n_994),
.B(n_1025),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1050),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_986),
.A2(n_1035),
.B(n_1049),
.C(n_1075),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1013),
.A2(n_1031),
.B(n_1018),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1013),
.A2(n_1018),
.B(n_1088),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1040),
.A2(n_1050),
.B1(n_1041),
.B2(n_981),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_979),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1070),
.B(n_996),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1022),
.A2(n_1013),
.A3(n_1101),
.B(n_1021),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_987),
.A2(n_1025),
.B(n_1098),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1006),
.A2(n_987),
.B(n_996),
.Y(n_1172)
);

CKINVDCx11_ASAP7_75t_R g1173 ( 
.A(n_979),
.Y(n_1173)
);

OAI22x1_ASAP7_75t_L g1174 ( 
.A1(n_1077),
.A2(n_1021),
.B1(n_1091),
.B2(n_1095),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1016),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1016),
.A2(n_867),
.B(n_697),
.C(n_964),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_994),
.B(n_970),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_985),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1039),
.B(n_896),
.Y(n_1179)
);

NAND2x1_ASAP7_75t_L g1180 ( 
.A(n_1025),
.B(n_773),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1060),
.A2(n_910),
.B(n_784),
.Y(n_1181)
);

AO21x1_ASAP7_75t_L g1182 ( 
.A1(n_1033),
.A2(n_867),
.B(n_961),
.Y(n_1182)
);

BUFx10_ASAP7_75t_L g1183 ( 
.A(n_1059),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_964),
.A2(n_867),
.B(n_781),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_970),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1060),
.A2(n_910),
.B(n_784),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_SL g1187 ( 
.A1(n_989),
.A2(n_910),
.B(n_781),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_970),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_970),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1079),
.A2(n_1029),
.A3(n_942),
.B(n_1080),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1060),
.A2(n_910),
.B(n_784),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1039),
.B(n_896),
.Y(n_1192)
);

AO21x1_ASAP7_75t_L g1193 ( 
.A1(n_1033),
.A2(n_867),
.B(n_961),
.Y(n_1193)
);

INVx3_ASAP7_75t_SL g1194 ( 
.A(n_1059),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_962),
.A2(n_867),
.B(n_603),
.C(n_877),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_962),
.B(n_603),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1079),
.A2(n_1029),
.A3(n_942),
.B(n_1080),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_982),
.A2(n_887),
.B(n_1081),
.Y(n_1198)
);

INVx5_ASAP7_75t_L g1199 ( 
.A(n_1016),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_1029),
.A2(n_972),
.B(n_1080),
.Y(n_1200)
);

AO21x2_ASAP7_75t_L g1201 ( 
.A1(n_1029),
.A2(n_1060),
.B(n_1080),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1039),
.B(n_896),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_978),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_984),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1039),
.B(n_867),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_970),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_982),
.A2(n_887),
.B(n_1081),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1079),
.A2(n_1029),
.A3(n_942),
.B(n_1080),
.Y(n_1208)
);

AO21x1_ASAP7_75t_L g1209 ( 
.A1(n_1033),
.A2(n_867),
.B(n_961),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1048),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_994),
.B(n_970),
.Y(n_1211)
);

NAND3xp33_ASAP7_75t_L g1212 ( 
.A(n_962),
.B(n_867),
.C(n_603),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_994),
.B(n_970),
.Y(n_1213)
);

AOI31xp67_ASAP7_75t_L g1214 ( 
.A1(n_972),
.A2(n_1042),
.A3(n_1089),
.B(n_1086),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_1062),
.A2(n_1057),
.B(n_807),
.C(n_791),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_973),
.A2(n_867),
.B1(n_804),
.B2(n_566),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_984),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1060),
.A2(n_910),
.B(n_784),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_SL g1219 ( 
.A(n_970),
.B(n_442),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1060),
.A2(n_910),
.B(n_784),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_964),
.A2(n_867),
.B1(n_788),
.B2(n_603),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_964),
.A2(n_867),
.B(n_781),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1060),
.A2(n_910),
.B(n_784),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1079),
.A2(n_1029),
.A3(n_942),
.B(n_1080),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1024),
.B(n_1001),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_962),
.B(n_867),
.C(n_603),
.Y(n_1226)
);

OR2x6_ASAP7_75t_L g1227 ( 
.A(n_1002),
.B(n_860),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_SL g1228 ( 
.A1(n_989),
.A2(n_910),
.B(n_781),
.Y(n_1228)
);

NOR2x1_ASAP7_75t_SL g1229 ( 
.A(n_1099),
.B(n_1102),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_964),
.A2(n_867),
.B1(n_788),
.B2(n_603),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1039),
.B(n_896),
.Y(n_1231)
);

BUFx8_ASAP7_75t_L g1232 ( 
.A(n_1002),
.Y(n_1232)
);

NAND3xp33_ASAP7_75t_L g1233 ( 
.A(n_962),
.B(n_867),
.C(n_603),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1060),
.A2(n_910),
.B(n_784),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1024),
.B(n_1001),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_970),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_SL g1237 ( 
.A1(n_963),
.A2(n_715),
.B1(n_838),
.B2(n_669),
.C(n_607),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_962),
.A2(n_867),
.B1(n_615),
.B2(n_839),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_982),
.A2(n_887),
.B(n_1081),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_964),
.A2(n_867),
.B(n_697),
.C(n_961),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_SL g1241 ( 
.A1(n_963),
.A2(n_715),
.B1(n_838),
.B2(n_669),
.C(n_607),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1210),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1238),
.A2(n_1221),
.B1(n_1230),
.B2(n_1122),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1196),
.A2(n_1212),
.B1(n_1226),
.B2(n_1233),
.Y(n_1244)
);

CKINVDCx16_ASAP7_75t_R g1245 ( 
.A(n_1132),
.Y(n_1245)
);

CKINVDCx11_ASAP7_75t_R g1246 ( 
.A(n_1194),
.Y(n_1246)
);

BUFx12f_ASAP7_75t_L g1247 ( 
.A(n_1173),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1216),
.A2(n_1193),
.B1(n_1209),
.B2(n_1182),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1232),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1232),
.Y(n_1250)
);

BUFx2_ASAP7_75t_SL g1251 ( 
.A(n_1159),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1203),
.Y(n_1252)
);

CKINVDCx6p67_ASAP7_75t_R g1253 ( 
.A(n_1183),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1217),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1184),
.A2(n_1222),
.B1(n_1205),
.B2(n_1179),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1192),
.A2(n_1231),
.B1(n_1202),
.B2(n_1133),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1240),
.A2(n_1135),
.B1(n_1176),
.B2(n_1195),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1108),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1183),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1140),
.A2(n_1103),
.B1(n_1139),
.B2(n_1113),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1229),
.A2(n_1126),
.B1(n_1152),
.B2(n_1112),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1204),
.A2(n_1136),
.B1(n_1111),
.B2(n_1235),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1138),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1225),
.A2(n_1145),
.B1(n_1128),
.B2(n_1127),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1104),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1178),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1146),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1107),
.Y(n_1268)
);

INVx8_ASAP7_75t_L g1269 ( 
.A(n_1199),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1138),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1241),
.A2(n_1237),
.B1(n_1153),
.B2(n_1158),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1148),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1153),
.A2(n_1201),
.B1(n_1105),
.B2(n_1200),
.Y(n_1273)
);

BUFx8_ASAP7_75t_L g1274 ( 
.A(n_1148),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1157),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1156),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1200),
.A2(n_1126),
.B1(n_1115),
.B2(n_1219),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1126),
.A2(n_1167),
.B1(n_1166),
.B2(n_1165),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1126),
.A2(n_1149),
.B1(n_1114),
.B2(n_1151),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1280)
);

CKINVDCx6p67_ASAP7_75t_R g1281 ( 
.A(n_1168),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1169),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1161),
.A2(n_1227),
.B1(n_1129),
.B2(n_1164),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1175),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1160),
.B(n_1163),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1227),
.A2(n_1154),
.B1(n_1134),
.B2(n_1130),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1199),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1174),
.A2(n_1142),
.B1(n_1117),
.B2(n_1234),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1177),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_SL g1290 ( 
.A1(n_1211),
.A2(n_1185),
.B1(n_1236),
.B2(n_1188),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1229),
.A2(n_1110),
.B1(n_1172),
.B2(n_1137),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1185),
.A2(n_1188),
.B1(n_1236),
.B2(n_1189),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1188),
.B(n_1236),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1131),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1190),
.Y(n_1295)
);

INVx3_ASAP7_75t_SL g1296 ( 
.A(n_1206),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1187),
.A2(n_1228),
.B1(n_1162),
.B2(n_1213),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1190),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1206),
.A2(n_1142),
.B1(n_1150),
.B2(n_1143),
.Y(n_1299)
);

CKINVDCx11_ASAP7_75t_R g1300 ( 
.A(n_1206),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1197),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1181),
.A2(n_1186),
.B1(n_1223),
.B2(n_1191),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1218),
.A2(n_1220),
.B1(n_1121),
.B2(n_1141),
.Y(n_1303)
);

CKINVDCx6p67_ASAP7_75t_R g1304 ( 
.A(n_1171),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1116),
.A2(n_1180),
.B1(n_1207),
.B2(n_1198),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1208),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1239),
.A2(n_1106),
.B1(n_1215),
.B2(n_1120),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1119),
.A2(n_1118),
.B(n_1144),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1208),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1214),
.A2(n_1147),
.B1(n_1109),
.B2(n_1224),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1224),
.A2(n_867),
.B1(n_1216),
.B2(n_1193),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1224),
.Y(n_1312)
);

BUFx2_ASAP7_75t_SL g1313 ( 
.A(n_1125),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1125),
.B(n_1170),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1170),
.A2(n_867),
.B1(n_1216),
.B2(n_1193),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1170),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1104),
.Y(n_1317)
);

INVx6_ASAP7_75t_L g1318 ( 
.A(n_1232),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1132),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1232),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1179),
.B(n_1039),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1232),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1199),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1196),
.A2(n_739),
.B1(n_962),
.B2(n_521),
.Y(n_1324)
);

BUFx4f_ASAP7_75t_SL g1325 ( 
.A(n_1132),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1216),
.A2(n_867),
.B1(n_1193),
.B2(n_1182),
.Y(n_1326)
);

INVx6_ASAP7_75t_L g1327 ( 
.A(n_1232),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1216),
.A2(n_867),
.B1(n_1193),
.B2(n_1182),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1232),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1196),
.A2(n_739),
.B1(n_962),
.B2(n_521),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1196),
.A2(n_739),
.B1(n_962),
.B2(n_521),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1194),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1232),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1194),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1216),
.A2(n_867),
.B1(n_1193),
.B2(n_1182),
.Y(n_1335)
);

INVx4_ASAP7_75t_L g1336 ( 
.A(n_1199),
.Y(n_1336)
);

INVxp67_ASAP7_75t_SL g1337 ( 
.A(n_1113),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1216),
.A2(n_867),
.B1(n_1193),
.B2(n_1182),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1196),
.A2(n_1216),
.B1(n_1238),
.B2(n_603),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1132),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1232),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1194),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1196),
.A2(n_1216),
.B1(n_1238),
.B2(n_603),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1199),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_1155),
.Y(n_1345)
);

INVx8_ASAP7_75t_L g1346 ( 
.A(n_1199),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1199),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1216),
.A2(n_867),
.B1(n_1193),
.B2(n_1182),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1210),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1295),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1263),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1301),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1270),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1309),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1254),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1321),
.B(n_1339),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1274),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1315),
.B(n_1311),
.Y(n_1358)
);

AND2x2_ASAP7_75t_SL g1359 ( 
.A(n_1248),
.B(n_1326),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1308),
.A2(n_1314),
.B(n_1294),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1306),
.B(n_1280),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1343),
.A2(n_1330),
.B1(n_1331),
.B2(n_1324),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_R g1363 ( 
.A(n_1247),
.B(n_1246),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1265),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1317),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1316),
.B(n_1298),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1274),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1255),
.B(n_1267),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1252),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1323),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1310),
.A2(n_1273),
.B(n_1315),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1311),
.B(n_1248),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1275),
.Y(n_1373)
);

BUFx2_ASAP7_75t_R g1374 ( 
.A(n_1251),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1312),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1304),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1283),
.A2(n_1257),
.B(n_1243),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1242),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1337),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1313),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1326),
.B(n_1328),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1243),
.A2(n_1338),
.B1(n_1348),
.B2(n_1335),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1244),
.A2(n_1286),
.B1(n_1335),
.B2(n_1328),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1262),
.B(n_1260),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1338),
.A2(n_1348),
.B(n_1256),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1262),
.B(n_1260),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1282),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1276),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1271),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1349),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1271),
.B(n_1256),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1305),
.A2(n_1307),
.B(n_1288),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1273),
.Y(n_1393)
);

INVx11_ASAP7_75t_L g1394 ( 
.A(n_1247),
.Y(n_1394)
);

CKINVDCx6p67_ASAP7_75t_R g1395 ( 
.A(n_1332),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1310),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1258),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1278),
.B(n_1288),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1278),
.B(n_1284),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1297),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1258),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1279),
.A2(n_1261),
.B1(n_1264),
.B2(n_1327),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1277),
.B(n_1264),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1272),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1302),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1303),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1299),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1307),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1291),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1277),
.A2(n_1346),
.B(n_1269),
.C(n_1345),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1305),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1345),
.A2(n_1293),
.B(n_1285),
.Y(n_1412)
);

BUFx2_ASAP7_75t_R g1413 ( 
.A(n_1322),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1290),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1383),
.B(n_1289),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1385),
.A2(n_1292),
.B(n_1287),
.Y(n_1416)
);

NAND2xp33_ASAP7_75t_R g1417 ( 
.A(n_1376),
.B(n_1259),
.Y(n_1417)
);

AOI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1382),
.A2(n_1362),
.B1(n_1381),
.B2(n_1377),
.C(n_1356),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1403),
.B(n_1266),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1379),
.B(n_1296),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1412),
.B(n_1296),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1368),
.B(n_1268),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1395),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1387),
.B(n_1250),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1392),
.A2(n_1336),
.B(n_1346),
.Y(n_1425)
);

AOI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1381),
.A2(n_1320),
.B1(n_1329),
.B2(n_1341),
.C(n_1322),
.Y(n_1426)
);

INVxp33_ASAP7_75t_SL g1427 ( 
.A(n_1363),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1412),
.B(n_1336),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1393),
.B(n_1327),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1377),
.A2(n_1253),
.B(n_1300),
.C(n_1281),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1359),
.A2(n_1319),
.B(n_1340),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1377),
.A2(n_1245),
.B1(n_1346),
.B2(n_1269),
.C(n_1347),
.Y(n_1432)
);

NOR2x1_ASAP7_75t_SL g1433 ( 
.A(n_1360),
.B(n_1347),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1369),
.B(n_1347),
.Y(n_1434)
);

OA21x2_ASAP7_75t_L g1435 ( 
.A1(n_1392),
.A2(n_1269),
.B(n_1344),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1355),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1375),
.B(n_1300),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1409),
.A2(n_1249),
.B(n_1318),
.C(n_1333),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1373),
.B(n_1318),
.Y(n_1439)
);

NOR2x1_ASAP7_75t_L g1440 ( 
.A(n_1376),
.B(n_1325),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1376),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1409),
.A2(n_1333),
.B(n_1272),
.C(n_1334),
.Y(n_1442)
);

BUFx4f_ASAP7_75t_SL g1443 ( 
.A(n_1395),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1397),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1405),
.B(n_1342),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1405),
.B(n_1325),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1359),
.A2(n_1372),
.B(n_1358),
.C(n_1398),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1359),
.B(n_1400),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1400),
.B(n_1399),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1410),
.A2(n_1384),
.B(n_1386),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1384),
.B(n_1386),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1350),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1399),
.B(n_1391),
.Y(n_1454)
);

NOR2x1_ASAP7_75t_SL g1455 ( 
.A(n_1360),
.B(n_1398),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1371),
.B(n_1358),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1371),
.B(n_1391),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1397),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1371),
.B(n_1411),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1401),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1454),
.B(n_1360),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1457),
.B(n_1456),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1455),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1418),
.A2(n_1372),
.B1(n_1402),
.B2(n_1406),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1420),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1459),
.B(n_1411),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1457),
.B(n_1351),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1453),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1459),
.B(n_1353),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1428),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1448),
.B(n_1406),
.C(n_1407),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1428),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1448),
.A2(n_1364),
.B1(n_1407),
.B2(n_1389),
.C(n_1365),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_1433),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1428),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1449),
.A2(n_1415),
.B1(n_1431),
.B2(n_1452),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1441),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1447),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1421),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1435),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1435),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1435),
.B(n_1352),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1450),
.B(n_1366),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1458),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1425),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1434),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1466),
.B(n_1396),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1461),
.B(n_1396),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1482),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1462),
.B(n_1361),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1468),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1470),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1474),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1462),
.B(n_1361),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1471),
.A2(n_1449),
.B1(n_1451),
.B2(n_1430),
.C(n_1416),
.Y(n_1495)
);

NOR2x1_ASAP7_75t_L g1496 ( 
.A(n_1484),
.B(n_1458),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1462),
.B(n_1429),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1481),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1470),
.B(n_1429),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1475),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1461),
.B(n_1419),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1470),
.B(n_1467),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1480),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1468),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1480),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1474),
.Y(n_1506)
);

AO21x1_ASAP7_75t_SL g1507 ( 
.A1(n_1481),
.A2(n_1380),
.B(n_1408),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1466),
.B(n_1408),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1477),
.Y(n_1509)
);

INVx5_ASAP7_75t_L g1510 ( 
.A(n_1480),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1467),
.B(n_1371),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1466),
.B(n_1354),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1469),
.B(n_1354),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1508),
.B(n_1483),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1513),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1502),
.B(n_1492),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1513),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1508),
.B(n_1483),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1502),
.B(n_1492),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1495),
.A2(n_1471),
.B1(n_1464),
.B2(n_1473),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1513),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1492),
.B(n_1475),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1496),
.B(n_1477),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1503),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1492),
.B(n_1475),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1511),
.B(n_1479),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1509),
.B(n_1472),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1472),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1508),
.B(n_1483),
.Y(n_1530)
);

NAND2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1496),
.B(n_1477),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1511),
.B(n_1472),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1488),
.B(n_1478),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1509),
.B(n_1463),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1488),
.B(n_1478),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1514),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1497),
.B(n_1465),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1514),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1497),
.B(n_1465),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1503),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1514),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1504),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1491),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1491),
.B(n_1478),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1517),
.B(n_1499),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1547),
.Y(n_1549)
);

NOR2x1_ASAP7_75t_L g1550 ( 
.A(n_1547),
.B(n_1423),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1517),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1515),
.B(n_1501),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1544),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1544),
.Y(n_1554)
);

NAND4xp25_ASAP7_75t_SL g1555 ( 
.A(n_1521),
.B(n_1495),
.C(n_1476),
.D(n_1473),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1521),
.B(n_1501),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1532),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1537),
.B(n_1490),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1534),
.B(n_1509),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1515),
.B(n_1487),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1519),
.B(n_1487),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1543),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_L g1563 ( 
.A(n_1528),
.B(n_1493),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1537),
.B(n_1490),
.Y(n_1564)
);

NAND2xp33_ASAP7_75t_SL g1565 ( 
.A(n_1540),
.B(n_1417),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1519),
.B(n_1487),
.Y(n_1566)
);

NAND4xp25_ASAP7_75t_L g1567 ( 
.A(n_1520),
.B(n_1476),
.C(n_1464),
.D(n_1426),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1499),
.Y(n_1568)
);

AO21x1_ASAP7_75t_L g1569 ( 
.A1(n_1524),
.A2(n_1498),
.B(n_1509),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1540),
.B(n_1490),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1534),
.B(n_1493),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1543),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1545),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1530),
.B(n_1494),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1494),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1533),
.B(n_1494),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1523),
.B(n_1499),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1532),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1523),
.B(n_1493),
.Y(n_1579)
);

NOR2x1_ASAP7_75t_L g1580 ( 
.A(n_1534),
.B(n_1423),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1533),
.B(n_1486),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1545),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1516),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1523),
.B(n_1506),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1535),
.B(n_1486),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1524),
.B(n_1438),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1516),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1518),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1526),
.B(n_1506),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1555),
.A2(n_1432),
.B1(n_1534),
.B2(n_1528),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1580),
.B(n_1550),
.Y(n_1591)
);

AOI21xp33_ASAP7_75t_L g1592 ( 
.A1(n_1556),
.A2(n_1417),
.B(n_1445),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1518),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1574),
.B(n_1536),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1562),
.Y(n_1595)
);

OAI21xp33_ASAP7_75t_L g1596 ( 
.A1(n_1567),
.A2(n_1535),
.B(n_1422),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1554),
.B(n_1549),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1548),
.B(n_1529),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1548),
.B(n_1529),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1568),
.B(n_1527),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1562),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1572),
.B(n_1522),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1571),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1551),
.B(n_1528),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1551),
.B(n_1559),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1575),
.B(n_1536),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1559),
.B(n_1568),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1582),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1563),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1588),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1588),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1552),
.B(n_1538),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1565),
.A2(n_1446),
.B1(n_1445),
.B2(n_1528),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1565),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1571),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1583),
.B(n_1522),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1587),
.B(n_1538),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1559),
.B(n_1527),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1560),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1558),
.B(n_1427),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1561),
.Y(n_1622)
);

NAND4xp25_ASAP7_75t_L g1623 ( 
.A(n_1579),
.B(n_1442),
.C(n_1415),
.D(n_1589),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1542),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1591),
.A2(n_1586),
.B(n_1569),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1611),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1612),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1596),
.B(n_1577),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1591),
.B(n_1577),
.Y(n_1629)
);

OAI211xp5_ASAP7_75t_L g1630 ( 
.A1(n_1615),
.A2(n_1589),
.B(n_1579),
.C(n_1584),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1605),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1621),
.B(n_1597),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1605),
.Y(n_1633)
);

OAI21xp33_ASAP7_75t_L g1634 ( 
.A1(n_1615),
.A2(n_1586),
.B(n_1584),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1606),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1620),
.B(n_1566),
.Y(n_1636)
);

AOI21xp33_ASAP7_75t_L g1637 ( 
.A1(n_1614),
.A2(n_1586),
.B(n_1571),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1604),
.B(n_1564),
.Y(n_1638)
);

OAI21xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1610),
.A2(n_1570),
.B(n_1557),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1616),
.B(n_1622),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1606),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1595),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1590),
.A2(n_1524),
.B1(n_1531),
.B2(n_1578),
.Y(n_1643)
);

AOI332xp33_ASAP7_75t_L g1644 ( 
.A1(n_1601),
.A2(n_1578),
.A3(n_1557),
.B1(n_1542),
.B2(n_1539),
.B3(n_1541),
.C1(n_1525),
.C2(n_1489),
.Y(n_1644)
);

NOR2x1_ASAP7_75t_SL g1645 ( 
.A(n_1603),
.B(n_1507),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1623),
.A2(n_1524),
.B1(n_1531),
.B2(n_1506),
.Y(n_1647)
);

AOI21xp33_ASAP7_75t_L g1648 ( 
.A1(n_1593),
.A2(n_1463),
.B(n_1446),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1610),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1630),
.A2(n_1592),
.B1(n_1593),
.B2(n_1608),
.C(n_1618),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1626),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1632),
.A2(n_1592),
.B1(n_1608),
.B2(n_1619),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1635),
.B(n_1600),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1625),
.B(n_1427),
.Y(n_1654)
);

OAI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1628),
.A2(n_1531),
.B1(n_1485),
.B2(n_1598),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1635),
.B(n_1599),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1626),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1629),
.B(n_1594),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1629),
.A2(n_1531),
.B1(n_1607),
.B2(n_1613),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_SL g1660 ( 
.A1(n_1634),
.A2(n_1624),
.B1(n_1618),
.B2(n_1617),
.C(n_1602),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1627),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1627),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1636),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1649),
.Y(n_1664)
);

AOI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1637),
.A2(n_1617),
.B(n_1602),
.C(n_1624),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1647),
.A2(n_1643),
.B(n_1640),
.Y(n_1666)
);

INVxp67_ASAP7_75t_SL g1667 ( 
.A(n_1649),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1641),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1654),
.B(n_1443),
.Y(n_1669)
);

NOR2x1_ASAP7_75t_L g1670 ( 
.A(n_1664),
.B(n_1641),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1663),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1654),
.B(n_1668),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1658),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1667),
.Y(n_1674)
);

AOI222xp33_ASAP7_75t_L g1675 ( 
.A1(n_1650),
.A2(n_1642),
.B1(n_1639),
.B2(n_1646),
.C1(n_1638),
.C2(n_1631),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1653),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1651),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1657),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1661),
.Y(n_1679)
);

AOI221x1_ASAP7_75t_L g1680 ( 
.A1(n_1674),
.A2(n_1662),
.B1(n_1659),
.B2(n_1656),
.C(n_1631),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1673),
.B(n_1633),
.Y(n_1681)
);

NOR3x1_ASAP7_75t_L g1682 ( 
.A(n_1676),
.B(n_1666),
.C(n_1636),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1669),
.B(n_1660),
.Y(n_1683)
);

AOI211xp5_ASAP7_75t_L g1684 ( 
.A1(n_1672),
.A2(n_1655),
.B(n_1665),
.C(n_1633),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1670),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1678),
.Y(n_1686)
);

NOR3xp33_ASAP7_75t_L g1687 ( 
.A(n_1673),
.B(n_1655),
.C(n_1648),
.Y(n_1687)
);

OAI211xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1675),
.A2(n_1652),
.B(n_1390),
.C(n_1378),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1671),
.B(n_1652),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1684),
.B(n_1677),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1688),
.A2(n_1678),
.B1(n_1679),
.B2(n_1440),
.C(n_1644),
.Y(n_1691)
);

AOI222xp33_ASAP7_75t_L g1692 ( 
.A1(n_1685),
.A2(n_1645),
.B1(n_1498),
.B2(n_1436),
.C1(n_1485),
.C2(n_1424),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1683),
.A2(n_1444),
.B1(n_1460),
.B2(n_1526),
.C(n_1546),
.Y(n_1693)
);

A2O1A1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1687),
.A2(n_1357),
.B(n_1645),
.C(n_1526),
.Y(n_1694)
);

NOR4xp25_ASAP7_75t_L g1695 ( 
.A(n_1689),
.B(n_1546),
.C(n_1541),
.D(n_1539),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1691),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1694),
.A2(n_1681),
.B1(n_1686),
.B2(n_1682),
.C(n_1692),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1690),
.A2(n_1680),
.B(n_1357),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_L g1699 ( 
.A(n_1693),
.B(n_1394),
.C(n_1404),
.Y(n_1699)
);

OAI222xp33_ASAP7_75t_L g1700 ( 
.A1(n_1695),
.A2(n_1441),
.B1(n_1510),
.B2(n_1585),
.C1(n_1581),
.C2(n_1500),
.Y(n_1700)
);

NOR4xp25_ASAP7_75t_L g1701 ( 
.A(n_1690),
.B(n_1394),
.C(n_1525),
.D(n_1539),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1692),
.B(n_1510),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1702),
.Y(n_1703)
);

INVxp33_ASAP7_75t_L g1704 ( 
.A(n_1698),
.Y(n_1704)
);

AO22x2_ASAP7_75t_L g1705 ( 
.A1(n_1699),
.A2(n_1525),
.B1(n_1541),
.B2(n_1532),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1696),
.Y(n_1706)
);

XNOR2xp5_ASAP7_75t_L g1707 ( 
.A(n_1701),
.B(n_1697),
.Y(n_1707)
);

NAND3xp33_ASAP7_75t_L g1708 ( 
.A(n_1707),
.B(n_1700),
.C(n_1404),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1706),
.Y(n_1709)
);

NAND2x1p5_ASAP7_75t_L g1710 ( 
.A(n_1703),
.B(n_1401),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1709),
.B(n_1704),
.Y(n_1711)
);

OAI22x1_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1708),
.B1(n_1710),
.B2(n_1705),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1705),
.B1(n_1367),
.B2(n_1510),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1712),
.A2(n_1413),
.B(n_1437),
.Y(n_1714)
);

OAI22x1_ASAP7_75t_L g1715 ( 
.A1(n_1714),
.A2(n_1441),
.B1(n_1437),
.B2(n_1414),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1713),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1716),
.B(n_1489),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1715),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1718),
.A2(n_1437),
.B(n_1439),
.Y(n_1719)
);

NAND2xp33_ASAP7_75t_SL g1720 ( 
.A(n_1719),
.B(n_1717),
.Y(n_1720)
);

XNOR2xp5_ASAP7_75t_L g1721 ( 
.A(n_1720),
.B(n_1367),
.Y(n_1721)
);

AOI221xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1503),
.B1(n_1505),
.B2(n_1512),
.C(n_1414),
.Y(n_1722)
);

AOI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1367),
.B(n_1374),
.C(n_1370),
.Y(n_1723)
);


endmodule