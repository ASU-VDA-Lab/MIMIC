module fake_jpeg_14913_n_353 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_45),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_34),
.B1(n_19),
.B2(n_21),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_46),
.B1(n_28),
.B2(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_17),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_20),
.B1(n_28),
.B2(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_28),
.Y(n_89)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_18),
.B1(n_48),
.B2(n_54),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_46),
.B1(n_33),
.B2(n_21),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_73),
.B1(n_71),
.B2(n_34),
.Y(n_108)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_91),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_34),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_63),
.Y(n_110)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_94),
.Y(n_118)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_102),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_98),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_49),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_51),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_110),
.B(n_115),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_18),
.B(n_27),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_124),
.B(n_126),
.Y(n_153)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_88),
.CI(n_52),
.CON(n_115),
.SN(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_41),
.C(n_56),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_41),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_65),
.B1(n_74),
.B2(n_62),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_123),
.B1(n_30),
.B2(n_26),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_18),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_96),
.B(n_86),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_83),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_75),
.B1(n_104),
.B2(n_48),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_127),
.B1(n_77),
.B2(n_93),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_22),
.B(n_24),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_59),
.B1(n_75),
.B2(n_70),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_68),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_131),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_81),
.A2(n_30),
.B(n_26),
.C(n_37),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_145),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_93),
.B1(n_102),
.B2(n_81),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_144),
.B1(n_146),
.B2(n_151),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_143),
.B(n_160),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_101),
.B1(n_97),
.B2(n_90),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_90),
.B1(n_86),
.B2(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_116),
.A2(n_101),
.B1(n_36),
.B2(n_37),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_36),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_99),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_158),
.Y(n_172)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_99),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_129),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_134),
.B1(n_120),
.B2(n_110),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_175),
.B(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_115),
.B1(n_127),
.B2(n_120),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_170),
.B1(n_177),
.B2(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_115),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_135),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_115),
.B1(n_120),
.B2(n_108),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_133),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_0),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_118),
.B(n_105),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_155),
.A2(n_130),
.B1(n_106),
.B2(n_121),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_186),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_105),
.B(n_133),
.Y(n_181)
);

NOR2x1_ASAP7_75t_R g182 ( 
.A(n_140),
.B(n_121),
.Y(n_182)
);

FAx1_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_147),
.CI(n_141),
.CON(n_196),
.SN(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_138),
.A2(n_132),
.B1(n_112),
.B2(n_107),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_112),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_188),
.B(n_129),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_137),
.A2(n_107),
.B1(n_117),
.B2(n_61),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_139),
.B1(n_148),
.B2(n_107),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_142),
.A3(n_146),
.B1(n_144),
.B2(n_152),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_191),
.B(n_197),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_142),
.C(n_170),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_194),
.C(n_201),
.Y(n_218)
);

OAI22x1_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_143),
.B1(n_145),
.B2(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_206),
.B1(n_215),
.B2(n_183),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_151),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_189),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_195),
.B(n_189),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_210),
.B(n_178),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_165),
.B1(n_171),
.B2(n_174),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_139),
.Y(n_201)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_175),
.C(n_164),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_214),
.C(n_192),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_117),
.B1(n_157),
.B2(n_61),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_129),
.B(n_162),
.C(n_16),
.D(n_15),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_168),
.B(n_162),
.CI(n_1),
.CON(n_211),
.SN(n_211)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_164),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_163),
.A2(n_76),
.B1(n_69),
.B2(n_162),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_237),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_184),
.C(n_167),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_242),
.C(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_188),
.B(n_163),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_174),
.B1(n_171),
.B2(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_214),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_187),
.B1(n_172),
.B2(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_172),
.B(n_185),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_185),
.B1(n_76),
.B2(n_69),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_204),
.A2(n_200),
.B1(n_196),
.B2(n_197),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_211),
.B1(n_191),
.B2(n_207),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_241),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_51),
.C(n_98),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_235),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_247),
.A2(n_254),
.B(n_3),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_258),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_213),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_241),
.B(n_224),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_235),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_264),
.C(n_242),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_207),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_216),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_266),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_219),
.B(n_210),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_262),
.B(n_227),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_215),
.B(n_1),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_243),
.B(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_51),
.C(n_84),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_238),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_0),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_267),
.A2(n_270),
.B(n_284),
.Y(n_290)
);

NOR3xp33_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_220),
.C(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_275),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_231),
.B(n_232),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_229),
.C(n_230),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_240),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_236),
.C(n_234),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_223),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_234),
.C(n_233),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_281),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_233),
.C(n_241),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_3),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_3),
.C(n_4),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_276),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_251),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_265),
.B1(n_266),
.B2(n_257),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_278),
.A2(n_259),
.B1(n_246),
.B2(n_260),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_268),
.B1(n_274),
.B2(n_272),
.Y(n_309)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_8),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_301),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_259),
.B1(n_246),
.B2(n_252),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_295),
.A2(n_303),
.B1(n_281),
.B2(n_283),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_245),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_300),
.C(n_294),
.Y(n_314)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_263),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_267),
.B(n_4),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_279),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_287),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_312),
.Y(n_325)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_317),
.B(n_9),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_273),
.B(n_286),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_311),
.B(n_300),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_286),
.B(n_7),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_5),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_8),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_314),
.Y(n_326)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_318),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_295),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_9),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_291),
.Y(n_318)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_319),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_293),
.B(n_303),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_11),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_309),
.B1(n_290),
.B2(n_308),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_11),
.C(n_12),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_288),
.B1(n_301),
.B2(n_10),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_304),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_8),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_330),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_328),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_313),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_305),
.A2(n_9),
.B(n_10),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_336),
.Y(n_345)
);

XNOR2x1_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_304),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_338),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_333),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_339),
.B(n_328),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_9),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_340),
.B(n_334),
.Y(n_346)
);

O2A1O1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_339),
.A2(n_321),
.B(n_323),
.C(n_324),
.Y(n_342)
);

AOI21xp33_ASAP7_75t_L g347 ( 
.A1(n_342),
.A2(n_343),
.B(n_325),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_325),
.B(n_326),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_347),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_11),
.C(n_12),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_341),
.B(n_345),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_350),
.A2(n_348),
.B(n_12),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_12),
.B(n_13),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_13),
.B(n_335),
.Y(n_353)
);


endmodule