module fake_jpeg_6103_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx6p67_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_15),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_22),
.B1(n_11),
.B2(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_1),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_30),
.C(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_24),
.B(n_16),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_38),
.B(n_16),
.C(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_13),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_34),
.B(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_52),
.B(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_61),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_47),
.B1(n_43),
.B2(n_21),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_34),
.B(n_27),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_51),
.B(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_71),
.C(n_55),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_49),
.B(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_74),
.Y(n_75)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_78),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_87),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_60),
.C(n_59),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_95),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_79),
.B1(n_78),
.B2(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_88),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_73),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_92),
.B(n_35),
.Y(n_102)
);

OAI31xp33_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_92),
.A3(n_17),
.B(n_8),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_102),
.Y(n_104)
);

AOI21x1_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_3),
.B(n_4),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_4),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_9),
.A3(n_19),
.B1(n_26),
.B2(n_58),
.C1(n_74),
.C2(n_102),
.Y(n_108)
);


endmodule