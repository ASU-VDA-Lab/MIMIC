module real_jpeg_13478_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_56),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_3),
.A2(n_56),
.B1(n_69),
.B2(n_71),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_56),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_6),
.A2(n_63),
.B1(n_69),
.B2(n_71),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_63),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_69),
.B1(n_71),
.B2(n_87),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_9),
.A2(n_33),
.B1(n_69),
.B2(n_71),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_11),
.A2(n_37),
.B(n_38),
.C(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_11),
.B(n_106),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_11),
.A2(n_40),
.B1(n_69),
.B2(n_71),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_11),
.A2(n_81),
.B1(n_85),
.B2(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_11),
.B(n_74),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_13),
.A2(n_59),
.B1(n_69),
.B2(n_71),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_59),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_14),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_14),
.A2(n_69),
.B1(n_71),
.B2(n_76),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_76),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_20),
.B(n_107),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_47),
.B1(n_48),
.B2(n_77),
.Y(n_21)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_25),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_25),
.A2(n_84),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_25),
.A2(n_30),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_26),
.A2(n_27),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_26),
.B(n_40),
.C(n_90),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_26),
.B(n_170),
.Y(n_169)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_30),
.B(n_135),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_32),
.A2(n_85),
.B(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g132 ( 
.A(n_40),
.B(n_42),
.CON(n_132),
.SN(n_132)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_40),
.B(n_85),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_40),
.B(n_89),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_42),
.B1(n_67),
.B2(n_68),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_41),
.B(n_68),
.C(n_69),
.Y(n_133)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_60),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_55),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_73),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_65),
.B1(n_74),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_64),
.A2(n_66),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_65),
.A2(n_74),
.B1(n_120),
.B2(n_132),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

OA22x2_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_67),
.A2(n_71),
.B(n_131),
.C(n_133),
.Y(n_130)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_69),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_71),
.B1(n_90),
.B2(n_91),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_71),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_98),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_81),
.A2(n_85),
.B1(n_164),
.B2(n_172),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_81),
.A2(n_166),
.B(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B(n_93),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_139),
.B1(n_141),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_96),
.A2(n_141),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_96),
.A2(n_141),
.B1(n_149),
.B2(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.C(n_104),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_112),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_108),
.B(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_110),
.B(n_112),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_118),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_195),
.B(n_199),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_150),
.B(n_194),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_145),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_127),
.B(n_145),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_142),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_129),
.B(n_136),
.C(n_142),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_134),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B(n_140),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.C(n_148),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_148),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_189),
.B(n_193),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_178),
.B(n_188),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_167),
.B(n_177),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_162),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_160),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_173),
.B(n_176),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_180),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_184),
.C(n_187),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_192),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_198),
.Y(n_199)
);


endmodule