module real_jpeg_25867_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_244;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_1),
.B(n_69),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_1),
.B(n_27),
.C(n_41),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_106),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_1),
.B(n_114),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_24),
.B1(n_125),
.B2(n_212),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_2),
.A2(n_46),
.B1(n_63),
.B2(n_64),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_3),
.A2(n_35),
.B1(n_63),
.B2(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_5),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_71),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_71),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_7),
.A2(n_56),
.B1(n_67),
.B2(n_79),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_79),
.Y(n_155)
);

INVx8_ASAP7_75t_SL g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_9),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_118),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_118),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_118),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_10),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_58),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_58),
.Y(n_205)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_148),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_147),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_20),
.B(n_120),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_95),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_21),
.B(n_82),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_22),
.B(n_54),
.C(n_72),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_23),
.B(n_38),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_33),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_24),
.A2(n_88),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_24),
.A2(n_85),
.B(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_24),
.A2(n_205),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_24),
.A2(n_33),
.B(n_88),
.Y(n_230)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_25),
.B(n_34),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_25),
.A2(n_31),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_25),
.A2(n_172),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_26),
.B(n_217),
.Y(n_216)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_29),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_36),
.Y(n_213)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_37),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_37),
.B(n_106),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B(n_47),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_39),
.B(n_52),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_39),
.A2(n_49),
.B1(n_191),
.B2(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_39),
.B(n_106),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_40),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_42),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_44),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_43),
.A2(n_76),
.B(n_226),
.C(n_228),
.Y(n_225)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_44),
.B(n_187),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_44),
.B(n_63),
.C(n_75),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_48),
.A2(n_129),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_48),
.A2(n_92),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_48),
.A2(n_92),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_49),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_49),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_72),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_69),
.B2(n_70),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_55),
.Y(n_119)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_59),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_59),
.A2(n_69),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_60),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_64),
.B(n_105),
.C(n_108),
.Y(n_104)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_63),
.C(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_64),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g227 ( 
.A(n_64),
.B(n_106),
.CON(n_227),
.SN(n_227)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_68),
.A2(n_105),
.B(n_106),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_69),
.B(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_70),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_78),
.B(n_80),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_73),
.B(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_73),
.A2(n_111),
.B1(n_114),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_73),
.A2(n_114),
.B1(n_177),
.B2(n_227),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_77),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_77),
.A2(n_112),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_90),
.B2(n_94),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_94),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_89),
.A2(n_101),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_92),
.B(n_155),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_93),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_95),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_109),
.C(n_115),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_96),
.A2(n_97),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_104),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_109),
.B(n_115),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B(n_113),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_117),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_146),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_131),
.B1(n_144),
.B2(n_145),
.Y(n_121)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_130),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_138),
.B1(n_139),
.B2(n_143),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_179),
.B(n_260),
.C(n_264),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_164),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_150),
.B(n_164),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_161),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_152),
.B(n_153),
.C(n_161),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_158),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_169),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_165),
.B(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_169),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_175),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_175),
.B(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_259),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_254),
.B(n_258),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_238),
.B(n_253),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_221),
.B(n_237),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_201),
.B(n_220),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_192),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_188),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_196),
.C(n_199),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_208),
.B(n_219),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_207),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_214),
.B(n_218),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_236),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_236),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_231),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_232),
.C(n_233),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_230),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_240),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_248),
.C(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_262),
.Y(n_264)
);


endmodule