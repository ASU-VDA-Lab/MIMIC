module fake_jpeg_16765_n_209 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_16),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_36),
.B(n_33),
.C(n_35),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_41),
.A2(n_15),
.B(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_39),
.Y(n_66)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_18),
.CI(n_25),
.CON(n_83),
.SN(n_83)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_56),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_16),
.B1(n_31),
.B2(n_19),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_19),
.Y(n_78)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_41),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_26),
.C(n_37),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_72),
.C(n_30),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_64),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_31),
.B1(n_55),
.B2(n_45),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_65),
.A2(n_81),
.B1(n_32),
.B2(n_23),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_68),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_38),
.Y(n_70)
);

XOR2x1_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_20),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_74),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_27),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_80),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_87),
.B(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_83),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_43),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_54),
.B1(n_31),
.B2(n_32),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_34),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_49),
.B(n_17),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_38),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_111),
.C(n_83),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_37),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_98),
.Y(n_119)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_106),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_28),
.C(n_20),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_37),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2x1p5_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_32),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_21),
.B1(n_30),
.B2(n_28),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_17),
.B(n_29),
.C(n_15),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_61),
.B1(n_74),
.B2(n_60),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_60),
.B1(n_59),
.B2(n_85),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_81),
.B1(n_87),
.B2(n_85),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_124),
.C(n_109),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_84),
.B1(n_71),
.B2(n_80),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_83),
.C(n_69),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_29),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_129),
.Y(n_147)
);

AOI22x1_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_71),
.B1(n_82),
.B2(n_23),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_132),
.B1(n_89),
.B2(n_94),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_28),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_93),
.A2(n_21),
.B1(n_24),
.B2(n_4),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_131),
.A2(n_109),
.B1(n_110),
.B2(n_93),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_20),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_30),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_98),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_120),
.B(n_30),
.C(n_4),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_145),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_118),
.C(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_104),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_143),
.A2(n_152),
.B(n_125),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_148),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_110),
.B1(n_101),
.B2(n_97),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_100),
.C(n_30),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_124),
.C(n_154),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_100),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_153),
.B(n_154),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_89),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_167),
.B1(n_138),
.B2(n_143),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_160),
.C(n_161),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_122),
.C(n_116),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_117),
.C(n_131),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_142),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_159),
.C(n_13),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_162),
.B(n_144),
.C(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_177),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_143),
.B1(n_152),
.B2(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_178),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_155),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_153),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_167),
.B(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_142),
.B1(n_146),
.B2(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_179),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

NAND4xp25_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_167),
.C(n_156),
.D(n_160),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_188),
.B(n_2),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_167),
.B(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_172),
.C(n_176),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_2),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_195),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_176),
.C(n_173),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_13),
.C(n_12),
.Y(n_197)
);

OA21x2_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_11),
.B(n_6),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_192),
.A3(n_189),
.B1(n_187),
.B2(n_186),
.C1(n_183),
.C2(n_10),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_5),
.B(n_6),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_202),
.Y(n_207)
);

NAND4xp25_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_11),
.C(n_12),
.D(n_7),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_204),
.A2(n_196),
.B(n_194),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_206),
.A2(n_205),
.B1(n_207),
.B2(n_203),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_9),
.Y(n_209)
);


endmodule