module fake_jpeg_25225_n_246 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_21),
.B1(n_33),
.B2(n_29),
.Y(n_56)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_20),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_55),
.B1(n_35),
.B2(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_38),
.B1(n_17),
.B2(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_32),
.B1(n_25),
.B2(n_3),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_57),
.B1(n_47),
.B2(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_68),
.B1(n_35),
.B2(n_39),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_27),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_40),
.C(n_41),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_26),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_4),
.B(n_5),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_32),
.B1(n_17),
.B2(n_3),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_81),
.B1(n_64),
.B2(n_46),
.Y(n_95)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_57),
.B1(n_60),
.B2(n_47),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_80),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_1),
.B(n_2),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_79),
.B(n_84),
.Y(n_100)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_52),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_39),
.B1(n_43),
.B2(n_40),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_89),
.C(n_64),
.Y(n_96)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_85),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_41),
.A3(n_40),
.B1(n_7),
.B2(n_8),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_50),
.B1(n_51),
.B2(n_62),
.Y(n_110)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_40),
.C(n_6),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_99),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_107),
.B1(n_111),
.B2(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_96),
.B(n_115),
.Y(n_116)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_109),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_59),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_86),
.B1(n_82),
.B2(n_80),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_61),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_112),
.B1(n_4),
.B2(n_6),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_50),
.B1(n_63),
.B2(n_62),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_62),
.B1(n_55),
.B2(n_49),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_88),
.B1(n_74),
.B2(n_62),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_49),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_65),
.Y(n_129)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_121),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_65),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_130),
.B(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_129),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_73),
.B1(n_91),
.B2(n_71),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_78),
.B1(n_83),
.B2(n_77),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_60),
.B1(n_40),
.B2(n_53),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_60),
.B1(n_53),
.B2(n_65),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_4),
.B(n_6),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_115),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_7),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_130),
.B(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_8),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_145),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_100),
.B(n_96),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_146),
.B(n_154),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_107),
.C(n_114),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_153),
.C(n_156),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_102),
.A3(n_100),
.B1(n_104),
.B2(n_103),
.C1(n_109),
.C2(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_149),
.Y(n_169)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_93),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_112),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_152),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_105),
.B(n_106),
.C(n_97),
.D(n_13),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_97),
.C(n_106),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_9),
.B(n_10),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_159),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_9),
.C(n_12),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_136),
.B1(n_123),
.B2(n_132),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_143),
.A2(n_136),
.B1(n_128),
.B2(n_134),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_176),
.B1(n_148),
.B2(n_157),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_146),
.B1(n_159),
.B2(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_174),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_154),
.B1(n_152),
.B2(n_138),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_139),
.C(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_122),
.B1(n_138),
.B2(n_119),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_121),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_139),
.C(n_156),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_133),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

XOR2x2_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_141),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_192),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_166),
.C(n_179),
.Y(n_203)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_170),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_181),
.B1(n_176),
.B2(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_198),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_148),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

AOI321xp33_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_169),
.A3(n_175),
.B1(n_168),
.B2(n_174),
.C(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_201),
.B(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_163),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_208),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_166),
.C(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_206),
.C(n_211),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_172),
.C(n_177),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_165),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_187),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_120),
.B(n_161),
.Y(n_228)
);

AO22x1_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_184),
.B1(n_191),
.B2(n_194),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_221),
.B(n_182),
.C(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_183),
.B1(n_195),
.B2(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_203),
.C(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_223),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_182),
.B(n_186),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_226),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_120),
.Y(n_227)
);

O2A1O1Ixp5_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_214),
.B(n_127),
.C(n_207),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_212),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_234),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_207),
.B(n_217),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_15),
.B(n_16),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_16),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_212),
.C(n_15),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_229),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_235),
.B(n_233),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_241),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_236),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_244),
.Y(n_246)
);


endmodule