module fake_ibex_591_n_583 (n_85, n_84, n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_583);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_583;

wire n_151;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_165;
wire n_452;
wire n_255;
wire n_175;
wire n_398;
wire n_304;
wire n_125;
wire n_191;
wire n_153;
wire n_545;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_578;
wire n_478;
wire n_239;
wire n_94;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_531;
wire n_556;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_122;
wire n_523;
wire n_116;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_355;
wire n_474;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_536;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_98;
wire n_129;
wire n_267;
wire n_245;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_554;
wire n_553;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_365;
wire n_539;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_516;
wire n_548;
wire n_567;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_582;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_320;
wire n_285;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_318;
wire n_291;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_118;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_311;
wire n_406;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_202;
wire n_159;
wire n_231;
wire n_298;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_63),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_83),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

BUFx8_ASAP7_75t_SL g101 ( 
.A(n_29),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_33),
.Y(n_105)
);

INVx4_ASAP7_75t_R g106 ( 
.A(n_28),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_10),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_66),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_24),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_25),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_15),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_58),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_64),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_47),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_73),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_68),
.B(n_31),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_6),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_11),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_39),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_52),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_12),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_15),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_48),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_56),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_80),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_91),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_57),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_22),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_38),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_27),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_4),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_23),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_0),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_97),
.B(n_0),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_101),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_94),
.A2(n_122),
.B(n_153),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_107),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_117),
.B(n_5),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_122),
.A2(n_36),
.B(n_89),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_5),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_7),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_35),
.B(n_85),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_107),
.B(n_7),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_119),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_132),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_144),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

BUFx8_ASAP7_75t_L g202 ( 
.A(n_134),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_9),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_126),
.B(n_13),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_145),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_135),
.B(n_16),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_138),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_102),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_98),
.B(n_18),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

AND3x2_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_104),
.C(n_136),
.Y(n_227)
);

OR2x6_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_109),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_198),
.B1(n_168),
.B2(n_179),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_111),
.B1(n_113),
.B2(n_116),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_130),
.C(n_154),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_223),
.B(n_105),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_96),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_95),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_174),
.B(n_182),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_159),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_111),
.B1(n_113),
.B2(n_116),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_R g246 ( 
.A(n_208),
.B(n_150),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_129),
.C(n_147),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_166),
.A2(n_136),
.B1(n_127),
.B2(n_146),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_159),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_165),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_202),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_199),
.B(n_131),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_177),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_177),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_201),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_163),
.A2(n_127),
.B1(n_149),
.B2(n_133),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_223),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_180),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_184),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_169),
.B(n_106),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_184),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

AOI22x1_ASAP7_75t_L g271 ( 
.A1(n_186),
.A2(n_196),
.B1(n_216),
.B2(n_189),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

NAND2xp33_ASAP7_75t_R g273 ( 
.A(n_178),
.B(n_19),
.Y(n_273)
);

OR2x6_ASAP7_75t_L g274 ( 
.A(n_164),
.B(n_20),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_205),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_181),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_176),
.B(n_41),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_251),
.B(n_187),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_240),
.A2(n_187),
.B1(n_176),
.B2(n_217),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_164),
.B1(n_209),
.B2(n_217),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_240),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_243),
.B(n_203),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_161),
.C(n_220),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_254),
.B(n_203),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_211),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_253),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_195),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_229),
.B(n_211),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_226),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_195),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_248),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_232),
.A2(n_200),
.B1(n_212),
.B2(n_210),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_172),
.C(n_221),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_240),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_194),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_253),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_239),
.B(n_191),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_247),
.B(n_196),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_256),
.B(n_189),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_245),
.B(n_192),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_247),
.B(n_207),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_242),
.B(n_207),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_266),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_245),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_228),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_228),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_240),
.B(n_192),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_162),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_236),
.B(n_200),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_L g322 ( 
.A(n_233),
.B(n_201),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_231),
.A2(n_170),
.B(n_173),
.C(n_215),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_183),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_278),
.B(n_170),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_228),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_278),
.B(n_170),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_249),
.B(n_204),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_237),
.B(n_183),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_264),
.B(n_204),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_261),
.A2(n_204),
.B1(n_215),
.B2(n_214),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_238),
.B(n_204),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_264),
.B(n_215),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_290),
.B(n_250),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_274),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_282),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_227),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_268),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_292),
.B(n_297),
.Y(n_340)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_274),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_274),
.B(n_269),
.C(n_270),
.Y(n_343)
);

AOI221xp5_ASAP7_75t_L g344 ( 
.A1(n_299),
.A2(n_300),
.B1(n_319),
.B2(n_283),
.C(n_314),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_302),
.B(n_274),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_276),
.Y(n_347)
);

BUFx8_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_305),
.B(n_263),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_309),
.B(n_277),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_281),
.B(n_271),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_302),
.A2(n_214),
.B1(n_175),
.B2(n_173),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_324),
.A2(n_235),
.B(n_230),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_175),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_175),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_287),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_318),
.B(n_175),
.Y(n_361)
);

O2A1O1Ixp5_ASAP7_75t_L g362 ( 
.A1(n_329),
.A2(n_285),
.B(n_288),
.C(n_326),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_173),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_291),
.B(n_21),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_26),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_SL g366 ( 
.A(n_301),
.B(n_206),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_30),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_304),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g372 ( 
.A(n_332),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_312),
.Y(n_373)
);

INVx11_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_280),
.B(n_289),
.Y(n_375)
);

AOI22x1_ASAP7_75t_SL g376 ( 
.A1(n_325),
.A2(n_34),
.B1(n_37),
.B2(n_59),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_296),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_317),
.A2(n_284),
.B1(n_307),
.B2(n_310),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_311),
.A2(n_265),
.B1(n_259),
.B2(n_258),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_359),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_343),
.A2(n_333),
.B(n_303),
.C(n_334),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_333),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_342),
.B(n_331),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_344),
.B(n_322),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

OAI22x1_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_338),
.B1(n_335),
.B2(n_336),
.Y(n_388)
);

NAND3x1_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_67),
.C(n_72),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_377),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_348),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_SL g393 ( 
.A1(n_353),
.A2(n_241),
.B(n_255),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_77),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_78),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_357),
.B(n_260),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_345),
.B(n_365),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_345),
.B(n_341),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_350),
.A2(n_375),
.B(n_362),
.C(n_378),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_348),
.Y(n_401)
);

OAI22x1_ASAP7_75t_L g402 ( 
.A1(n_368),
.A2(n_365),
.B1(n_376),
.B2(n_341),
.Y(n_402)
);

NAND2x1_ASAP7_75t_L g403 ( 
.A(n_352),
.B(n_373),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_373),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_SL g405 ( 
.A(n_352),
.B(n_372),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_361),
.A2(n_363),
.B(n_358),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_346),
.A2(n_367),
.B(n_351),
.C(n_349),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_374),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_379),
.A2(n_354),
.B(n_366),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_340),
.Y(n_410)
);

OA22x2_ASAP7_75t_L g411 ( 
.A1(n_342),
.A2(n_228),
.B1(n_244),
.B2(n_283),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_340),
.B(n_344),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_336),
.B(n_279),
.Y(n_413)
);

CKINVDCx6p67_ASAP7_75t_R g414 ( 
.A(n_337),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_371),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_345),
.A2(n_299),
.B1(n_344),
.B2(n_300),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_348),
.Y(n_418)
);

AOI211x1_ASAP7_75t_L g419 ( 
.A1(n_356),
.A2(n_286),
.B(n_364),
.C(n_299),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_337),
.B(n_244),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_371),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_336),
.B(n_279),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_340),
.B(n_344),
.Y(n_423)
);

AO31x2_ASAP7_75t_L g424 ( 
.A1(n_356),
.A2(n_324),
.A3(n_330),
.B(n_353),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_371),
.A2(n_281),
.B1(n_374),
.B2(n_340),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_337),
.Y(n_426)
);

NOR4xp25_ASAP7_75t_L g427 ( 
.A(n_343),
.B(n_299),
.C(n_344),
.D(n_323),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_340),
.B(n_344),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_360),
.Y(n_429)
);

OR2x6_ASAP7_75t_L g430 ( 
.A(n_342),
.B(n_244),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_371),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_337),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_337),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_377),
.Y(n_434)
);

OAI21x1_ASAP7_75t_SL g435 ( 
.A1(n_343),
.A2(n_290),
.B(n_281),
.Y(n_435)
);

BUFx12f_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_377),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_429),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_411),
.A2(n_417),
.B1(n_430),
.B2(n_412),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_423),
.B(n_428),
.C(n_400),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

INVx5_ASAP7_75t_L g444 ( 
.A(n_390),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_396),
.B(n_413),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_383),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_391),
.Y(n_448)
);

NAND2x1p5_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_431),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_430),
.A2(n_402),
.B1(n_425),
.B2(n_408),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_436),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_414),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_430),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_415),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_384),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_409),
.A2(n_389),
.B(n_398),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_416),
.B(n_431),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_409),
.A2(n_403),
.B(n_435),
.Y(n_460)
);

BUFx12f_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

AND3x4_ASAP7_75t_L g462 ( 
.A(n_392),
.B(n_394),
.C(n_401),
.Y(n_462)
);

AOI21x1_ASAP7_75t_L g463 ( 
.A1(n_388),
.A2(n_386),
.B(n_399),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_419),
.B(n_421),
.Y(n_464)
);

AO31x2_ASAP7_75t_L g465 ( 
.A1(n_381),
.A2(n_407),
.A3(n_393),
.B(n_424),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_406),
.A2(n_404),
.B(n_410),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_420),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

AOI22x1_ASAP7_75t_L g472 ( 
.A1(n_395),
.A2(n_397),
.B1(n_434),
.B2(n_437),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_405),
.A2(n_437),
.B(n_419),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_424),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_424),
.B(n_412),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_412),
.B(n_423),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_418),
.Y(n_477)
);

NAND3xp33_ASAP7_75t_L g478 ( 
.A(n_419),
.B(n_202),
.C(n_417),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_385),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_423),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_466),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_448),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_443),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_443),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_480),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_460),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_445),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_441),
.B(n_453),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_475),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_442),
.Y(n_492)
);

INVx8_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_468),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_444),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_467),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_450),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_462),
.Y(n_498)
);

INVx8_ASAP7_75t_L g499 ( 
.A(n_493),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_482),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_460),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_468),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_465),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_486),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_483),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_465),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_487),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_484),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_465),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_464),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_464),
.Y(n_512)
);

NOR2x1_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_462),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_458),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_493),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_507),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_506),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_509),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_507),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_488),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_496),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_508),
.Y(n_522)
);

O2A1O1Ixp33_ASAP7_75t_SL g523 ( 
.A1(n_522),
.A2(n_515),
.B(n_500),
.C(n_502),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_519),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_512),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_511),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_517),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_511),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_505),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_509),
.Y(n_530)
);

NAND2x1_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_513),
.Y(n_531)
);

OAI21xp33_ASAP7_75t_L g532 ( 
.A1(n_522),
.A2(n_513),
.B(n_492),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_527),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_529),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_524),
.B(n_518),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_521),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_521),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_525),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_520),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_528),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_530),
.Y(n_542)
);

AOI32xp33_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_498),
.A3(n_540),
.B1(n_532),
.B2(n_539),
.Y(n_543)
);

AOI31xp33_ASAP7_75t_L g544 ( 
.A1(n_535),
.A2(n_523),
.A3(n_515),
.B(n_503),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_533),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_533),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_539),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_534),
.Y(n_548)
);

A2O1A1Ixp33_ASAP7_75t_L g549 ( 
.A1(n_544),
.A2(n_531),
.B(n_499),
.C(n_536),
.Y(n_549)
);

AOI32xp33_ASAP7_75t_L g550 ( 
.A1(n_542),
.A2(n_518),
.A3(n_525),
.B1(n_492),
.B2(n_520),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_545),
.Y(n_551)
);

AOI221xp5_ASAP7_75t_L g552 ( 
.A1(n_544),
.A2(n_455),
.B1(n_454),
.B2(n_447),
.C(n_478),
.Y(n_552)
);

AOI221xp5_ASAP7_75t_L g553 ( 
.A1(n_550),
.A2(n_543),
.B1(n_548),
.B2(n_542),
.C(n_547),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_549),
.B(n_541),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_SL g555 ( 
.A(n_552),
.B(n_477),
.C(n_452),
.Y(n_555)
);

NOR3xp33_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_451),
.C(n_456),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_554),
.B(n_461),
.Y(n_557)
);

NOR3xp33_ASAP7_75t_L g558 ( 
.A(n_556),
.B(n_553),
.C(n_456),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_L g559 ( 
.A(n_557),
.B(n_473),
.C(n_440),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_558),
.B(n_477),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_R g561 ( 
.A(n_559),
.B(n_461),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_560),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_561),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_562),
.B(n_551),
.Y(n_564)
);

AND3x1_ASAP7_75t_L g565 ( 
.A(n_563),
.B(n_489),
.C(n_470),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_563),
.A2(n_494),
.B1(n_546),
.B2(n_545),
.Y(n_566)
);

NOR2x1_ASAP7_75t_L g567 ( 
.A(n_564),
.B(n_439),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_566),
.A2(n_442),
.B(n_458),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_503),
.Y(n_569)
);

XOR2x1_ASAP7_75t_L g570 ( 
.A(n_565),
.B(n_472),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_495),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_567),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_569),
.A2(n_514),
.B1(n_471),
.B2(n_444),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_568),
.A2(n_493),
.B1(n_499),
.B2(n_514),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_567),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_571),
.B(n_499),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_572),
.B(n_484),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_575),
.A2(n_493),
.B(n_499),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_576),
.A2(n_574),
.B(n_573),
.Y(n_579)
);

AOI21xp33_ASAP7_75t_L g580 ( 
.A1(n_577),
.A2(n_499),
.B(n_444),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_578),
.A2(n_463),
.B(n_444),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_579),
.A2(n_497),
.B(n_514),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_582),
.A2(n_580),
.B1(n_581),
.B2(n_474),
.Y(n_583)
);


endmodule