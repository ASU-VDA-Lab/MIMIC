module fake_netlist_1_2380_n_1583 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_383, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_384, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_381, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_382, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_385, n_257, n_269, n_1583);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_383;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_384;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_381;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_382;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_385;
input n_257;
input n_269;
output n_1583;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1460;
wire n_1372;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_1570;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1486;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1291;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_600;
wire n_1531;
wire n_1548;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1442;
INVx1_ASAP7_75t_L g386 ( .A(n_213), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_368), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_15), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_33), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_224), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_14), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_131), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_173), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_365), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_270), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_58), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_246), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_316), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_186), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_1), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_70), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_65), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_46), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_218), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_245), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_380), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_94), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_5), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_227), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_327), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_0), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_313), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_129), .B(n_299), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_280), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_278), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_361), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_315), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_2), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_267), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_363), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_48), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_317), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_125), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_336), .Y(n_424) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_142), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_201), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_183), .Y(n_427) );
CKINVDCx14_ASAP7_75t_R g428 ( .A(n_124), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_351), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_279), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_92), .Y(n_431) );
NOR2xp67_ASAP7_75t_L g432 ( .A(n_134), .B(n_127), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_70), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_135), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_28), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_367), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_268), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_346), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_288), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_220), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_109), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_210), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_300), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_42), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_78), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_303), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_337), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_196), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_301), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_214), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_119), .B(n_178), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_117), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_130), .B(n_182), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_304), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_110), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_334), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_296), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_160), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_379), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_118), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_341), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_140), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_322), .Y(n_463) );
NOR2xp67_ASAP7_75t_L g464 ( .A(n_373), .B(n_235), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_222), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_143), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_203), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_124), .B(n_159), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_243), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_311), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_22), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_332), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_305), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_31), .Y(n_474) );
BUFx10_ASAP7_75t_L g475 ( .A(n_291), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_233), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_369), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_383), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_293), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_287), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_116), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_74), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_378), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_381), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_160), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_325), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_360), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_211), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_323), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_331), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_73), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_145), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_298), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_190), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_105), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_297), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_81), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_206), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_69), .Y(n_499) );
BUFx10_ASAP7_75t_L g500 ( .A(n_371), .Y(n_500) );
CKINVDCx14_ASAP7_75t_R g501 ( .A(n_384), .Y(n_501) );
NOR2xp67_ASAP7_75t_L g502 ( .A(n_132), .B(n_105), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_147), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_98), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_187), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_28), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_312), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_168), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_290), .Y(n_509) );
BUFx2_ASAP7_75t_L g510 ( .A(n_50), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_302), .Y(n_511) );
INVxp33_ASAP7_75t_SL g512 ( .A(n_326), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_321), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_116), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_294), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_111), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_241), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_174), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_126), .B(n_32), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_61), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_69), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_274), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_134), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_230), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_263), .B(n_333), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_320), .Y(n_526) );
NOR2xp67_ASAP7_75t_L g527 ( .A(n_231), .B(n_68), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_132), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_149), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_353), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_97), .Y(n_531) );
BUFx3_ASAP7_75t_L g532 ( .A(n_318), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_286), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_277), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_364), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_342), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_237), .Y(n_537) );
XOR2xp5_ASAP7_75t_L g538 ( .A(n_314), .B(n_129), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_180), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_65), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_52), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_309), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_223), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_377), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_330), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_4), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_215), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_64), .Y(n_548) );
CKINVDCx14_ASAP7_75t_R g549 ( .A(n_54), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_244), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_113), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_88), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_207), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_61), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_306), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_329), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_198), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_184), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_254), .Y(n_559) );
CKINVDCx14_ASAP7_75t_R g560 ( .A(n_38), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_58), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_27), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g563 ( .A(n_43), .B(n_257), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_152), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_202), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_41), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_19), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_93), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_362), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_112), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_352), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_80), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_262), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_295), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_292), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_119), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_366), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_370), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_77), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_27), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_171), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_199), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_67), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_165), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_50), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_348), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_236), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_118), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_289), .Y(n_589) );
CKINVDCx16_ASAP7_75t_R g590 ( .A(n_108), .Y(n_590) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_48), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_212), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_283), .Y(n_593) );
BUFx6f_ASAP7_75t_SL g594 ( .A(n_338), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_276), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_392), .Y(n_596) );
INVx3_ASAP7_75t_L g597 ( .A(n_475), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_406), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_456), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_456), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_428), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_392), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_428), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_456), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_549), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_555), .B(n_3), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_567), .B(n_6), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_456), .Y(n_608) );
BUFx12f_ASAP7_75t_L g609 ( .A(n_475), .Y(n_609) );
NAND2xp33_ASAP7_75t_L g610 ( .A(n_425), .B(n_163), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_396), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_396), .B(n_6), .Y(n_612) );
INVx5_ASAP7_75t_L g613 ( .A(n_398), .Y(n_613) );
AND2x2_ASAP7_75t_SL g614 ( .A(n_525), .B(n_164), .Y(n_614) );
AND2x4_ASAP7_75t_L g615 ( .A(n_441), .B(n_7), .Y(n_615) );
OA21x2_ASAP7_75t_L g616 ( .A1(n_437), .A2(n_167), .B(n_166), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_475), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_441), .B(n_7), .Y(n_618) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_437), .A2(n_170), .B(n_169), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_586), .B(n_8), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_549), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_489), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_455), .B(n_8), .Y(n_623) );
INVx6_ASAP7_75t_L g624 ( .A(n_500), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_504), .B(n_9), .Y(n_625) );
AOI22x1_ASAP7_75t_SL g626 ( .A1(n_401), .A2(n_11), .B1(n_9), .B2(n_10), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_446), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_446), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_500), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_483), .B(n_10), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_497), .Y(n_631) );
INVx6_ASAP7_75t_L g632 ( .A(n_500), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_497), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g634 ( .A(n_425), .B(n_172), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_523), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_398), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_470), .B(n_11), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_560), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_510), .B(n_12), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_597), .B(n_526), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_627), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_597), .B(n_470), .Y(n_642) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_601), .A2(n_403), .B1(n_590), .B2(n_458), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_603), .B(n_501), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_597), .B(n_476), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_612), .A2(n_560), .B1(n_400), .B2(n_402), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_636), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_627), .Y(n_648) );
NOR2xp33_ASAP7_75t_SL g649 ( .A(n_614), .B(n_594), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_597), .B(n_404), .Y(n_650) );
AO22x2_ASAP7_75t_L g651 ( .A1(n_626), .A2(n_538), .B1(n_591), .B2(n_488), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_627), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_612), .A2(n_408), .B1(n_411), .B2(n_388), .Y(n_653) );
INVx3_ASAP7_75t_L g654 ( .A(n_612), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_636), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_612), .A2(n_421), .B1(n_423), .B2(n_418), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_636), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_612), .B(n_387), .C(n_386), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_597), .B(n_404), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_624), .B(n_416), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_617), .B(n_476), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_603), .B(n_501), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_619), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_636), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_621), .B(n_391), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_628), .Y(n_666) );
OR2x6_ASAP7_75t_L g667 ( .A(n_609), .B(n_432), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_617), .B(n_391), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_628), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_617), .B(n_488), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_621), .B(n_407), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_615), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_617), .B(n_412), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_636), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_624), .B(n_479), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_628), .Y(n_676) );
INVxp67_ASAP7_75t_SL g677 ( .A(n_638), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_617), .B(n_412), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_638), .B(n_433), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_629), .B(n_517), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_629), .B(n_517), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_649), .A2(n_614), .B1(n_606), .B2(n_615), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_647), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_640), .B(n_644), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_649), .B(n_614), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_640), .B(n_629), .Y(n_686) );
BUFx8_ASAP7_75t_L g687 ( .A(n_644), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_644), .B(n_629), .Y(n_688) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_662), .A2(n_626), .B1(n_614), .B2(n_499), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_662), .B(n_629), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_647), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_654), .A2(n_606), .B1(n_672), .B2(n_658), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_677), .A2(n_606), .B1(n_625), .B2(n_623), .Y(n_693) );
AND2x4_ASAP7_75t_SL g694 ( .A(n_667), .B(n_394), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_677), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_663), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_679), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_665), .B(n_624), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_665), .B(n_609), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_679), .B(n_623), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_665), .B(n_623), .Y(n_701) );
BUFx2_ASAP7_75t_L g702 ( .A(n_671), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_642), .A2(n_619), .B(n_610), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_671), .B(n_624), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_671), .B(n_624), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_650), .B(n_609), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_646), .A2(n_606), .B1(n_639), .B2(n_625), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_663), .B(n_606), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_668), .B(n_632), .Y(n_709) );
BUFx3_ASAP7_75t_L g710 ( .A(n_654), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_668), .B(n_632), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_668), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_668), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_660), .B(n_632), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_675), .B(n_632), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_659), .B(n_632), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_642), .B(n_632), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_645), .B(n_625), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_663), .B(n_615), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_654), .A2(n_615), .B1(n_618), .B2(n_639), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_645), .B(n_639), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_653), .B(n_630), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_654), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_672), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_672), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_672), .A2(n_618), .B1(n_630), .B2(n_620), .Y(n_726) );
NAND2x1p5_ASAP7_75t_L g727 ( .A(n_673), .B(n_618), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_661), .B(n_620), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_663), .B(n_618), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_658), .A2(n_619), .B(n_616), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_653), .B(n_622), .C(n_598), .Y(n_731) );
AND2x2_ASAP7_75t_SL g732 ( .A(n_656), .B(n_618), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_655), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_678), .B(n_607), .Y(n_734) );
O2A1O1Ixp5_ASAP7_75t_L g735 ( .A1(n_661), .A2(n_637), .B(n_607), .C(n_507), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_655), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_641), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_670), .B(n_417), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_680), .B(n_419), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_667), .B(n_512), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_655), .Y(n_741) );
INVx3_ASAP7_75t_L g742 ( .A(n_641), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_680), .B(n_419), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_681), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_663), .B(n_393), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_681), .B(n_465), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_643), .B(n_605), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_643), .A2(n_601), .B1(n_605), .B2(n_394), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_648), .Y(n_749) );
INVxp67_ASAP7_75t_L g750 ( .A(n_667), .Y(n_750) );
BUFx3_ASAP7_75t_L g751 ( .A(n_652), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_657), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_667), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_667), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_652), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g756 ( .A1(n_666), .A2(n_602), .B(n_611), .C(n_596), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_666), .B(n_530), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_663), .A2(n_637), .B1(n_512), .B2(n_407), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_669), .A2(n_434), .B1(n_435), .B2(n_431), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_667), .A2(n_439), .B1(n_505), .B2(n_426), .Y(n_760) );
O2A1O1Ixp33_ASAP7_75t_L g761 ( .A1(n_676), .A2(n_519), .B(n_602), .C(n_596), .Y(n_761) );
O2A1O1Ixp33_ASAP7_75t_L g762 ( .A1(n_676), .A2(n_631), .B(n_633), .C(n_611), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_657), .Y(n_763) );
BUFx2_ASAP7_75t_L g764 ( .A(n_651), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_657), .B(n_530), .Y(n_765) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_751), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_708), .A2(n_616), .B(n_634), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g768 ( .A1(n_730), .A2(n_616), .B(n_664), .Y(n_768) );
AND2x4_ASAP7_75t_L g769 ( .A(n_695), .B(n_468), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_712), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_703), .A2(n_616), .B(n_664), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_718), .B(n_462), .Y(n_772) );
A2O1A1Ixp33_ASAP7_75t_L g773 ( .A1(n_682), .A2(n_445), .B(n_452), .C(n_444), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_708), .A2(n_616), .B(n_664), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_685), .A2(n_439), .B1(n_505), .B2(n_426), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_732), .A2(n_508), .B1(n_401), .B2(n_499), .Y(n_776) );
NOR3xp33_ASAP7_75t_L g777 ( .A(n_689), .B(n_495), .C(n_389), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_732), .A2(n_651), .B1(n_520), .B2(n_508), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_SL g779 ( .A1(n_745), .A2(n_397), .B(n_399), .C(n_395), .Y(n_779) );
OR2x6_ASAP7_75t_L g780 ( .A(n_747), .B(n_651), .Y(n_780) );
INVx5_ASAP7_75t_L g781 ( .A(n_742), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_742), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_721), .B(n_466), .Y(n_783) );
BUFx4f_ASAP7_75t_L g784 ( .A(n_694), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_SL g785 ( .A1(n_706), .A2(n_674), .B(n_453), .C(n_413), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_728), .B(n_466), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_742), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g788 ( .A(n_687), .B(n_536), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_701), .B(n_471), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g790 ( .A(n_687), .B(n_697), .Y(n_790) );
BUFx8_ASAP7_75t_L g791 ( .A(n_764), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_685), .A2(n_520), .B1(n_651), .B2(n_531), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_701), .B(n_471), .Y(n_793) );
INVx2_ASAP7_75t_SL g794 ( .A(n_687), .Y(n_794) );
NOR2xp33_ASAP7_75t_SL g795 ( .A(n_694), .B(n_531), .Y(n_795) );
BUFx6f_ASAP7_75t_L g796 ( .A(n_696), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_693), .B(n_548), .Y(n_797) );
A2O1A1Ixp33_ASAP7_75t_L g798 ( .A1(n_734), .A2(n_485), .B(n_492), .C(n_491), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_722), .B(n_548), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_722), .B(n_561), .Y(n_800) );
INVxp33_ASAP7_75t_SL g801 ( .A(n_760), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_707), .A2(n_651), .B1(n_572), .B2(n_561), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_750), .B(n_572), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_747), .B(n_474), .Y(n_804) );
INVx6_ASAP7_75t_L g805 ( .A(n_710), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_686), .B(n_481), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_699), .B(n_503), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_738), .B(n_536), .Y(n_808) );
AND2x2_ASAP7_75t_SL g809 ( .A(n_748), .B(n_523), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_739), .B(n_583), .Y(n_810) );
NOR2xp33_ASAP7_75t_SL g811 ( .A(n_753), .B(n_594), .Y(n_811) );
NOR2xp33_ASAP7_75t_SL g812 ( .A(n_753), .B(n_543), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_723), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g814 ( .A(n_743), .B(n_746), .Y(n_814) );
AOI21x1_ASAP7_75t_L g815 ( .A1(n_719), .A2(n_464), .B(n_409), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_726), .B(n_543), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_719), .A2(n_410), .B(n_405), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_729), .A2(n_415), .B(n_414), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_740), .A2(n_547), .B1(n_550), .B2(n_544), .Y(n_819) );
O2A1O1Ixp33_ASAP7_75t_SL g820 ( .A1(n_745), .A2(n_430), .B(n_436), .C(n_420), .Y(n_820) );
AO22x1_ASAP7_75t_L g821 ( .A1(n_754), .A2(n_702), .B1(n_547), .B2(n_550), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_723), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_731), .B(n_506), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_720), .A2(n_553), .B1(n_556), .B2(n_544), .Y(n_824) );
O2A1O1Ixp5_ASAP7_75t_L g825 ( .A1(n_735), .A2(n_582), .B(n_559), .C(n_438), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_710), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_688), .B(n_514), .Y(n_827) );
OR2x6_ASAP7_75t_L g828 ( .A(n_690), .B(n_502), .Y(n_828) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_696), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_698), .B(n_553), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g831 ( .A1(n_729), .A2(n_443), .B(n_442), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_717), .A2(n_449), .B(n_448), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_714), .A2(n_454), .B(n_450), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_713), .Y(n_834) );
OR2x6_ASAP7_75t_L g835 ( .A(n_727), .B(n_568), .Y(n_835) );
NAND3xp33_ASAP7_75t_L g836 ( .A(n_758), .B(n_569), .C(n_558), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_713), .Y(n_837) );
OAI21xp5_ASAP7_75t_L g838 ( .A1(n_724), .A2(n_459), .B(n_457), .Y(n_838) );
A2O1A1Ixp33_ASAP7_75t_L g839 ( .A1(n_762), .A2(n_516), .B(n_528), .C(n_521), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_704), .B(n_540), .Y(n_840) );
OR2x6_ASAP7_75t_L g841 ( .A(n_727), .B(n_761), .Y(n_841) );
O2A1O1Ixp33_ASAP7_75t_SL g842 ( .A1(n_756), .A2(n_467), .B(n_469), .C(n_463), .Y(n_842) );
A2O1A1Ixp33_ASAP7_75t_L g843 ( .A1(n_725), .A2(n_546), .B(n_551), .C(n_541), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_705), .B(n_552), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_692), .B(n_554), .Y(n_845) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_709), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_757), .B(n_562), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_737), .Y(n_848) );
NAND2xp5_ASAP7_75t_SL g849 ( .A(n_711), .B(n_390), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_749), .A2(n_566), .B1(n_570), .B2(n_564), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_755), .B(n_579), .Y(n_851) );
A2O1A1Ixp33_ASAP7_75t_SL g852 ( .A1(n_716), .A2(n_633), .B(n_635), .C(n_631), .Y(n_852) );
BUFx6f_ASAP7_75t_L g853 ( .A(n_696), .Y(n_853) );
NAND3xp33_ASAP7_75t_L g854 ( .A(n_759), .B(n_613), .C(n_477), .Y(n_854) );
AOI21xp5_ASAP7_75t_L g855 ( .A1(n_715), .A2(n_478), .B(n_473), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_756), .B(n_580), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g857 ( .A1(n_683), .A2(n_484), .B(n_480), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_765), .B(n_588), .Y(n_858) );
OA22x2_ASAP7_75t_L g859 ( .A1(n_683), .A2(n_635), .B1(n_576), .B2(n_585), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_691), .Y(n_860) );
A2O1A1Ixp33_ASAP7_75t_L g861 ( .A1(n_691), .A2(n_527), .B(n_563), .C(n_451), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_733), .A2(n_460), .B1(n_482), .B2(n_425), .Y(n_862) );
OR2x2_ASAP7_75t_L g863 ( .A(n_736), .B(n_12), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_736), .B(n_422), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_741), .B(n_460), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_752), .A2(n_482), .B1(n_529), .B2(n_460), .Y(n_866) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_752), .A2(n_487), .B(n_486), .Y(n_867) );
O2A1O1Ixp33_ASAP7_75t_L g868 ( .A1(n_763), .A2(n_493), .B(n_496), .C(n_490), .Y(n_868) );
INVx1_ASAP7_75t_SL g869 ( .A(n_700), .Y(n_869) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_730), .A2(n_518), .B(n_511), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_712), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_730), .A2(n_524), .B(n_522), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_694), .Y(n_873) );
OAI21xp33_ASAP7_75t_L g874 ( .A1(n_697), .A2(n_427), .B(n_424), .Y(n_874) );
INVx4_ASAP7_75t_L g875 ( .A(n_751), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_712), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_712), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_708), .A2(n_535), .B(n_533), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_682), .A2(n_529), .B1(n_482), .B2(n_537), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_682), .A2(n_529), .B1(n_542), .B2(n_539), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_712), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_682), .A2(n_529), .B1(n_557), .B2(n_545), .Y(n_882) );
BUFx4f_ASAP7_75t_SL g883 ( .A(n_687), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_697), .B(n_534), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_684), .B(n_440), .Y(n_885) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_751), .Y(n_886) );
AND2x4_ASAP7_75t_L g887 ( .A(n_695), .B(n_565), .Y(n_887) );
A2O1A1Ixp33_ASAP7_75t_L g888 ( .A1(n_682), .A2(n_575), .B(n_581), .C(n_571), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_732), .A2(n_636), .B1(n_587), .B2(n_589), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_708), .A2(n_592), .B(n_584), .Y(n_890) );
NAND2xp5_ASAP7_75t_SL g891 ( .A(n_744), .B(n_461), .Y(n_891) );
BUFx2_ASAP7_75t_L g892 ( .A(n_687), .Y(n_892) );
AOI21xp5_ASAP7_75t_L g893 ( .A1(n_708), .A2(n_595), .B(n_613), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_682), .A2(n_494), .B1(n_513), .B2(n_472), .Y(n_894) );
NAND2xp5_ASAP7_75t_SL g895 ( .A(n_744), .B(n_515), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_802), .A2(n_636), .B1(n_574), .B2(n_577), .C(n_573), .Y(n_896) );
OAI21x1_ASAP7_75t_L g897 ( .A1(n_771), .A2(n_600), .B(n_599), .Y(n_897) );
O2A1O1Ixp5_ASAP7_75t_L g898 ( .A1(n_785), .A2(n_600), .B(n_604), .C(n_599), .Y(n_898) );
BUFx3_ASAP7_75t_L g899 ( .A(n_883), .Y(n_899) );
OAI22x1_ASAP7_75t_L g900 ( .A1(n_775), .A2(n_593), .B1(n_578), .B2(n_15), .Y(n_900) );
AO32x2_ASAP7_75t_L g901 ( .A1(n_880), .A2(n_882), .A3(n_879), .B1(n_792), .B2(n_850), .Y(n_901) );
AOI21xp5_ASAP7_75t_L g902 ( .A1(n_774), .A2(n_613), .B(n_447), .Y(n_902) );
OR2x2_ASAP7_75t_L g903 ( .A(n_776), .B(n_13), .Y(n_903) );
OAI21x1_ASAP7_75t_L g904 ( .A1(n_768), .A2(n_608), .B(n_604), .Y(n_904) );
OAI21xp5_ASAP7_75t_L g905 ( .A1(n_870), .A2(n_613), .B(n_608), .Y(n_905) );
AOI21xp5_ASAP7_75t_L g906 ( .A1(n_767), .A2(n_613), .B(n_447), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_848), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_801), .B(n_14), .Y(n_908) );
AO31x2_ASAP7_75t_L g909 ( .A1(n_888), .A2(n_498), .A3(n_509), .B(n_429), .Y(n_909) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_780), .A2(n_498), .B1(n_509), .B2(n_429), .Y(n_910) );
AOI21xp5_ASAP7_75t_L g911 ( .A1(n_814), .A2(n_613), .B(n_532), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_851), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_804), .B(n_780), .Y(n_913) );
AOI21xp5_ASAP7_75t_L g914 ( .A1(n_872), .A2(n_613), .B(n_175), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_863), .Y(n_915) );
AOI22xp5_ASAP7_75t_L g916 ( .A1(n_777), .A2(n_18), .B1(n_16), .B2(n_17), .Y(n_916) );
AO31x2_ASAP7_75t_L g917 ( .A1(n_861), .A2(n_19), .A3(n_17), .B(n_18), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g918 ( .A1(n_796), .A2(n_177), .B(n_176), .Y(n_918) );
AND2x4_ASAP7_75t_L g919 ( .A(n_794), .B(n_20), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_770), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_871), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_786), .B(n_21), .Y(n_922) );
OAI21xp5_ASAP7_75t_L g923 ( .A1(n_825), .A2(n_181), .B(n_179), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_860), .Y(n_924) );
OAI221xp5_ASAP7_75t_L g925 ( .A1(n_778), .A2(n_24), .B1(n_22), .B2(n_23), .C(n_25), .Y(n_925) );
A2O1A1Ixp33_ASAP7_75t_L g926 ( .A1(n_847), .A2(n_26), .B(n_23), .C(n_24), .Y(n_926) );
AOI221xp5_ASAP7_75t_SL g927 ( .A1(n_798), .A2(n_26), .B1(n_29), .B2(n_30), .C(n_31), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_876), .Y(n_928) );
AOI221xp5_ASAP7_75t_SL g929 ( .A1(n_773), .A2(n_29), .B1(n_30), .B2(n_32), .C(n_33), .Y(n_929) );
BUFx3_ASAP7_75t_L g930 ( .A(n_892), .Y(n_930) );
BUFx3_ASAP7_75t_L g931 ( .A(n_784), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_795), .A2(n_36), .B1(n_34), .B2(n_35), .Y(n_932) );
OAI21xp5_ASAP7_75t_L g933 ( .A1(n_839), .A2(n_34), .B(n_35), .Y(n_933) );
AO21x2_ASAP7_75t_L g934 ( .A1(n_852), .A2(n_188), .B(n_185), .Y(n_934) );
CKINVDCx8_ASAP7_75t_R g935 ( .A(n_873), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_796), .A2(n_191), .B(n_189), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_877), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_799), .B(n_36), .Y(n_938) );
INVx3_ASAP7_75t_L g939 ( .A(n_875), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g940 ( .A1(n_796), .A2(n_193), .B(n_192), .Y(n_940) );
OA21x2_ASAP7_75t_L g941 ( .A1(n_838), .A2(n_195), .B(n_194), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_881), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_865), .Y(n_943) );
AND2x2_ASAP7_75t_L g944 ( .A(n_784), .B(n_37), .Y(n_944) );
OAI21x1_ASAP7_75t_L g945 ( .A1(n_893), .A2(n_200), .B(n_197), .Y(n_945) );
OAI21x1_ASAP7_75t_SL g946 ( .A1(n_875), .A2(n_38), .B(n_39), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_800), .B(n_39), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_829), .A2(n_205), .B(n_204), .Y(n_948) );
NOR2xp33_ASAP7_75t_L g949 ( .A(n_790), .B(n_40), .Y(n_949) );
BUFx3_ASAP7_75t_L g950 ( .A(n_766), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_772), .B(n_40), .Y(n_951) );
INVx5_ASAP7_75t_L g952 ( .A(n_766), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_889), .A2(n_43), .B1(n_41), .B2(n_42), .Y(n_953) );
O2A1O1Ixp33_ASAP7_75t_L g954 ( .A1(n_843), .A2(n_46), .B(n_44), .C(n_45), .Y(n_954) );
AND2x4_ASAP7_75t_L g955 ( .A(n_781), .B(n_44), .Y(n_955) );
AND2x4_ASAP7_75t_L g956 ( .A(n_781), .B(n_45), .Y(n_956) );
AO21x2_ASAP7_75t_L g957 ( .A1(n_842), .A2(n_209), .B(n_208), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g958 ( .A1(n_823), .A2(n_841), .B1(n_807), .B2(n_827), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_884), .B(n_47), .Y(n_959) );
AO31x2_ASAP7_75t_L g960 ( .A1(n_858), .A2(n_51), .A3(n_47), .B(n_49), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_829), .A2(n_217), .B(n_216), .Y(n_961) );
INVx3_ASAP7_75t_L g962 ( .A(n_781), .Y(n_962) );
INVx4_ASAP7_75t_L g963 ( .A(n_766), .Y(n_963) );
AOI21xp5_ASAP7_75t_L g964 ( .A1(n_829), .A2(n_221), .B(n_219), .Y(n_964) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_853), .A2(n_226), .B(n_225), .Y(n_965) );
AOI21xp5_ASAP7_75t_L g966 ( .A1(n_853), .A2(n_229), .B(n_228), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_841), .A2(n_52), .B1(n_49), .B2(n_51), .Y(n_967) );
AOI21xp5_ASAP7_75t_L g968 ( .A1(n_853), .A2(n_234), .B(n_232), .Y(n_968) );
CKINVDCx5p33_ASAP7_75t_R g969 ( .A(n_791), .Y(n_969) );
A2O1A1Ixp33_ASAP7_75t_L g970 ( .A1(n_868), .A2(n_55), .B(n_53), .C(n_54), .Y(n_970) );
INVx2_ASAP7_75t_SL g971 ( .A(n_835), .Y(n_971) );
A2O1A1Ixp33_ASAP7_75t_L g972 ( .A1(n_832), .A2(n_56), .B(n_53), .C(n_55), .Y(n_972) );
O2A1O1Ixp33_ASAP7_75t_L g973 ( .A1(n_789), .A2(n_59), .B(n_56), .C(n_57), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_783), .B(n_57), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_886), .Y(n_975) );
OA21x2_ASAP7_75t_L g976 ( .A1(n_856), .A2(n_239), .B(n_238), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_797), .B(n_59), .Y(n_977) );
NAND3xp33_ASAP7_75t_L g978 ( .A(n_828), .B(n_60), .C(n_62), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g979 ( .A1(n_835), .A2(n_63), .B1(n_60), .B2(n_62), .Y(n_979) );
INVx1_ASAP7_75t_SL g980 ( .A(n_886), .Y(n_980) );
OAI21x1_ASAP7_75t_L g981 ( .A1(n_857), .A2(n_242), .B(n_240), .Y(n_981) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_793), .B(n_63), .Y(n_982) );
OAI21xp5_ASAP7_75t_L g983 ( .A1(n_878), .A2(n_248), .B(n_247), .Y(n_983) );
AOI31xp67_ASAP7_75t_L g984 ( .A1(n_840), .A2(n_385), .A3(n_382), .B(n_376), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_887), .B(n_803), .Y(n_985) );
AO21x2_ASAP7_75t_L g986 ( .A1(n_779), .A2(n_250), .B(n_249), .Y(n_986) );
OAI22x1_ASAP7_75t_L g987 ( .A1(n_788), .A2(n_64), .B1(n_66), .B2(n_67), .Y(n_987) );
OAI21xp5_ASAP7_75t_L g988 ( .A1(n_890), .A2(n_252), .B(n_251), .Y(n_988) );
O2A1O1Ixp33_ASAP7_75t_SL g989 ( .A1(n_787), .A2(n_375), .B(n_374), .C(n_372), .Y(n_989) );
BUFx6f_ASAP7_75t_L g990 ( .A(n_886), .Y(n_990) );
OAI21xp5_ASAP7_75t_L g991 ( .A1(n_817), .A2(n_255), .B(n_253), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_887), .B(n_66), .Y(n_992) );
OAI21xp5_ASAP7_75t_L g993 ( .A1(n_818), .A2(n_68), .B(n_71), .Y(n_993) );
INVx2_ASAP7_75t_SL g994 ( .A(n_791), .Y(n_994) );
NAND2x1p5_ASAP7_75t_L g995 ( .A(n_782), .B(n_71), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_844), .B(n_72), .Y(n_996) );
CKINVDCx11_ASAP7_75t_R g997 ( .A(n_828), .Y(n_997) );
OAI21xp5_ASAP7_75t_SL g998 ( .A1(n_819), .A2(n_72), .B(n_73), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_782), .A2(n_846), .B1(n_845), .B2(n_885), .Y(n_999) );
OAI21xp5_ASAP7_75t_L g1000 ( .A1(n_831), .A2(n_258), .B(n_256), .Y(n_1000) );
INVx2_ASAP7_75t_SL g1001 ( .A(n_821), .Y(n_1001) );
OAI21xp5_ASAP7_75t_L g1002 ( .A1(n_833), .A2(n_260), .B(n_259), .Y(n_1002) );
NAND2xp33_ASAP7_75t_L g1003 ( .A(n_826), .B(n_261), .Y(n_1003) );
BUFx6f_ASAP7_75t_L g1004 ( .A(n_805), .Y(n_1004) );
BUFx10_ASAP7_75t_L g1005 ( .A(n_769), .Y(n_1005) );
A2O1A1Ixp33_ASAP7_75t_L g1006 ( .A1(n_855), .A2(n_75), .B(n_76), .C(n_77), .Y(n_1006) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_826), .B(n_78), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g1008 ( .A1(n_816), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_1008) );
AOI21xp5_ASAP7_75t_L g1009 ( .A1(n_864), .A2(n_265), .B(n_264), .Y(n_1009) );
NAND2xp5_ASAP7_75t_SL g1010 ( .A(n_812), .B(n_79), .Y(n_1010) );
AO21x2_ASAP7_75t_L g1011 ( .A1(n_820), .A2(n_269), .B(n_266), .Y(n_1011) );
OAI21x1_ASAP7_75t_L g1012 ( .A1(n_867), .A2(n_272), .B(n_271), .Y(n_1012) );
INVx1_ASAP7_75t_SL g1013 ( .A(n_834), .Y(n_1013) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_824), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_806), .B(n_82), .Y(n_1015) );
BUFx3_ASAP7_75t_L g1016 ( .A(n_813), .Y(n_1016) );
AOI21xp5_ASAP7_75t_L g1017 ( .A1(n_810), .A2(n_275), .B(n_273), .Y(n_1017) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_874), .B(n_82), .Y(n_1018) );
AOI21xp5_ASAP7_75t_L g1019 ( .A1(n_808), .A2(n_282), .B(n_281), .Y(n_1019) );
A2O1A1Ixp33_ASAP7_75t_L g1020 ( .A1(n_837), .A2(n_83), .B(n_84), .C(n_85), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_830), .B(n_83), .Y(n_1021) );
NAND2x1p5_ASAP7_75t_L g1022 ( .A(n_891), .B(n_84), .Y(n_1022) );
AOI211x1_ASAP7_75t_L g1023 ( .A1(n_854), .A2(n_86), .B(n_87), .C(n_88), .Y(n_1023) );
OAI21x1_ASAP7_75t_L g1024 ( .A1(n_822), .A2(n_359), .B(n_358), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_894), .B(n_86), .Y(n_1025) );
AOI21x1_ASAP7_75t_L g1026 ( .A1(n_862), .A2(n_357), .B(n_356), .Y(n_1026) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_849), .A2(n_355), .B(n_354), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_811), .B(n_87), .Y(n_1028) );
INVx2_ASAP7_75t_L g1029 ( .A(n_866), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_895), .Y(n_1030) );
AOI21xp5_ASAP7_75t_L g1031 ( .A1(n_836), .A2(n_319), .B(n_349), .Y(n_1031) );
OAI21xp33_ASAP7_75t_SL g1032 ( .A1(n_859), .A2(n_89), .B(n_90), .Y(n_1032) );
O2A1O1Ixp33_ASAP7_75t_SL g1033 ( .A1(n_785), .A2(n_350), .B(n_347), .C(n_345), .Y(n_1033) );
AOI21x1_ASAP7_75t_L g1034 ( .A1(n_815), .A2(n_344), .B(n_343), .Y(n_1034) );
A2O1A1Ixp33_ASAP7_75t_L g1035 ( .A1(n_847), .A2(n_90), .B(n_91), .C(n_92), .Y(n_1035) );
NOR2xp33_ASAP7_75t_SL g1036 ( .A(n_784), .B(n_284), .Y(n_1036) );
A2O1A1Ixp33_ASAP7_75t_L g1037 ( .A1(n_847), .A2(n_91), .B(n_93), .C(n_94), .Y(n_1037) );
AO21x1_ASAP7_75t_L g1038 ( .A1(n_870), .A2(n_340), .B(n_339), .Y(n_1038) );
A2O1A1Ixp33_ASAP7_75t_L g1039 ( .A1(n_847), .A2(n_95), .B(n_96), .C(n_97), .Y(n_1039) );
NOR2xp67_ASAP7_75t_L g1040 ( .A(n_781), .B(n_285), .Y(n_1040) );
AOI21xp5_ASAP7_75t_L g1041 ( .A1(n_774), .A2(n_310), .B(n_335), .Y(n_1041) );
NOR2x1_ASAP7_75t_L g1042 ( .A(n_875), .B(n_95), .Y(n_1042) );
INVx2_ASAP7_75t_SL g1043 ( .A(n_883), .Y(n_1043) );
INVx1_ASAP7_75t_SL g1044 ( .A(n_766), .Y(n_1044) );
AO32x2_ASAP7_75t_L g1045 ( .A1(n_880), .A2(n_96), .A3(n_98), .B1(n_99), .B2(n_100), .Y(n_1045) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_883), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_859), .Y(n_1047) );
BUFx3_ASAP7_75t_L g1048 ( .A(n_883), .Y(n_1048) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_883), .Y(n_1049) );
AO31x2_ASAP7_75t_L g1050 ( .A1(n_767), .A2(n_99), .A3(n_100), .B(n_101), .Y(n_1050) );
INVx3_ASAP7_75t_L g1051 ( .A(n_875), .Y(n_1051) );
NOR2x1_ASAP7_75t_SL g1052 ( .A(n_835), .B(n_101), .Y(n_1052) );
AOI21xp5_ASAP7_75t_L g1053 ( .A1(n_774), .A2(n_328), .B(n_324), .Y(n_1053) );
INVx2_ASAP7_75t_L g1054 ( .A(n_848), .Y(n_1054) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_883), .Y(n_1055) );
NAND2xp5_ASAP7_75t_SL g1056 ( .A(n_795), .B(n_102), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_971), .B(n_102), .Y(n_1057) );
BUFx2_ASAP7_75t_SL g1058 ( .A(n_899), .Y(n_1058) );
OAI21xp5_ASAP7_75t_L g1059 ( .A1(n_898), .A2(n_103), .B(n_104), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1054), .Y(n_1060) );
AO21x2_ASAP7_75t_L g1061 ( .A1(n_923), .A2(n_308), .B(n_307), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_924), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_912), .B(n_104), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_952), .Y(n_1064) );
O2A1O1Ixp33_ASAP7_75t_L g1065 ( .A1(n_998), .A2(n_106), .B(n_107), .C(n_108), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_920), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_921), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_928), .Y(n_1068) );
OAI21xp5_ASAP7_75t_L g1069 ( .A1(n_905), .A2(n_106), .B(n_107), .Y(n_1069) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_952), .Y(n_1070) );
INVx2_ASAP7_75t_L g1071 ( .A(n_937), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_913), .B(n_109), .Y(n_1072) );
OAI21x1_ASAP7_75t_L g1073 ( .A1(n_1041), .A2(n_111), .B(n_112), .Y(n_1073) );
A2O1A1Ixp33_ASAP7_75t_L g1074 ( .A1(n_998), .A2(n_113), .B(n_114), .C(n_115), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_942), .Y(n_1075) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_903), .B(n_114), .Y(n_1076) );
AOI21xp5_ASAP7_75t_L g1077 ( .A1(n_902), .A2(n_117), .B(n_120), .Y(n_1077) );
NAND2x1p5_ASAP7_75t_L g1078 ( .A(n_952), .B(n_120), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_908), .B(n_121), .Y(n_1079) );
AO31x2_ASAP7_75t_L g1080 ( .A1(n_1038), .A2(n_121), .A3(n_122), .B(n_123), .Y(n_1080) );
OAI21x1_ASAP7_75t_L g1081 ( .A1(n_1053), .A2(n_123), .B(n_125), .Y(n_1081) );
BUFx2_ASAP7_75t_L g1082 ( .A(n_930), .Y(n_1082) );
AND2x4_ASAP7_75t_SL g1083 ( .A(n_1043), .B(n_126), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_919), .Y(n_1084) );
INVx3_ASAP7_75t_L g1085 ( .A(n_962), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_919), .Y(n_1086) );
AOI21xp5_ASAP7_75t_L g1087 ( .A1(n_1033), .A2(n_128), .B(n_130), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1047), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_1007), .Y(n_1089) );
BUFx8_ASAP7_75t_L g1090 ( .A(n_1046), .Y(n_1090) );
A2O1A1Ixp33_ASAP7_75t_L g1091 ( .A1(n_1032), .A2(n_131), .B(n_133), .C(n_135), .Y(n_1091) );
OA21x2_ASAP7_75t_L g1092 ( .A1(n_914), .A2(n_133), .B(n_136), .Y(n_1092) );
OAI21xp5_ASAP7_75t_L g1093 ( .A1(n_1032), .A2(n_136), .B(n_137), .Y(n_1093) );
NAND2x1p5_ASAP7_75t_L g1094 ( .A(n_962), .B(n_137), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_958), .B(n_138), .Y(n_1095) );
INVx2_ASAP7_75t_L g1096 ( .A(n_1050), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_925), .A2(n_138), .B1(n_139), .B2(n_140), .Y(n_1097) );
NOR2xp33_ASAP7_75t_L g1098 ( .A(n_985), .B(n_139), .Y(n_1098) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_1001), .B(n_944), .Y(n_1099) );
AO31x2_ASAP7_75t_L g1100 ( .A1(n_970), .A2(n_141), .A3(n_142), .B(n_143), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1050), .Y(n_1101) );
AOI21xp5_ASAP7_75t_L g1102 ( .A1(n_1021), .A2(n_141), .B(n_144), .Y(n_1102) );
AOI21xp5_ASAP7_75t_L g1103 ( .A1(n_1015), .A2(n_144), .B(n_145), .Y(n_1103) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_1003), .A2(n_146), .B(n_148), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_958), .B(n_150), .Y(n_1105) );
OAI21x1_ASAP7_75t_L g1106 ( .A1(n_1024), .A2(n_150), .B(n_151), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1050), .Y(n_1107) );
OAI21x1_ASAP7_75t_L g1108 ( .A1(n_945), .A2(n_153), .B(n_154), .Y(n_1108) );
OAI21x1_ASAP7_75t_L g1109 ( .A1(n_1034), .A2(n_153), .B(n_155), .Y(n_1109) );
AOI21xp5_ASAP7_75t_L g1110 ( .A1(n_922), .A2(n_155), .B(n_156), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_979), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_1014), .A2(n_157), .B1(n_158), .B2(n_159), .Y(n_1112) );
OAI21x1_ASAP7_75t_L g1113 ( .A1(n_981), .A2(n_157), .B(n_158), .Y(n_1113) );
AO21x2_ASAP7_75t_L g1114 ( .A1(n_934), .A2(n_161), .B(n_162), .Y(n_1114) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_939), .B(n_162), .Y(n_1115) );
OA21x2_ASAP7_75t_L g1116 ( .A1(n_927), .A2(n_929), .B(n_1012), .Y(n_1116) );
INVxp67_ASAP7_75t_SL g1117 ( .A(n_915), .Y(n_1117) );
OAI21x1_ASAP7_75t_L g1118 ( .A1(n_1009), .A2(n_948), .B(n_936), .Y(n_1118) );
AO21x2_ASAP7_75t_L g1119 ( .A1(n_934), .A2(n_957), .B(n_910), .Y(n_1119) );
AOI21xp5_ASAP7_75t_L g1120 ( .A1(n_938), .A2(n_947), .B(n_999), .Y(n_1120) );
OAI21xp5_ASAP7_75t_L g1121 ( .A1(n_977), .A2(n_951), .B(n_974), .Y(n_1121) );
OAI21x1_ASAP7_75t_L g1122 ( .A1(n_918), .A2(n_968), .B(n_966), .Y(n_1122) );
AOI21xp5_ASAP7_75t_L g1123 ( .A1(n_996), .A2(n_1029), .B(n_911), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_982), .B(n_1013), .Y(n_1124) );
AOI21xp5_ASAP7_75t_L g1125 ( .A1(n_1017), .A2(n_989), .B(n_1013), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_910), .A2(n_932), .B1(n_1008), .B2(n_995), .Y(n_1126) );
INVx1_ASAP7_75t_SL g1127 ( .A(n_980), .Y(n_1127) );
OAI21x1_ASAP7_75t_SL g1128 ( .A1(n_1052), .A2(n_933), .B(n_1042), .Y(n_1128) );
BUFx4f_ASAP7_75t_L g1129 ( .A(n_994), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1130 ( .A1(n_941), .A2(n_1002), .B(n_957), .Y(n_1130) );
NAND2xp33_ASAP7_75t_SL g1131 ( .A(n_900), .B(n_955), .Y(n_1131) );
AND2x4_ASAP7_75t_L g1132 ( .A(n_939), .B(n_1051), .Y(n_1132) );
AND2x4_ASAP7_75t_L g1133 ( .A(n_1051), .B(n_1048), .Y(n_1133) );
INVx2_ASAP7_75t_L g1134 ( .A(n_990), .Y(n_1134) );
NAND4xp25_ASAP7_75t_SL g1135 ( .A(n_916), .B(n_932), .C(n_929), .D(n_1008), .Y(n_1135) );
INVx1_ASAP7_75t_SL g1136 ( .A(n_980), .Y(n_1136) );
HB1xp67_ASAP7_75t_L g1137 ( .A(n_1007), .Y(n_1137) );
INVx2_ASAP7_75t_L g1138 ( .A(n_975), .Y(n_1138) );
BUFx3_ASAP7_75t_L g1139 ( .A(n_1049), .Y(n_1139) );
INVx3_ASAP7_75t_L g1140 ( .A(n_963), .Y(n_1140) );
OA21x2_ASAP7_75t_L g1141 ( .A1(n_983), .A2(n_991), .B(n_988), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1030), .B(n_959), .Y(n_1142) );
OAI21x1_ASAP7_75t_L g1143 ( .A1(n_940), .A2(n_965), .B(n_961), .Y(n_1143) );
INVx2_ASAP7_75t_SL g1144 ( .A(n_1055), .Y(n_1144) );
OA21x2_ASAP7_75t_L g1145 ( .A1(n_1000), .A2(n_1031), .B(n_993), .Y(n_1145) );
AND2x4_ASAP7_75t_L g1146 ( .A(n_1016), .B(n_963), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1042), .Y(n_1147) );
BUFx12f_ASAP7_75t_L g1148 ( .A(n_969), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_943), .Y(n_1149) );
OAI21xp5_ASAP7_75t_L g1150 ( .A1(n_933), .A2(n_993), .B(n_972), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1025), .B(n_896), .Y(n_1151) );
OAI21xp5_ASAP7_75t_L g1152 ( .A1(n_1006), .A2(n_1019), .B(n_1027), .Y(n_1152) );
INVx1_ASAP7_75t_L g1153 ( .A(n_955), .Y(n_1153) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_949), .A2(n_997), .B1(n_916), .B2(n_992), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_909), .B(n_1044), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_956), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_909), .B(n_1044), .Y(n_1157) );
NAND2x1p5_ASAP7_75t_L g1158 ( .A(n_956), .B(n_950), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_987), .Y(n_1159) );
AOI21xp5_ASAP7_75t_L g1160 ( .A1(n_941), .A2(n_976), .B(n_986), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_909), .B(n_1022), .Y(n_1161) );
AO21x2_ASAP7_75t_L g1162 ( .A1(n_986), .A2(n_1011), .B(n_1040), .Y(n_1162) );
O2A1O1Ixp33_ASAP7_75t_L g1163 ( .A1(n_926), .A2(n_1039), .B(n_1037), .C(n_1035), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1045), .Y(n_1164) );
BUFx12f_ASAP7_75t_L g1165 ( .A(n_1005), .Y(n_1165) );
AO21x2_ASAP7_75t_L g1166 ( .A1(n_1011), .A2(n_1040), .B(n_946), .Y(n_1166) );
HB1xp67_ASAP7_75t_SL g1167 ( .A(n_935), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1004), .B(n_953), .Y(n_1168) );
OAI21x1_ASAP7_75t_L g1169 ( .A1(n_964), .A2(n_976), .B(n_1026), .Y(n_1169) );
A2O1A1Ixp33_ASAP7_75t_L g1170 ( .A1(n_954), .A2(n_973), .B(n_978), .C(n_1020), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_978), .A2(n_967), .B1(n_1018), .B2(n_1023), .Y(n_1171) );
INVx4_ASAP7_75t_L g1172 ( .A(n_1004), .Y(n_1172) );
OAI21xp5_ASAP7_75t_L g1173 ( .A1(n_984), .A2(n_1010), .B(n_1056), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_1028), .A2(n_1036), .B1(n_901), .B2(n_1045), .Y(n_1174) );
A2O1A1Ixp33_ASAP7_75t_L g1175 ( .A1(n_901), .A2(n_1023), .B(n_917), .C(n_960), .Y(n_1175) );
OAI21x1_ASAP7_75t_L g1176 ( .A1(n_901), .A2(n_960), .B(n_917), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_960), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_917), .B(n_912), .Y(n_1178) );
BUFx8_ASAP7_75t_L g1179 ( .A(n_1043), .Y(n_1179) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_930), .Y(n_1180) );
BUFx6f_ASAP7_75t_L g1181 ( .A(n_990), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_925), .A2(n_780), .B1(n_809), .B2(n_764), .Y(n_1182) );
INVx3_ASAP7_75t_L g1183 ( .A(n_952), .Y(n_1183) );
A2O1A1Ixp33_ASAP7_75t_L g1184 ( .A1(n_998), .A2(n_1032), .B(n_933), .C(n_685), .Y(n_1184) );
A2O1A1Ixp33_ASAP7_75t_L g1185 ( .A1(n_998), .A2(n_958), .B(n_1032), .C(n_982), .Y(n_1185) );
AND2x4_ASAP7_75t_L g1186 ( .A(n_931), .B(n_912), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1054), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_907), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_907), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g1190 ( .A(n_990), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_907), .Y(n_1191) );
AO21x2_ASAP7_75t_L g1192 ( .A1(n_897), .A2(n_904), .B(n_771), .Y(n_1192) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1054), .Y(n_1193) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_952), .Y(n_1194) );
AOI21xp5_ASAP7_75t_L g1195 ( .A1(n_906), .A2(n_767), .B(n_771), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_907), .Y(n_1196) );
OR2x2_ASAP7_75t_L g1197 ( .A(n_971), .B(n_869), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_907), .Y(n_1198) );
AO21x2_ASAP7_75t_L g1199 ( .A1(n_897), .A2(n_904), .B(n_771), .Y(n_1199) );
AND2x4_ASAP7_75t_L g1200 ( .A(n_931), .B(n_912), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_907), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1066), .Y(n_1202) );
OR2x6_ASAP7_75t_L g1203 ( .A(n_1158), .B(n_1089), .Y(n_1203) );
INVx2_ASAP7_75t_SL g1204 ( .A(n_1129), .Y(n_1204) );
INVx4_ASAP7_75t_L g1205 ( .A(n_1129), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1067), .Y(n_1206) );
HB1xp67_ASAP7_75t_L g1207 ( .A(n_1089), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1068), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1076), .B(n_1197), .Y(n_1209) );
OA21x2_ASAP7_75t_L g1210 ( .A1(n_1160), .A2(n_1130), .B(n_1176), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1071), .Y(n_1211) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1117), .B(n_1082), .Y(n_1212) );
BUFx3_ASAP7_75t_L g1213 ( .A(n_1180), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1075), .Y(n_1214) );
INVx2_ASAP7_75t_L g1215 ( .A(n_1096), .Y(n_1215) );
BUFx2_ASAP7_75t_SL g1216 ( .A(n_1139), .Y(n_1216) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1101), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1188), .Y(n_1218) );
OR2x6_ASAP7_75t_L g1219 ( .A(n_1158), .B(n_1137), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1117), .B(n_1189), .Y(n_1220) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_1151), .B(n_1111), .Y(n_1221) );
INVx3_ASAP7_75t_L g1222 ( .A(n_1183), .Y(n_1222) );
INVxp67_ASAP7_75t_SL g1223 ( .A(n_1137), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1191), .Y(n_1224) );
AO21x2_ASAP7_75t_L g1225 ( .A1(n_1160), .A2(n_1130), .B(n_1195), .Y(n_1225) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1107), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1062), .Y(n_1227) );
OAI221xp5_ASAP7_75t_L g1228 ( .A1(n_1154), .A2(n_1151), .B1(n_1074), .B2(n_1185), .C(n_1182), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1196), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1198), .Y(n_1230) );
OAI21xp5_ASAP7_75t_L g1231 ( .A1(n_1170), .A2(n_1120), .B(n_1163), .Y(n_1231) );
INVx3_ASAP7_75t_L g1232 ( .A(n_1183), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1201), .Y(n_1233) );
OA21x2_ASAP7_75t_L g1234 ( .A1(n_1175), .A2(n_1161), .B(n_1177), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1098), .B(n_1072), .Y(n_1235) );
INVx2_ASAP7_75t_SL g1236 ( .A(n_1064), .Y(n_1236) );
NAND3xp33_ASAP7_75t_L g1237 ( .A(n_1131), .B(n_1074), .C(n_1159), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1098), .B(n_1186), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1088), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1063), .Y(n_1240) );
OAI21xp5_ASAP7_75t_L g1241 ( .A1(n_1170), .A2(n_1120), .B(n_1163), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1186), .B(n_1200), .Y(n_1242) );
AND2x4_ASAP7_75t_L g1243 ( .A(n_1153), .B(n_1156), .Y(n_1243) );
BUFx2_ASAP7_75t_L g1244 ( .A(n_1064), .Y(n_1244) );
AO21x1_ASAP7_75t_SL g1245 ( .A1(n_1093), .A2(n_1194), .B(n_1070), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1200), .B(n_1079), .Y(n_1246) );
OR2x6_ASAP7_75t_L g1247 ( .A(n_1078), .B(n_1115), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1057), .B(n_1060), .Y(n_1248) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1116), .Y(n_1249) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1187), .B(n_1193), .Y(n_1250) );
NAND2x1p5_ASAP7_75t_L g1251 ( .A(n_1115), .B(n_1146), .Y(n_1251) );
CKINVDCx20_ASAP7_75t_R g1252 ( .A(n_1090), .Y(n_1252) );
HB1xp67_ASAP7_75t_L g1253 ( .A(n_1155), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1149), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1095), .B(n_1105), .Y(n_1255) );
BUFx6f_ASAP7_75t_L g1256 ( .A(n_1181), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1094), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1084), .B(n_1086), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1094), .Y(n_1259) );
INVx2_ASAP7_75t_SL g1260 ( .A(n_1070), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_1126), .A2(n_1182), .B1(n_1184), .B2(n_1124), .Y(n_1261) );
HB1xp67_ASAP7_75t_L g1262 ( .A(n_1155), .Y(n_1262) );
INVx2_ASAP7_75t_SL g1263 ( .A(n_1194), .Y(n_1263) );
INVx2_ASAP7_75t_SL g1264 ( .A(n_1146), .Y(n_1264) );
INVx2_ASAP7_75t_SL g1265 ( .A(n_1179), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1078), .Y(n_1266) );
BUFx2_ASAP7_75t_L g1267 ( .A(n_1133), .Y(n_1267) );
INVxp67_ASAP7_75t_SL g1268 ( .A(n_1157), .Y(n_1268) );
BUFx6f_ASAP7_75t_L g1269 ( .A(n_1181), .Y(n_1269) );
AO21x2_ASAP7_75t_L g1270 ( .A1(n_1087), .A2(n_1157), .B(n_1178), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1099), .B(n_1083), .Y(n_1271) );
AO21x2_ASAP7_75t_L g1272 ( .A1(n_1178), .A2(n_1162), .B(n_1123), .Y(n_1272) );
AOI21xp5_ASAP7_75t_SL g1273 ( .A1(n_1065), .A2(n_1091), .B(n_1093), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1142), .Y(n_1274) );
AND2x4_ASAP7_75t_L g1275 ( .A(n_1140), .B(n_1132), .Y(n_1275) );
INVx3_ASAP7_75t_L g1276 ( .A(n_1140), .Y(n_1276) );
INVx2_ASAP7_75t_L g1277 ( .A(n_1192), .Y(n_1277) );
INVxp67_ASAP7_75t_SL g1278 ( .A(n_1174), .Y(n_1278) );
INVx2_ASAP7_75t_SL g1279 ( .A(n_1179), .Y(n_1279) );
INVx4_ASAP7_75t_L g1280 ( .A(n_1165), .Y(n_1280) );
CKINVDCx20_ASAP7_75t_R g1281 ( .A(n_1090), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g1282 ( .A(n_1127), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1085), .B(n_1172), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1147), .Y(n_1284) );
OAI21xp33_ASAP7_75t_L g1285 ( .A1(n_1091), .A2(n_1184), .B(n_1135), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1174), .B(n_1112), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1102), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1102), .Y(n_1288) );
INVx2_ASAP7_75t_L g1289 ( .A(n_1199), .Y(n_1289) );
OA21x2_ASAP7_75t_L g1290 ( .A1(n_1123), .A2(n_1169), .B(n_1164), .Y(n_1290) );
BUFx6f_ASAP7_75t_L g1291 ( .A(n_1181), .Y(n_1291) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1171), .B(n_1168), .Y(n_1292) );
INVx3_ASAP7_75t_L g1293 ( .A(n_1172), .Y(n_1293) );
INVx3_ASAP7_75t_L g1294 ( .A(n_1190), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1058), .B(n_1112), .Y(n_1295) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1199), .Y(n_1296) );
OAI21xp5_ASAP7_75t_L g1297 ( .A1(n_1059), .A2(n_1121), .B(n_1150), .Y(n_1297) );
OR2x6_ASAP7_75t_L g1298 ( .A(n_1128), .B(n_1065), .Y(n_1298) );
AO21x2_ASAP7_75t_L g1299 ( .A1(n_1162), .A2(n_1119), .B(n_1150), .Y(n_1299) );
AOI21xp5_ASAP7_75t_SL g1300 ( .A1(n_1104), .A2(n_1069), .B(n_1171), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1110), .Y(n_1301) );
INVxp67_ASAP7_75t_L g1302 ( .A(n_1127), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1144), .B(n_1136), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1110), .Y(n_1304) );
INVx2_ASAP7_75t_SL g1305 ( .A(n_1136), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1103), .B(n_1069), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1103), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1097), .B(n_1121), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1138), .B(n_1168), .Y(n_1309) );
BUFx2_ASAP7_75t_L g1310 ( .A(n_1148), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1097), .B(n_1100), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1077), .B(n_1104), .Y(n_1312) );
INVx2_ASAP7_75t_SL g1313 ( .A(n_1134), .Y(n_1313) );
OR2x6_ASAP7_75t_L g1314 ( .A(n_1077), .B(n_1106), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1113), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1316 ( .A(n_1212), .B(n_1080), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1292), .B(n_1080), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1292), .B(n_1080), .Y(n_1318) );
HB1xp67_ASAP7_75t_L g1319 ( .A(n_1244), .Y(n_1319) );
INVxp67_ASAP7_75t_SL g1320 ( .A(n_1220), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1278), .B(n_1114), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1202), .Y(n_1322) );
BUFx3_ASAP7_75t_L g1323 ( .A(n_1213), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_1228), .A2(n_1059), .B1(n_1152), .B2(n_1141), .Y(n_1324) );
INVx2_ASAP7_75t_SL g1325 ( .A(n_1236), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1206), .Y(n_1326) );
OAI22xp5_ASAP7_75t_SL g1327 ( .A1(n_1252), .A2(n_1167), .B1(n_1092), .B2(n_1141), .Y(n_1327) );
INVxp67_ASAP7_75t_L g1328 ( .A(n_1216), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1278), .B(n_1114), .Y(n_1329) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1215), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1227), .B(n_1119), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1231), .B(n_1166), .Y(n_1332) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_1221), .A2(n_1152), .B1(n_1145), .B2(n_1173), .Y(n_1333) );
AND2x4_ASAP7_75t_L g1334 ( .A(n_1298), .B(n_1166), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1217), .Y(n_1335) );
INVx3_ASAP7_75t_L g1336 ( .A(n_1256), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1241), .B(n_1145), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1282), .B(n_1073), .Y(n_1338) );
AND2x4_ASAP7_75t_L g1339 ( .A(n_1298), .B(n_1108), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1218), .Y(n_1340) );
NOR2x1_ASAP7_75t_SL g1341 ( .A(n_1247), .B(n_1061), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1342 ( .A(n_1282), .B(n_1081), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1226), .Y(n_1343) );
INVxp67_ASAP7_75t_SL g1344 ( .A(n_1223), .Y(n_1344) );
AND2x4_ASAP7_75t_L g1345 ( .A(n_1298), .B(n_1109), .Y(n_1345) );
OR2x6_ASAP7_75t_L g1346 ( .A(n_1247), .B(n_1125), .Y(n_1346) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1249), .Y(n_1347) );
BUFx2_ASAP7_75t_L g1348 ( .A(n_1247), .Y(n_1348) );
BUFx3_ASAP7_75t_L g1349 ( .A(n_1213), .Y(n_1349) );
BUFx3_ASAP7_75t_L g1350 ( .A(n_1251), .Y(n_1350) );
BUFx2_ASAP7_75t_L g1351 ( .A(n_1253), .Y(n_1351) );
INVx2_ASAP7_75t_SL g1352 ( .A(n_1260), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1224), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1229), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1230), .Y(n_1355) );
NOR2x1_ASAP7_75t_SL g1356 ( .A(n_1245), .B(n_1122), .Y(n_1356) );
INVxp67_ASAP7_75t_L g1357 ( .A(n_1263), .Y(n_1357) );
HB1xp67_ASAP7_75t_L g1358 ( .A(n_1263), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1233), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1274), .B(n_1118), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1254), .B(n_1143), .Y(n_1361) );
INVx4_ASAP7_75t_R g1362 ( .A(n_1265), .Y(n_1362) );
NOR3xp33_ASAP7_75t_L g1363 ( .A(n_1237), .B(n_1257), .C(n_1259), .Y(n_1363) );
NOR2x1_ASAP7_75t_SL g1364 ( .A(n_1203), .B(n_1219), .Y(n_1364) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_1205), .B(n_1280), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1285), .B(n_1297), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1284), .B(n_1208), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1211), .B(n_1214), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1261), .B(n_1239), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1309), .Y(n_1370) );
OR2x6_ASAP7_75t_L g1371 ( .A(n_1273), .B(n_1251), .Y(n_1371) );
BUFx6f_ASAP7_75t_L g1372 ( .A(n_1256), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1253), .B(n_1262), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1262), .B(n_1287), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1288), .B(n_1301), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1304), .B(n_1307), .Y(n_1376) );
INVx5_ASAP7_75t_SL g1377 ( .A(n_1203), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1234), .B(n_1268), .Y(n_1378) );
INVx1_ASAP7_75t_SL g1379 ( .A(n_1242), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1250), .Y(n_1380) );
AOI22xp5_ASAP7_75t_L g1381 ( .A1(n_1295), .A2(n_1235), .B1(n_1238), .B2(n_1308), .Y(n_1381) );
BUFx3_ASAP7_75t_L g1382 ( .A(n_1275), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1234), .B(n_1302), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1302), .B(n_1240), .Y(n_1384) );
BUFx2_ASAP7_75t_L g1385 ( .A(n_1223), .Y(n_1385) );
INVx2_ASAP7_75t_SL g1386 ( .A(n_1275), .Y(n_1386) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1207), .B(n_1209), .Y(n_1387) );
BUFx3_ASAP7_75t_L g1388 ( .A(n_1275), .Y(n_1388) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1305), .B(n_1255), .Y(n_1389) );
HB1xp67_ASAP7_75t_L g1390 ( .A(n_1303), .Y(n_1390) );
BUFx2_ASAP7_75t_L g1391 ( .A(n_1269), .Y(n_1391) );
INVx2_ASAP7_75t_SL g1392 ( .A(n_1264), .Y(n_1392) );
BUFx2_ASAP7_75t_L g1393 ( .A(n_1385), .Y(n_1393) );
INVx2_ASAP7_75t_L g1394 ( .A(n_1347), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1375), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1322), .Y(n_1396) );
OR2x2_ASAP7_75t_L g1397 ( .A(n_1387), .B(n_1286), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1337), .B(n_1270), .Y(n_1398) );
INVx3_ASAP7_75t_L g1399 ( .A(n_1339), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1332), .B(n_1299), .Y(n_1400) );
NAND2x1p5_ASAP7_75t_L g1401 ( .A(n_1348), .B(n_1266), .Y(n_1401) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_1328), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1326), .Y(n_1403) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_1385), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1332), .B(n_1299), .Y(n_1405) );
NAND2x1_ASAP7_75t_SL g1406 ( .A(n_1334), .B(n_1276), .Y(n_1406) );
BUFx2_ASAP7_75t_L g1407 ( .A(n_1344), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1374), .B(n_1277), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1374), .B(n_1289), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1317), .B(n_1289), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1340), .Y(n_1411) );
OAI21xp33_ASAP7_75t_L g1412 ( .A1(n_1366), .A2(n_1300), .B(n_1311), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1376), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1317), .B(n_1318), .Y(n_1414) );
OR2x2_ASAP7_75t_L g1415 ( .A(n_1387), .B(n_1296), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1353), .Y(n_1416) );
NAND2x1p5_ASAP7_75t_L g1417 ( .A(n_1348), .B(n_1276), .Y(n_1417) );
OR2x2_ASAP7_75t_L g1418 ( .A(n_1320), .B(n_1306), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1419 ( .A(n_1351), .B(n_1225), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1354), .Y(n_1420) );
AND2x4_ASAP7_75t_L g1421 ( .A(n_1339), .B(n_1315), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1383), .B(n_1290), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1383), .B(n_1290), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1376), .B(n_1290), .Y(n_1424) );
NAND2xp5_ASAP7_75t_SL g1425 ( .A(n_1325), .B(n_1265), .Y(n_1425) );
OR2x2_ASAP7_75t_L g1426 ( .A(n_1351), .B(n_1272), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1355), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1366), .B(n_1272), .Y(n_1428) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1359), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1321), .B(n_1210), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_1389), .B(n_1312), .Y(n_1431) );
NOR2xp33_ASAP7_75t_R g1432 ( .A(n_1365), .B(n_1281), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1321), .B(n_1210), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1380), .B(n_1264), .Y(n_1434) );
AND2x4_ASAP7_75t_L g1435 ( .A(n_1345), .B(n_1356), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1329), .B(n_1373), .Y(n_1436) );
INVx4_ASAP7_75t_L g1437 ( .A(n_1350), .Y(n_1437) );
BUFx2_ASAP7_75t_L g1438 ( .A(n_1323), .Y(n_1438) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1367), .Y(n_1439) );
NOR2xp67_ASAP7_75t_L g1440 ( .A(n_1319), .B(n_1279), .Y(n_1440) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1368), .Y(n_1441) );
NAND2xp5_ASAP7_75t_L g1442 ( .A(n_1368), .B(n_1246), .Y(n_1442) );
INVx1_ASAP7_75t_SL g1443 ( .A(n_1349), .Y(n_1443) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1384), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1384), .Y(n_1445) );
AND2x4_ASAP7_75t_L g1446 ( .A(n_1345), .B(n_1314), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1329), .B(n_1210), .Y(n_1447) );
OR2x2_ASAP7_75t_L g1448 ( .A(n_1389), .B(n_1248), .Y(n_1448) );
HB1xp67_ASAP7_75t_L g1449 ( .A(n_1358), .Y(n_1449) );
INVx3_ASAP7_75t_L g1450 ( .A(n_1345), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1396), .Y(n_1451) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1403), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1436), .B(n_1390), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1436), .B(n_1379), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1414), .B(n_1378), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1414), .B(n_1378), .Y(n_1456) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1411), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1416), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1420), .Y(n_1459) );
AOI22xp5_ASAP7_75t_L g1460 ( .A1(n_1440), .A2(n_1363), .B1(n_1369), .B2(n_1381), .Y(n_1460) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1427), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1429), .Y(n_1462) );
AND2x4_ASAP7_75t_L g1463 ( .A(n_1435), .B(n_1356), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1439), .B(n_1349), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1444), .B(n_1352), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1445), .B(n_1352), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1441), .B(n_1370), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1468 ( .A(n_1395), .B(n_1370), .Y(n_1468) );
HB1xp67_ASAP7_75t_L g1469 ( .A(n_1407), .Y(n_1469) );
OR2x2_ASAP7_75t_L g1470 ( .A(n_1418), .B(n_1316), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1471 ( .A(n_1448), .B(n_1316), .Y(n_1471) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1424), .Y(n_1472) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_1448), .B(n_1335), .Y(n_1473) );
AND2x4_ASAP7_75t_L g1474 ( .A(n_1435), .B(n_1346), .Y(n_1474) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1397), .B(n_1343), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1428), .B(n_1331), .Y(n_1476) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1413), .Y(n_1477) );
OR2x2_ASAP7_75t_L g1478 ( .A(n_1407), .B(n_1343), .Y(n_1478) );
NAND2x1_ASAP7_75t_L g1479 ( .A(n_1438), .B(n_1362), .Y(n_1479) );
AND2x4_ASAP7_75t_SL g1480 ( .A(n_1437), .B(n_1371), .Y(n_1480) );
AND2x4_ASAP7_75t_L g1481 ( .A(n_1435), .B(n_1346), .Y(n_1481) );
INVx2_ASAP7_75t_L g1482 ( .A(n_1424), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1428), .B(n_1331), .Y(n_1483) );
NOR2x1_ASAP7_75t_L g1484 ( .A(n_1425), .B(n_1252), .Y(n_1484) );
OR3x2_ASAP7_75t_L g1485 ( .A(n_1432), .B(n_1281), .C(n_1364), .Y(n_1485) );
INVx2_ASAP7_75t_L g1486 ( .A(n_1394), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1410), .B(n_1361), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_1449), .B(n_1357), .Y(n_1488) );
OR2x2_ASAP7_75t_L g1489 ( .A(n_1431), .B(n_1330), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1443), .B(n_1386), .Y(n_1490) );
AOI22xp5_ASAP7_75t_L g1491 ( .A1(n_1412), .A2(n_1371), .B1(n_1327), .B2(n_1386), .Y(n_1491) );
INVxp67_ASAP7_75t_L g1492 ( .A(n_1393), .Y(n_1492) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_1431), .B(n_1330), .Y(n_1493) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_1485), .A2(n_1371), .B1(n_1446), .B2(n_1405), .Y(n_1494) );
INVx2_ASAP7_75t_L g1495 ( .A(n_1486), .Y(n_1495) );
AO21x1_ASAP7_75t_L g1496 ( .A1(n_1479), .A2(n_1437), .B(n_1401), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1472), .B(n_1426), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1472), .B(n_1400), .Y(n_1498) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1451), .Y(n_1499) );
NAND2x1_ASAP7_75t_SL g1500 ( .A(n_1463), .B(n_1485), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1452), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1482), .B(n_1430), .Y(n_1502) );
INVxp67_ASAP7_75t_L g1503 ( .A(n_1469), .Y(n_1503) );
INVxp67_ASAP7_75t_SL g1504 ( .A(n_1469), .Y(n_1504) );
OR2x2_ASAP7_75t_L g1505 ( .A(n_1482), .B(n_1426), .Y(n_1505) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1486), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1455), .B(n_1430), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1508 ( .A(n_1470), .B(n_1419), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1455), .B(n_1433), .Y(n_1509) );
HB1xp67_ASAP7_75t_L g1510 ( .A(n_1492), .Y(n_1510) );
OAI22xp5_ASAP7_75t_L g1511 ( .A1(n_1460), .A2(n_1377), .B1(n_1401), .B2(n_1402), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1456), .B(n_1433), .Y(n_1512) );
OR2x2_ASAP7_75t_L g1513 ( .A(n_1471), .B(n_1415), .Y(n_1513) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1457), .Y(n_1514) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1458), .Y(n_1515) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1459), .Y(n_1516) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1461), .Y(n_1517) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1462), .Y(n_1518) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1477), .Y(n_1519) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1473), .Y(n_1520) );
INVx1_ASAP7_75t_SL g1521 ( .A(n_1513), .Y(n_1521) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1497), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1507), .B(n_1454), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1507), .B(n_1453), .Y(n_1524) );
AOI31xp33_ASAP7_75t_L g1525 ( .A1(n_1496), .A2(n_1484), .A3(n_1511), .B(n_1402), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1509), .B(n_1476), .Y(n_1526) );
OAI22xp33_ASAP7_75t_SL g1527 ( .A1(n_1504), .A2(n_1488), .B1(n_1492), .B2(n_1463), .Y(n_1527) );
OAI21xp33_ASAP7_75t_L g1528 ( .A1(n_1500), .A2(n_1491), .B(n_1483), .Y(n_1528) );
NAND2xp5_ASAP7_75t_SL g1529 ( .A(n_1503), .B(n_1463), .Y(n_1529) );
OAI32xp33_ASAP7_75t_L g1530 ( .A1(n_1510), .A2(n_1401), .A3(n_1417), .B1(n_1478), .B2(n_1442), .Y(n_1530) );
INVx3_ASAP7_75t_L g1531 ( .A(n_1495), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_1494), .A2(n_1480), .B1(n_1474), .B2(n_1481), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1499), .Y(n_1533) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1501), .Y(n_1534) );
NAND2xp5_ASAP7_75t_L g1535 ( .A(n_1520), .B(n_1476), .Y(n_1535) );
INVxp67_ASAP7_75t_SL g1536 ( .A(n_1500), .Y(n_1536) );
NOR2xp33_ASAP7_75t_R g1537 ( .A(n_1521), .B(n_1310), .Y(n_1537) );
AOI21xp5_ASAP7_75t_L g1538 ( .A1(n_1525), .A2(n_1364), .B(n_1474), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_1536), .A2(n_1508), .B1(n_1512), .B2(n_1474), .Y(n_1539) );
INVx1_ASAP7_75t_SL g1540 ( .A(n_1523), .Y(n_1540) );
OAI21xp33_ASAP7_75t_L g1541 ( .A1(n_1527), .A2(n_1505), .B(n_1497), .Y(n_1541) );
AOI21xp5_ASAP7_75t_L g1542 ( .A1(n_1529), .A2(n_1481), .B(n_1490), .Y(n_1542) );
OAI221xp5_ASAP7_75t_L g1543 ( .A1(n_1532), .A2(n_1505), .B1(n_1516), .B2(n_1518), .C(n_1517), .Y(n_1543) );
OAI32xp33_ASAP7_75t_L g1544 ( .A1(n_1529), .A2(n_1417), .A3(n_1515), .B1(n_1514), .B2(n_1475), .Y(n_1544) );
AOI22xp33_ASAP7_75t_L g1545 ( .A1(n_1522), .A2(n_1446), .B1(n_1481), .B2(n_1450), .Y(n_1545) );
AOI221xp5_ASAP7_75t_L g1546 ( .A1(n_1530), .A2(n_1519), .B1(n_1498), .B2(n_1502), .C(n_1467), .Y(n_1546) );
OAI22xp33_ASAP7_75t_L g1547 ( .A1(n_1524), .A2(n_1404), .B1(n_1393), .B2(n_1417), .Y(n_1547) );
INVxp67_ASAP7_75t_L g1548 ( .A(n_1533), .Y(n_1548) );
AOI21xp5_ASAP7_75t_L g1549 ( .A1(n_1530), .A2(n_1468), .B(n_1404), .Y(n_1549) );
AOI221xp5_ASAP7_75t_L g1550 ( .A1(n_1534), .A2(n_1464), .B1(n_1466), .B2(n_1465), .C(n_1483), .Y(n_1550) );
NAND4xp25_ASAP7_75t_L g1551 ( .A(n_1535), .B(n_1271), .C(n_1324), .D(n_1434), .Y(n_1551) );
NAND3xp33_ASAP7_75t_SL g1552 ( .A(n_1526), .B(n_1333), .C(n_1267), .Y(n_1552) );
AOI221xp5_ASAP7_75t_L g1553 ( .A1(n_1526), .A2(n_1487), .B1(n_1506), .B2(n_1398), .C(n_1450), .Y(n_1553) );
O2A1O1Ixp33_ASAP7_75t_L g1554 ( .A1(n_1531), .A2(n_1204), .B(n_1346), .C(n_1392), .Y(n_1554) );
AOI22xp33_ASAP7_75t_SL g1555 ( .A1(n_1531), .A2(n_1399), .B1(n_1446), .B2(n_1377), .Y(n_1555) );
NOR3xp33_ASAP7_75t_L g1556 ( .A(n_1525), .B(n_1204), .C(n_1232), .Y(n_1556) );
AOI322xp5_ASAP7_75t_L g1557 ( .A1(n_1528), .A2(n_1447), .A3(n_1422), .B1(n_1423), .B2(n_1410), .C1(n_1409), .C2(n_1408), .Y(n_1557) );
NAND4xp25_ASAP7_75t_L g1558 ( .A(n_1556), .B(n_1538), .C(n_1557), .D(n_1546), .Y(n_1558) );
NAND4xp25_ASAP7_75t_SL g1559 ( .A(n_1543), .B(n_1542), .C(n_1553), .D(n_1545), .Y(n_1559) );
NAND3xp33_ASAP7_75t_SL g1560 ( .A(n_1537), .B(n_1541), .C(n_1549), .Y(n_1560) );
OAI211xp5_ASAP7_75t_L g1561 ( .A1(n_1552), .A2(n_1544), .B(n_1551), .C(n_1555), .Y(n_1561) );
NOR2x1_ASAP7_75t_L g1562 ( .A(n_1539), .B(n_1547), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1562), .B(n_1540), .Y(n_1563) );
NOR3xp33_ASAP7_75t_L g1564 ( .A(n_1560), .B(n_1554), .C(n_1548), .Y(n_1564) );
NOR3xp33_ASAP7_75t_L g1565 ( .A(n_1561), .B(n_1550), .C(n_1222), .Y(n_1565) );
OAI221xp5_ASAP7_75t_SL g1566 ( .A1(n_1558), .A2(n_1203), .B1(n_1219), .B2(n_1493), .C(n_1489), .Y(n_1566) );
NOR4xp25_ASAP7_75t_L g1567 ( .A(n_1559), .B(n_1258), .C(n_1293), .D(n_1283), .Y(n_1567) );
INVx2_ASAP7_75t_SL g1568 ( .A(n_1563), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1564), .Y(n_1569) );
XNOR2x1_ASAP7_75t_L g1570 ( .A(n_1567), .B(n_1243), .Y(n_1570) );
INVx2_ASAP7_75t_SL g1571 ( .A(n_1566), .Y(n_1571) );
NOR3xp33_ASAP7_75t_L g1572 ( .A(n_1569), .B(n_1571), .C(n_1568), .Y(n_1572) );
XOR2xp5_ASAP7_75t_L g1573 ( .A(n_1570), .B(n_1565), .Y(n_1573) );
AND3x2_ASAP7_75t_L g1574 ( .A(n_1572), .B(n_1243), .C(n_1391), .Y(n_1574) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_1573), .A2(n_1421), .B1(n_1388), .B2(n_1382), .Y(n_1575) );
XNOR2x1_ASAP7_75t_SL g1576 ( .A(n_1574), .B(n_1294), .Y(n_1576) );
OAI22xp5_ASAP7_75t_L g1577 ( .A1(n_1575), .A2(n_1388), .B1(n_1415), .B2(n_1338), .Y(n_1577) );
OAI21xp5_ASAP7_75t_SL g1578 ( .A1(n_1577), .A2(n_1391), .B(n_1336), .Y(n_1578) );
NOR2xp67_ASAP7_75t_L g1579 ( .A(n_1576), .B(n_1342), .Y(n_1579) );
OAI21xp5_ASAP7_75t_L g1580 ( .A1(n_1579), .A2(n_1406), .B(n_1360), .Y(n_1580) );
AOI21xp5_ASAP7_75t_L g1581 ( .A1(n_1578), .A2(n_1341), .B(n_1314), .Y(n_1581) );
OAI22xp33_ASAP7_75t_L g1582 ( .A1(n_1580), .A2(n_1269), .B1(n_1291), .B2(n_1372), .Y(n_1582) );
AOI21xp5_ASAP7_75t_L g1583 ( .A1(n_1582), .A2(n_1581), .B(n_1313), .Y(n_1583) );
endmodule