module fake_netlist_6_3707_n_85 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_85);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_85;

wire n_52;
wire n_46;
wire n_21;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_77;
wire n_42;
wire n_24;
wire n_54;
wire n_32;
wire n_66;
wire n_78;
wire n_84;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_80;
wire n_41;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_2),
.A2(n_15),
.B1(n_3),
.B2(n_10),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_2),
.Y(n_22)
);

AND2x4_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_15),
.Y(n_27)
);

AND2x4_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_11),
.A2(n_12),
.B1(n_9),
.B2(n_5),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_0),
.B1(n_8),
.B2(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_14),
.B1(n_13),
.B2(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_21),
.A2(n_5),
.B1(n_10),
.B2(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_23),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_20),
.B1(n_31),
.B2(n_29),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_27),
.B(n_24),
.C(n_33),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_26),
.B(n_33),
.C(n_22),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_20),
.B(n_26),
.Y(n_46)
);

AO21x2_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_23),
.B(n_31),
.Y(n_47)
);

NOR2x1_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_43),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_23),
.Y(n_57)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_34),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_56),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_47),
.B1(n_53),
.B2(n_52),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_57),
.B(n_52),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_53),
.B1(n_42),
.B2(n_58),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_53),
.B(n_58),
.Y(n_72)
);

AOI222xp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.C1(n_58),
.C2(n_42),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_34),
.C(n_30),
.Y(n_74)
);

NAND5xp2_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_32),
.C(n_72),
.D(n_71),
.E(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR4xp25_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_42),
.C(n_45),
.D(n_43),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_45),
.C(n_31),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_78),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_77),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_74),
.B(n_82),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_75),
.B(n_80),
.Y(n_85)
);


endmodule