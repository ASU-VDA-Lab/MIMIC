module fake_jpeg_8492_n_178 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_35),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_0),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_39),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_16),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_29),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_27),
.B1(n_19),
.B2(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_53),
.B1(n_20),
.B2(n_24),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_19),
.B1(n_27),
.B2(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_19),
.Y(n_59)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_34),
.B1(n_41),
.B2(n_37),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_66),
.B1(n_18),
.B2(n_30),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_17),
.B1(n_23),
.B2(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_79),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_23),
.B(n_20),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_6),
.C(n_7),
.Y(n_92)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_9),
.Y(n_95)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_15),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_25),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_24),
.B(n_25),
.C(n_18),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_81),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_26),
.Y(n_83)
);

OA21x2_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_84),
.B(n_92),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_1),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_88),
.B1(n_70),
.B2(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_2),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_5),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_101),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_6),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_66),
.C(n_68),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_9),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_106),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_71),
.B1(n_69),
.B2(n_60),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_116),
.B1(n_105),
.B2(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_110),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_57),
.C(n_75),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_93),
.C(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_79),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_88),
.B1(n_87),
.B2(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_81),
.B1(n_98),
.B2(n_74),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_94),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_56),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_85),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_82),
.B(n_90),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_135),
.B(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_128),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_133),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_101),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_89),
.B(n_92),
.C(n_99),
.D(n_84),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_99),
.B(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_98),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_108),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_155)
);

OAI322xp33_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_142),
.A3(n_122),
.B1(n_125),
.B2(n_136),
.C1(n_131),
.C2(n_130),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_107),
.C(n_117),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_110),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_106),
.C(n_109),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_144),
.A2(n_123),
.B(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_131),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_95),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_148),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_12),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_153),
.Y(n_164)
);

OA21x2_ASAP7_75t_SL g153 ( 
.A1(n_147),
.A2(n_123),
.B(n_132),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_143),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_138),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_130),
.B(n_7),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_78),
.B1(n_7),
.B2(n_8),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_14),
.B(n_6),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_161),
.B(n_151),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_145),
.B(n_137),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_151),
.B(n_150),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_12),
.C(n_14),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_157),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_167),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_162),
.C(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_164),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_174),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_172),
.B(n_173),
.C(n_158),
.Y(n_177)
);


endmodule