module fake_jpeg_17080_n_305 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_51;
wire n_47;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_13;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_21),
.B1(n_16),
.B2(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_48),
.B1(n_30),
.B2(n_21),
.Y(n_53)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_50),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_15),
.B(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_21),
.B1(n_27),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_58),
.B1(n_66),
.B2(n_48),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_33),
.B(n_20),
.C(n_32),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_35),
.B1(n_32),
.B2(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_16),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_23),
.B(n_14),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_64),
.B1(n_39),
.B2(n_46),
.Y(n_71)
);

AOI22x1_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_35),
.B1(n_28),
.B2(n_18),
.Y(n_64)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_31),
.B1(n_15),
.B2(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_18),
.B1(n_17),
.B2(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_36),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_71),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_39),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_59),
.B1(n_65),
.B2(n_56),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_84),
.B1(n_88),
.B2(n_48),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_80),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_77),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_39),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_48),
.B1(n_44),
.B2(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_99),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_93),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_64),
.B1(n_61),
.B2(n_50),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_101),
.B1(n_102),
.B2(n_107),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_109),
.B(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_51),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_54),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_68),
.B1(n_67),
.B2(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_68),
.B1(n_67),
.B2(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_65),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_65),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_79),
.B1(n_88),
.B2(n_74),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_69),
.B1(n_76),
.B2(n_71),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_121),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_92),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_99),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_106),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_75),
.C(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_125),
.B(n_128),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_94),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_74),
.B(n_79),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_103),
.B(n_109),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_131),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_86),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_103),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_144),
.C(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_126),
.B(n_114),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_96),
.CI(n_102),
.CON(n_143),
.SN(n_143)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_143),
.B(n_145),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_86),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_105),
.C(n_78),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_109),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_105),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_114),
.B(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_72),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_122),
.B(n_97),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_147),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_159),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_78),
.C(n_71),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_97),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_169),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_134),
.B1(n_130),
.B2(n_113),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_187),
.B1(n_152),
.B2(n_137),
.Y(n_195)
);

NAND4xp25_ASAP7_75t_SL g171 ( 
.A(n_158),
.B(n_116),
.C(n_120),
.D(n_44),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_97),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_126),
.B(n_69),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_173),
.A2(n_153),
.B(n_146),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_113),
.B1(n_120),
.B2(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_117),
.B1(n_69),
.B2(n_97),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_136),
.Y(n_181)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_142),
.C(n_138),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_72),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_141),
.A2(n_87),
.B1(n_44),
.B2(n_58),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_188),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_149),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_206),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_148),
.C(n_162),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_7),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_177),
.B1(n_175),
.B2(n_168),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_186),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_208),
.B(n_209),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_139),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_207),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_156),
.B(n_143),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_165),
.B(n_187),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_144),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_137),
.B(n_150),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_210),
.A2(n_176),
.B(n_202),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_229),
.B(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_167),
.C(n_178),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_219),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_170),
.B1(n_184),
.B2(n_178),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_231),
.B1(n_227),
.B2(n_222),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_177),
.C(n_168),
.Y(n_219)
);

AOI22x1_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_182),
.B1(n_179),
.B2(n_163),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_10),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_195),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_181),
.C(n_165),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_228),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_66),
.C(n_47),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_227),
.B(n_228),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_66),
.C(n_47),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_25),
.B(n_23),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_47),
.C(n_46),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_0),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_204),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_243),
.B(n_8),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_245),
.C(n_247),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_224),
.A2(n_198),
.B1(n_192),
.B2(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_212),
.B(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

AOI322xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_198),
.A3(n_211),
.B1(n_189),
.B2(n_200),
.C1(n_47),
.C2(n_44),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_240),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_242),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_25),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_12),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_17),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_222),
.B(n_215),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_215),
.C(n_18),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_251),
.C(n_256),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_17),
.C(n_18),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_23),
.B1(n_14),
.B2(n_12),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_8),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_7),
.Y(n_274)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_24),
.C(n_19),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_24),
.C(n_19),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_241),
.C(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_236),
.C(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_24),
.C(n_19),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_13),
.C(n_6),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_262),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_272),
.A2(n_262),
.B1(n_251),
.B2(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_13),
.C(n_7),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_257),
.C(n_256),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_5),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_277),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_279),
.B(n_283),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_281),
.C(n_282),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_13),
.C(n_4),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_269),
.B(n_4),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_280),
.C(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_R g286 ( 
.A(n_279),
.B(n_274),
.C(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_288),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_284),
.A2(n_271),
.B(n_4),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_3),
.B(n_5),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_0),
.C(n_1),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_5),
.C(n_8),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_292),
.B(n_287),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_295),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_297),
.B(n_9),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_0),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_1),
.C(n_2),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_1),
.B(n_9),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_9),
.B(n_1),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_1),
.Y(n_305)
);


endmodule