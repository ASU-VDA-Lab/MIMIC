module real_aes_1398_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_0), .B(n_120), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_1), .A2(n_129), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_2), .B(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_3), .B(n_120), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_4), .B(n_136), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_5), .B(n_136), .Y(n_506) );
INVx1_ASAP7_75t_L g127 ( .A(n_6), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_7), .B(n_136), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g763 ( .A(n_8), .Y(n_763) );
NAND2xp33_ASAP7_75t_L g487 ( .A(n_9), .B(n_138), .Y(n_487) );
AND2x2_ASAP7_75t_L g156 ( .A(n_10), .B(n_145), .Y(n_156) );
AND2x2_ASAP7_75t_L g165 ( .A(n_11), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
AOI221x1_ASAP7_75t_L g528 ( .A1(n_13), .A2(n_24), .B1(n_120), .B2(n_129), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_14), .B(n_136), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_15), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_16), .B(n_120), .Y(n_483) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_17), .A2(n_145), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_18), .B(n_140), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_19), .B(n_136), .Y(n_466) );
AO21x1_ASAP7_75t_L g501 ( .A1(n_20), .A2(n_120), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_21), .B(n_120), .Y(n_190) );
INVx1_ASAP7_75t_L g453 ( .A(n_22), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_23), .A2(n_91), .B1(n_120), .B2(n_229), .Y(n_228) );
NAND2x1_ASAP7_75t_L g515 ( .A(n_25), .B(n_136), .Y(n_515) );
NAND2x1_ASAP7_75t_L g476 ( .A(n_26), .B(n_138), .Y(n_476) );
OR2x2_ASAP7_75t_L g143 ( .A(n_27), .B(n_88), .Y(n_143) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_27), .A2(n_88), .B(n_142), .Y(n_146) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_28), .A2(n_103), .B1(n_756), .B2(n_767), .C1(n_785), .C2(n_789), .Y(n_102) );
OAI22x1_ASAP7_75t_R g775 ( .A1(n_28), .A2(n_776), .B1(n_777), .B2(n_780), .Y(n_775) );
INVx1_ASAP7_75t_L g780 ( .A(n_28), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_29), .B(n_138), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_30), .B(n_136), .Y(n_486) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_31), .A2(n_166), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_32), .B(n_138), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_33), .A2(n_129), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_34), .B(n_136), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_35), .A2(n_129), .B(n_547), .Y(n_546) );
XNOR2x2_ASAP7_75t_SL g104 ( .A(n_36), .B(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g126 ( .A(n_37), .B(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g130 ( .A(n_37), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g237 ( .A(n_37), .Y(n_237) );
OR2x6_ASAP7_75t_L g451 ( .A(n_38), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_39), .B(n_120), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_40), .B(n_120), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_41), .B(n_136), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_42), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_43), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_44), .B(n_138), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_45), .B(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_46), .A2(n_129), .B(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_47), .A2(n_129), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_48), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_49), .B(n_138), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_50), .B(n_120), .Y(n_172) );
INVx1_ASAP7_75t_L g123 ( .A(n_51), .Y(n_123) );
INVx1_ASAP7_75t_L g133 ( .A(n_51), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_52), .A2(n_68), .B1(n_778), .B2(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_52), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_53), .B(n_136), .Y(n_163) );
AND2x2_ASAP7_75t_L g201 ( .A(n_54), .B(n_140), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_55), .B(n_138), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_56), .B(n_136), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_57), .B(n_138), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_58), .A2(n_129), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_59), .B(n_120), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_60), .B(n_120), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_61), .A2(n_129), .B(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g196 ( .A(n_62), .B(n_141), .Y(n_196) );
AO21x1_ASAP7_75t_L g503 ( .A1(n_63), .A2(n_129), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_64), .B(n_120), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_65), .A2(n_82), .B1(n_106), .B2(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_65), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_66), .B(n_138), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_67), .B(n_120), .Y(n_478) );
INVx1_ASAP7_75t_L g779 ( .A(n_68), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_69), .B(n_138), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_70), .A2(n_96), .B1(n_129), .B2(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_71), .B(n_136), .Y(n_193) );
AND2x2_ASAP7_75t_L g551 ( .A(n_72), .B(n_141), .Y(n_551) );
INVx1_ASAP7_75t_L g125 ( .A(n_73), .Y(n_125) );
INVx1_ASAP7_75t_L g131 ( .A(n_73), .Y(n_131) );
AND2x2_ASAP7_75t_L g479 ( .A(n_74), .B(n_166), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_75), .B(n_138), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_76), .A2(n_129), .B(n_205), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_77), .A2(n_129), .B(n_134), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_78), .A2(n_129), .B(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g187 ( .A(n_79), .B(n_141), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_80), .B(n_140), .Y(n_226) );
INVx1_ASAP7_75t_L g454 ( .A(n_81), .Y(n_454) );
INVx1_ASAP7_75t_L g107 ( .A(n_82), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_83), .B(n_120), .Y(n_468) );
AND2x2_ASAP7_75t_L g489 ( .A(n_84), .B(n_166), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_85), .A2(n_104), .B1(n_748), .B2(n_752), .Y(n_747) );
AND2x2_ASAP7_75t_L g144 ( .A(n_86), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g502 ( .A(n_87), .B(n_177), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_89), .B(n_138), .Y(n_467) );
AND2x2_ASAP7_75t_L g518 ( .A(n_90), .B(n_166), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_92), .B(n_136), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_93), .A2(n_129), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_94), .B(n_138), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_95), .A2(n_129), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_97), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_98), .B(n_136), .Y(n_494) );
BUFx2_ASAP7_75t_L g195 ( .A(n_99), .Y(n_195) );
BUFx2_ASAP7_75t_L g764 ( .A(n_100), .Y(n_764) );
BUFx2_ASAP7_75t_SL g793 ( .A(n_100), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_101), .A2(n_129), .B(n_485), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_108), .B(n_747), .Y(n_103) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OAI22xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_446), .B1(n_455), .B2(n_745), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_111), .A2(n_448), .B1(n_749), .B2(n_750), .Y(n_748) );
OAI22x1_ASAP7_75t_SL g772 ( .A1(n_111), .A2(n_773), .B1(n_774), .B2(n_775), .Y(n_772) );
INVx5_ASAP7_75t_L g773 ( .A(n_111), .Y(n_773) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_350), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_275), .C(n_311), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_249), .Y(n_113) );
AOI211xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_167), .B(n_197), .C(n_222), .Y(n_114) );
AND2x2_ASAP7_75t_L g340 ( .A(n_115), .B(n_199), .Y(n_340) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_147), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_116), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g373 ( .A(n_116), .B(n_255), .Y(n_373) );
AND2x2_ASAP7_75t_L g389 ( .A(n_116), .B(n_214), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_116), .B(n_399), .Y(n_398) );
NAND2x1p5_ASAP7_75t_L g422 ( .A(n_116), .B(n_423), .Y(n_422) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_SL g209 ( .A(n_117), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g244 ( .A(n_117), .Y(n_244) );
AND2x2_ASAP7_75t_L g291 ( .A(n_117), .B(n_224), .Y(n_291) );
AND2x2_ASAP7_75t_L g310 ( .A(n_117), .B(n_147), .Y(n_310) );
BUFx2_ASAP7_75t_L g315 ( .A(n_117), .Y(n_315) );
AND2x2_ASAP7_75t_L g359 ( .A(n_117), .B(n_157), .Y(n_359) );
AND2x4_ASAP7_75t_L g431 ( .A(n_117), .B(n_432), .Y(n_431) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_117), .B(n_213), .Y(n_443) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_144), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_128), .B(n_140), .Y(n_118) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_126), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
AND2x6_ASAP7_75t_L g138 ( .A(n_122), .B(n_131), .Y(n_138) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g136 ( .A(n_124), .B(n_133), .Y(n_136) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx5_ASAP7_75t_L g139 ( .A(n_126), .Y(n_139) );
AND2x2_ASAP7_75t_L g132 ( .A(n_127), .B(n_133), .Y(n_132) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_127), .Y(n_232) );
AND2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
BUFx3_ASAP7_75t_L g233 ( .A(n_130), .Y(n_233) );
INVx2_ASAP7_75t_L g239 ( .A(n_131), .Y(n_239) );
AND2x4_ASAP7_75t_L g235 ( .A(n_132), .B(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g231 ( .A(n_133), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_137), .B(n_139), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_138), .B(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_139), .A2(n_153), .B(n_154), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_139), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_139), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_139), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_139), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_139), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_139), .A2(n_466), .B(n_467), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_139), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_139), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_139), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_139), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_139), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_139), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_139), .A2(n_548), .B(n_549), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_140), .Y(n_149) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_140), .A2(n_228), .B(n_234), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_140), .A2(n_491), .B(n_492), .Y(n_490) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_140), .A2(n_528), .B(n_532), .Y(n_527) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_140), .A2(n_528), .B(n_532), .Y(n_539) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x4_ASAP7_75t_L g177 ( .A(n_142), .B(n_143), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_145), .A2(n_190), .B(n_191), .Y(n_189) );
BUFx4f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_147), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g362 ( .A(n_147), .Y(n_362) );
BUFx2_ASAP7_75t_L g411 ( .A(n_147), .Y(n_411) );
INVx1_ASAP7_75t_L g433 ( .A(n_147), .Y(n_433) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_157), .Y(n_147) );
INVx3_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_148), .Y(n_399) );
AOI21x1_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_156), .Y(n_148) );
AO21x2_ASAP7_75t_L g472 ( .A1(n_149), .A2(n_473), .B(n_479), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
INVx2_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_157), .B(n_210), .Y(n_214) );
INVx2_ASAP7_75t_L g299 ( .A(n_157), .Y(n_299) );
OR2x2_ASAP7_75t_L g306 ( .A(n_157), .B(n_255), .Y(n_306) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_165), .Y(n_157) );
INVx4_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
INVx3_ASAP7_75t_L g180 ( .A(n_166), .Y(n_180) );
AND2x2_ASAP7_75t_L g261 ( .A(n_167), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g295 ( .A(n_167), .B(n_258), .Y(n_295) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_178), .Y(n_167) );
AND2x2_ASAP7_75t_L g331 ( .A(n_168), .B(n_220), .Y(n_331) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g288 ( .A(n_169), .B(n_179), .Y(n_288) );
AND2x2_ASAP7_75t_L g407 ( .A(n_169), .B(n_188), .Y(n_407) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
INVx1_ASAP7_75t_L g247 ( .A(n_170), .Y(n_247) );
AND2x2_ASAP7_75t_L g303 ( .A(n_170), .B(n_179), .Y(n_303) );
AND2x2_ASAP7_75t_L g308 ( .A(n_170), .B(n_200), .Y(n_308) );
OR2x2_ASAP7_75t_L g371 ( .A(n_170), .B(n_188), .Y(n_371) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_170), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_177), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_177), .A2(n_203), .B(n_204), .Y(n_202) );
INVx1_ASAP7_75t_SL g462 ( .A(n_177), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_177), .A2(n_483), .B(n_484), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_177), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g199 ( .A(n_178), .B(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g248 ( .A(n_178), .Y(n_248) );
NOR2x1_ASAP7_75t_SL g178 ( .A(n_179), .B(n_188), .Y(n_178) );
AO21x1_ASAP7_75t_SL g179 ( .A1(n_180), .A2(n_181), .B(n_187), .Y(n_179) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_180), .A2(n_181), .B(n_187), .Y(n_221) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_180), .A2(n_512), .B(n_518), .Y(n_511) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_180), .A2(n_545), .B(n_551), .Y(n_544) );
AO21x2_ASAP7_75t_L g580 ( .A1(n_180), .A2(n_545), .B(n_551), .Y(n_580) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_180), .A2(n_512), .B(n_518), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_186), .Y(n_181) );
AND2x2_ASAP7_75t_L g216 ( .A(n_188), .B(n_217), .Y(n_216) );
INVx2_ASAP7_75t_SL g274 ( .A(n_188), .Y(n_274) );
NAND2x1_ASAP7_75t_L g284 ( .A(n_188), .B(n_200), .Y(n_284) );
OR2x2_ASAP7_75t_L g289 ( .A(n_188), .B(n_217), .Y(n_289) );
BUFx2_ASAP7_75t_L g345 ( .A(n_188), .Y(n_345) );
AND2x2_ASAP7_75t_L g381 ( .A(n_188), .B(n_260), .Y(n_381) );
AND2x2_ASAP7_75t_L g392 ( .A(n_188), .B(n_220), .Y(n_392) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_196), .Y(n_188) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_208), .B1(n_214), .B2(n_215), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_199), .A2(n_389), .B1(n_439), .B2(n_444), .Y(n_438) );
INVx4_ASAP7_75t_L g217 ( .A(n_200), .Y(n_217) );
INVx2_ASAP7_75t_L g258 ( .A(n_200), .Y(n_258) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_200), .Y(n_329) );
OR2x2_ASAP7_75t_L g344 ( .A(n_200), .B(n_220), .Y(n_344) );
OR2x2_ASAP7_75t_SL g370 ( .A(n_200), .B(n_371), .Y(n_370) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_209), .B(n_211), .Y(n_208) );
INVx2_ASAP7_75t_SL g251 ( .A(n_209), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_209), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g319 ( .A(n_209), .B(n_267), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_209), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g241 ( .A(n_210), .Y(n_241) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
AND2x2_ASAP7_75t_L g322 ( .A(n_210), .B(n_299), .Y(n_322) );
INVx1_ASAP7_75t_L g432 ( .A(n_210), .Y(n_432) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_212), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_212), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g240 ( .A(n_213), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_214), .B(n_373), .Y(n_372) );
AOI321xp33_ASAP7_75t_L g394 ( .A1(n_215), .A2(n_296), .A3(n_364), .B1(n_395), .B2(n_396), .C(n_400), .Y(n_394) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_218), .Y(n_215) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_216), .Y(n_293) );
AND2x2_ASAP7_75t_L g318 ( .A(n_216), .B(n_247), .Y(n_318) );
AND2x2_ASAP7_75t_L g393 ( .A(n_216), .B(n_303), .Y(n_393) );
INVx1_ASAP7_75t_L g262 ( .A(n_217), .Y(n_262) );
BUFx2_ASAP7_75t_L g272 ( .A(n_217), .Y(n_272) );
NOR2xp67_ASAP7_75t_L g379 ( .A(n_217), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g317 ( .A(n_218), .Y(n_317) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
BUFx2_ASAP7_75t_L g324 ( .A(n_219), .Y(n_324) );
INVx2_ASAP7_75t_L g260 ( .A(n_220), .Y(n_260) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_220), .Y(n_283) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AOI21xp33_ASAP7_75t_SL g222 ( .A1(n_223), .A2(n_242), .B(n_245), .Y(n_222) );
NOR2xp67_ASAP7_75t_L g376 ( .A(n_223), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_240), .Y(n_224) );
INVx3_ASAP7_75t_L g267 ( .A(n_225), .Y(n_267) );
AND2x2_ASAP7_75t_L g298 ( .A(n_225), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
AND2x4_ASAP7_75t_L g255 ( .A(n_226), .B(n_227), .Y(n_255) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_233), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
NOR2x1p5_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g338 ( .A(n_240), .Y(n_338) );
INVx1_ASAP7_75t_SL g423 ( .A(n_241), .Y(n_423) );
INVxp33_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_244), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g349 ( .A(n_244), .B(n_306), .Y(n_349) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
AND2x2_ASAP7_75t_L g353 ( .A(n_246), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_246), .B(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_247), .B(n_284), .Y(n_339) );
NOR4xp25_ASAP7_75t_L g434 ( .A(n_247), .B(n_278), .C(n_435), .D(n_436), .Y(n_434) );
OR2x2_ASAP7_75t_L g402 ( .A(n_248), .B(n_403), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_256), .B1(n_261), .B2(n_263), .C(n_268), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_L g277 ( .A(n_252), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g314 ( .A(n_253), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g334 ( .A(n_254), .Y(n_334) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx3_ASAP7_75t_L g357 ( .A(n_255), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_255), .B(n_365), .Y(n_364) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OR2x2_ASAP7_75t_L g301 ( .A(n_258), .B(n_302), .Y(n_301) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_260), .B(n_274), .Y(n_273) );
INVxp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx2_ASAP7_75t_L g278 ( .A(n_265), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_265), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g270 ( .A(n_267), .Y(n_270) );
OAI321xp33_ASAP7_75t_L g382 ( .A1(n_267), .A2(n_375), .A3(n_383), .B1(n_388), .B2(n_390), .C(n_394), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
OR2x2_ASAP7_75t_L g337 ( .A(n_270), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g437 ( .A(n_273), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_274), .B(n_317), .Y(n_316) );
NAND2xp33_ASAP7_75t_SL g417 ( .A(n_274), .B(n_288), .Y(n_417) );
OAI211xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .B(n_290), .C(n_294), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2x1_ASAP7_75t_L g279 ( .A(n_280), .B(n_285), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g386 ( .A(n_283), .Y(n_386) );
INVx3_ASAP7_75t_L g325 ( .A(n_284), .Y(n_325) );
OR2x2_ASAP7_75t_L g428 ( .A(n_284), .B(n_302), .Y(n_428) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_286), .A2(n_370), .B1(n_372), .B2(n_374), .Y(n_369) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_SL g368 ( .A(n_289), .Y(n_368) );
OR2x2_ASAP7_75t_L g445 ( .A(n_289), .B(n_302), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI21xp5_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_296), .B(n_300), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_298), .B(n_315), .Y(n_414) );
AND2x2_ASAP7_75t_L g420 ( .A(n_298), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g365 ( .A(n_299), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B1(n_307), .B2(n_309), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g346 ( .A1(n_302), .A2(n_345), .B(n_347), .C(n_349), .Y(n_346) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_305), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_305), .B(n_397), .Y(n_419) );
INVx2_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g391 ( .A(n_308), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_310), .A2(n_342), .B(n_345), .C(n_346), .Y(n_341) );
NAND3xp33_ASAP7_75t_SL g311 ( .A(n_312), .B(n_326), .C(n_341), .Y(n_311) );
AOI222xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B1(n_318), .B2(n_319), .C1(n_320), .C2(n_323), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g375 ( .A(n_315), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_315), .B(n_348), .Y(n_401) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g335 ( .A(n_322), .Y(n_335) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
OR2x2_ASAP7_75t_L g440 ( .A(n_324), .B(n_357), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_325), .A2(n_416), .B1(n_418), .B2(n_420), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_332), .B1(n_336), .B2(n_339), .C(n_340), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI21xp5_ASAP7_75t_SL g400 ( .A1(n_333), .A2(n_401), .B(n_402), .Y(n_400) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx2_ASAP7_75t_L g348 ( .A(n_334), .Y(n_348) );
AND2x2_ASAP7_75t_L g442 ( .A(n_334), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g426 ( .A(n_338), .Y(n_426) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g355 ( .A(n_344), .B(n_345), .Y(n_355) );
INVx1_ASAP7_75t_L g408 ( .A(n_344), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_382), .C(n_404), .Y(n_350) );
OAI211xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_356), .B(n_358), .C(n_363), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_353), .A2(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI211xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B(n_369), .C(n_376), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g387 ( .A(n_370), .Y(n_387) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_371), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_373), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g435 ( .A(n_373), .Y(n_435) );
AND2x2_ASAP7_75t_L g425 ( .A(n_375), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g395 ( .A(n_377), .Y(n_395) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_391), .A2(n_425), .B1(n_427), .B2(n_429), .C(n_434), .Y(n_424) );
OAI21xp33_ASAP7_75t_SL g439 ( .A1(n_396), .A2(n_440), .B(n_441), .Y(n_439) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_415), .C(n_424), .D(n_438), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B1(n_412), .B2(n_413), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_433), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
CKINVDCx6p67_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
AND2x6_ASAP7_75t_SL g449 ( .A(n_450), .B(n_451), .Y(n_449) );
OR2x6_ASAP7_75t_SL g745 ( .A(n_450), .B(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g755 ( .A(n_450), .B(n_451), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_450), .B(n_746), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_451), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx2_ASAP7_75t_L g749 ( .A(n_455), .Y(n_749) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_643), .Y(n_455) );
NAND3xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_555), .C(n_610), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_496), .B1(n_519), .B2(n_523), .C(n_533), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_480), .Y(n_458) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_459), .B(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g554 ( .A(n_459), .Y(n_554) );
AND2x2_ASAP7_75t_L g599 ( .A(n_459), .B(n_536), .Y(n_599) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g587 ( .A(n_461), .Y(n_587) );
INVx1_ASAP7_75t_L g597 ( .A(n_461), .Y(n_597) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_469), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_462), .B(n_470), .Y(n_469) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_462), .A2(n_463), .B(n_469), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_468), .Y(n_463) );
OR2x2_ASAP7_75t_L g576 ( .A(n_471), .B(n_481), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_471), .B(n_522), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_471), .B(n_488), .Y(n_620) );
INVx2_ASAP7_75t_L g629 ( .A(n_471), .Y(n_629) );
AND2x2_ASAP7_75t_L g650 ( .A(n_471), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g734 ( .A(n_471), .B(n_553), .Y(n_734) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g562 ( .A(n_472), .B(n_488), .Y(n_562) );
AND2x2_ASAP7_75t_L g695 ( .A(n_472), .B(n_522), .Y(n_695) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_472), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
AND2x4_ASAP7_75t_L g649 ( .A(n_480), .B(n_650), .Y(n_649) );
AOI321xp33_ASAP7_75t_L g663 ( .A1(n_480), .A2(n_592), .A3(n_593), .B1(n_625), .B2(n_664), .C(n_667), .Y(n_663) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_488), .Y(n_480) );
BUFx3_ASAP7_75t_L g520 ( .A(n_481), .Y(n_520) );
INVx2_ASAP7_75t_L g553 ( .A(n_481), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_481), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g586 ( .A(n_481), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g619 ( .A(n_481), .Y(n_619) );
INVx5_ASAP7_75t_L g522 ( .A(n_488), .Y(n_522) );
NOR2x1_ASAP7_75t_SL g571 ( .A(n_488), .B(n_561), .Y(n_571) );
BUFx2_ASAP7_75t_L g666 ( .A(n_488), .Y(n_666) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVxp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_509), .Y(n_497) );
NOR2xp33_ASAP7_75t_SL g564 ( .A(n_498), .B(n_565), .Y(n_564) );
NOR4xp25_ASAP7_75t_L g667 ( .A(n_498), .B(n_661), .C(n_665), .D(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g705 ( .A(n_498), .Y(n_705) );
AND2x2_ASAP7_75t_L g739 ( .A(n_498), .B(n_679), .Y(n_739) );
BUFx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g540 ( .A(n_499), .Y(n_540) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g594 ( .A(n_500), .Y(n_594) );
OAI21x1_ASAP7_75t_SL g500 ( .A1(n_501), .A2(n_503), .B(n_507), .Y(n_500) );
INVx1_ASAP7_75t_L g508 ( .A(n_502), .Y(n_508) );
AOI33xp33_ASAP7_75t_L g735 ( .A1(n_509), .A2(n_537), .A3(n_568), .B1(n_584), .B2(n_690), .B3(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g525 ( .A(n_510), .B(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g535 ( .A(n_510), .B(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g542 ( .A(n_511), .Y(n_542) );
INVxp67_ASAP7_75t_L g623 ( .A(n_511), .Y(n_623) );
AND2x2_ASAP7_75t_L g679 ( .A(n_511), .B(n_544), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_519), .A2(n_701), .B(n_702), .Y(n_700) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AND2x2_ASAP7_75t_L g688 ( .A(n_520), .B(n_562), .Y(n_688) );
AND3x2_ASAP7_75t_L g690 ( .A(n_520), .B(n_574), .C(n_629), .Y(n_690) );
INVx3_ASAP7_75t_SL g642 ( .A(n_521), .Y(n_642) );
INVx4_ASAP7_75t_L g536 ( .A(n_522), .Y(n_536) );
AND2x2_ASAP7_75t_L g574 ( .A(n_522), .B(n_561), .Y(n_574) );
INVxp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g568 ( .A(n_526), .Y(n_568) );
AND2x4_ASAP7_75t_L g593 ( .A(n_526), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g656 ( .A(n_526), .B(n_544), .Y(n_656) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g626 ( .A(n_527), .Y(n_626) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_527), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_R g533 ( .A1(n_534), .A2(n_537), .B(n_541), .C(n_552), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g585 ( .A(n_536), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_536), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_536), .B(n_553), .Y(n_714) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g696 ( .A(n_538), .B(n_686), .Y(n_696) );
AND2x2_ASAP7_75t_SL g538 ( .A(n_539), .B(n_540), .Y(n_538) );
AND2x2_ASAP7_75t_L g543 ( .A(n_539), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g565 ( .A(n_539), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g581 ( .A(n_539), .B(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_L g614 ( .A(n_539), .B(n_594), .Y(n_614) );
AND2x4_ASAP7_75t_L g579 ( .A(n_540), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g603 ( .A(n_540), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g641 ( .A(n_540), .B(n_566), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
AND2x2_ASAP7_75t_L g569 ( .A(n_542), .B(n_566), .Y(n_569) );
AND2x2_ASAP7_75t_L g584 ( .A(n_542), .B(n_544), .Y(n_584) );
BUFx2_ASAP7_75t_L g640 ( .A(n_542), .Y(n_640) );
AND2x2_ASAP7_75t_L g654 ( .A(n_542), .B(n_565), .Y(n_654) );
INVx2_ASAP7_75t_L g566 ( .A(n_544), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_550), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_552), .A2(n_603), .B1(n_605), .B2(n_609), .Y(n_602) );
INVx2_ASAP7_75t_SL g633 ( .A(n_552), .Y(n_633) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x2_ASAP7_75t_L g608 ( .A(n_553), .B(n_561), .Y(n_608) );
INVx1_ASAP7_75t_L g715 ( .A(n_554), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_588), .C(n_602), .Y(n_555) );
OAI221xp5_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_563), .B1(n_567), .B2(n_570), .C(n_572), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g616 ( .A(n_560), .Y(n_616) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_560), .Y(n_744) );
INVx1_ASAP7_75t_L g707 ( .A(n_562), .Y(n_707) );
AND2x2_ASAP7_75t_SL g717 ( .A(n_562), .B(n_586), .Y(n_717) );
INVxp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_566), .B(n_594), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OR2x2_ASAP7_75t_L g600 ( .A(n_568), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g678 ( .A(n_568), .Y(n_678) );
AND2x2_ASAP7_75t_L g613 ( .A(n_569), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g659 ( .A(n_571), .B(n_619), .Y(n_659) );
AND2x2_ASAP7_75t_L g736 ( .A(n_571), .B(n_734), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .B1(n_584), .B2(n_585), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g595 ( .A(n_576), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx2_ASAP7_75t_L g601 ( .A(n_579), .Y(n_601) );
AND2x4_ASAP7_75t_L g625 ( .A(n_579), .B(n_626), .Y(n_625) );
OAI21xp33_ASAP7_75t_SL g655 ( .A1(n_579), .A2(n_656), .B(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g682 ( .A(n_579), .B(n_640), .Y(n_682) );
INVx2_ASAP7_75t_L g604 ( .A(n_580), .Y(n_604) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_580), .Y(n_637) );
INVx1_ASAP7_75t_SL g661 ( .A(n_581), .Y(n_661) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g592 ( .A(n_583), .Y(n_592) );
AND2x4_ASAP7_75t_SL g686 ( .A(n_583), .B(n_604), .Y(n_686) );
AND2x2_ASAP7_75t_L g683 ( .A(n_586), .B(n_629), .Y(n_683) );
AND2x2_ASAP7_75t_L g709 ( .A(n_586), .B(n_695), .Y(n_709) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_587), .Y(n_631) );
INVx1_ASAP7_75t_L g651 ( .A(n_587), .Y(n_651) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_595), .B1(n_598), .B2(n_600), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_593), .B(n_604), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_593), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g732 ( .A(n_593), .Y(n_732) );
INVx2_ASAP7_75t_SL g657 ( .A(n_595), .Y(n_657) );
AND2x2_ASAP7_75t_L g669 ( .A(n_597), .B(n_629), .Y(n_669) );
INVx2_ASAP7_75t_L g675 ( .A(n_597), .Y(n_675) );
INVxp33_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g634 ( .A(n_600), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_603), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g725 ( .A(n_603), .Y(n_725) );
INVx1_ASAP7_75t_L g653 ( .A(n_605), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_606), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g664 ( .A(n_608), .B(n_665), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_608), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_632), .C(n_635), .Y(n_610) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B1(n_617), .B2(n_621), .C(n_624), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g730 ( .A(n_615), .Y(n_730) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g699 ( .A(n_616), .B(n_665), .Y(n_699) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g630 ( .A(n_619), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g701 ( .A(n_621), .Y(n_701) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g698 ( .A(n_622), .Y(n_698) );
INVx1_ASAP7_75t_L g704 ( .A(n_623), .Y(n_704) );
OR2x2_ASAP7_75t_L g727 ( .A(n_623), .B(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_SL g636 ( .A(n_626), .Y(n_636) );
AND2x2_ASAP7_75t_L g706 ( .A(n_626), .B(n_686), .Y(n_706) );
AND2x2_ASAP7_75t_SL g738 ( .A(n_626), .B(n_639), .Y(n_738) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g743 ( .A(n_629), .Y(n_743) );
INVx1_ASAP7_75t_L g693 ( .A(n_631), .Y(n_693) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_638), .C(n_642), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_636), .B(n_686), .Y(n_710) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_639), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g647 ( .A(n_641), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g728 ( .A(n_641), .Y(n_728) );
NAND4xp75_ASAP7_75t_L g643 ( .A(n_644), .B(n_700), .C(n_716), .D(n_737), .Y(n_643) );
NOR3x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_662), .C(n_684), .Y(n_644) );
NAND4xp75_ASAP7_75t_L g645 ( .A(n_646), .B(n_652), .C(n_655), .D(n_658), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_647), .B(n_649), .Y(n_646) );
AND2x2_ASAP7_75t_L g697 ( .A(n_648), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g722 ( .A(n_649), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_SL g711 ( .A(n_654), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_670), .Y(n_662) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_666), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_676), .B(n_680), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI322xp33_ASAP7_75t_L g702 ( .A1(n_674), .A2(n_703), .A3(n_707), .B1(n_708), .B2(n_710), .C1(n_711), .C2(n_712), .Y(n_702) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_675), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_678), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_679), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_689), .C(n_691), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_696), .B1(n_697), .B2(n_699), .Y(n_691) );
NOR2xp33_ASAP7_75t_SL g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B(n_706), .Y(n_703) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_709), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_713), .B(n_715), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g719 ( .A(n_714), .B(n_720), .Y(n_719) );
O2A1O1Ixp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B(n_723), .C(n_726), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_719), .B(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI221xp5_ASAP7_75t_SL g726 ( .A1(n_727), .A2(n_729), .B1(n_731), .B2(n_733), .C(n_735), .Y(n_726) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
CKINVDCx11_ASAP7_75t_R g751 ( .A(n_745), .Y(n_751) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
INVx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_765), .Y(n_758) );
INVxp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_761), .B(n_764), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_SL g788 ( .A(n_762), .B(n_764), .Y(n_788) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_762), .A2(n_791), .B(n_794), .Y(n_790) );
BUFx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
BUFx2_ASAP7_75t_R g771 ( .A(n_766), .Y(n_771) );
BUFx3_ASAP7_75t_L g783 ( .A(n_766), .Y(n_783) );
BUFx2_ASAP7_75t_L g795 ( .A(n_766), .Y(n_795) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AOI21xp33_ASAP7_75t_SL g768 ( .A1(n_769), .A2(n_772), .B(n_781), .Y(n_768) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
NOR2xp33_ASAP7_75t_SL g781 ( .A(n_782), .B(n_784), .Y(n_781) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
CKINVDCx9p33_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
CKINVDCx8_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
endmodule