module fake_jpeg_29568_n_140 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_8),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_48),
.B1(n_52),
.B2(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_15),
.B1(n_28),
.B2(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_15),
.B1(n_28),
.B2(n_17),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_25),
.B(n_17),
.C(n_15),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_25),
.B1(n_24),
.B2(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_41),
.B1(n_35),
.B2(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_65),
.Y(n_90)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_78),
.B1(n_51),
.B2(n_49),
.Y(n_85)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_36),
.B1(n_35),
.B2(n_37),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_53),
.B1(n_62),
.B2(n_3),
.Y(n_89)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_77),
.B1(n_62),
.B2(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_76),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_38),
.B1(n_24),
.B2(n_18),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_2),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_5),
.B(n_6),
.C(n_10),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_18),
.Y(n_81)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_53),
.A3(n_51),
.B1(n_49),
.B2(n_62),
.Y(n_83)
);

OAI31xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_68),
.A3(n_64),
.B(n_76),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_89),
.B1(n_66),
.B2(n_80),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_69),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_91),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_6),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_71),
.B(n_73),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_89),
.B(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_105),
.B1(n_92),
.B2(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_65),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_67),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_93),
.C(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_70),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_114),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_115),
.B1(n_97),
.B2(n_82),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_92),
.C(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_113),
.Y(n_118)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_101),
.C(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_113),
.C(n_109),
.Y(n_124)
);

AOI222xp33_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_97),
.B1(n_105),
.B2(n_99),
.C1(n_96),
.C2(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_123),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_128),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_123),
.B(n_121),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_11),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_120),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_127),
.B(n_116),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_131),
.B(n_12),
.Y(n_136)
);

AOI21x1_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_128),
.B(n_131),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_136),
.B(n_11),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_13),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_13),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);


endmodule