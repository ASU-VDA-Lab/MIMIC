module real_jpeg_3660_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_32),
.B1(n_34),
.B2(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_32),
.B1(n_38),
.B2(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_38),
.B1(n_46),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_34),
.B1(n_51),
.B2(n_60),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_51),
.Y(n_123)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_7),
.B(n_37),
.C(n_38),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_34),
.B1(n_60),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_7),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_7),
.B(n_57),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_7),
.B(n_24),
.C(n_47),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_7),
.A2(n_38),
.B1(n_46),
.B2(n_62),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_7),
.B(n_21),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_7),
.B(n_71),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_8),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_38),
.B1(n_46),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_53),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_10),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_92),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_91),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_65),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_17),
.B(n_65),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_42),
.C(n_54),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_18),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_18)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_19),
.B(n_41),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B(n_28),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_24),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_20),
.A2(n_22),
.B1(n_30),
.B2(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_20),
.B(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_20),
.A2(n_30),
.B1(n_97),
.B2(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_21),
.A2(n_29),
.B(n_123),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_30),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_37),
.B1(n_58),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_34),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_34),
.A2(n_60),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_38),
.B1(n_46),
.B2(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_38),
.B(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_42),
.B(n_54),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_43),
.A2(n_70),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_68),
.B(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_44),
.B(n_72),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_49),
.A2(n_50),
.B(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_63),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_62),
.A2(n_99),
.B(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_74),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_73),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_87),
.B2(n_88),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_133),
.B(n_137),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_114),
.B(n_132),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_108),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_108),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_106),
.B2(n_107),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_103),
.C(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_126),
.B(n_131),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_121),
.B(n_125),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_124),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_129),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);


endmodule