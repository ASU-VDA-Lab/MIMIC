module fake_jpeg_3446_n_54 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_54);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_25),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_20),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_21),
.B(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_18),
.B1(n_20),
.B2(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_32),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_27),
.B(n_18),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.C(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_23),
.B(n_2),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_0),
.C(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_36),
.B1(n_31),
.B2(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_4),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_14),
.C(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_5),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_46),
.B1(n_6),
.B2(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_49),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_50),
.B(n_6),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_5),
.C(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_8),
.Y(n_54)
);


endmodule