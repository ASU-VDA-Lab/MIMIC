module real_aes_1881_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_0), .B(n_147), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_1), .A2(n_141), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_2), .B(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_3), .B(n_158), .Y(n_233) );
INVx1_ASAP7_75t_L g146 ( .A(n_4), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_5), .B(n_158), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_6), .B(n_210), .Y(n_498) );
INVx1_ASAP7_75t_L g541 ( .A(n_7), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g810 ( .A(n_8), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_9), .Y(n_555) );
NAND2xp33_ASAP7_75t_L g209 ( .A(n_10), .B(n_156), .Y(n_209) );
INVx2_ASAP7_75t_L g138 ( .A(n_11), .Y(n_138) );
AOI221x1_ASAP7_75t_L g140 ( .A1(n_12), .A2(n_24), .B1(n_141), .B2(n_147), .C(n_154), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_13), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g808 ( .A(n_13), .B(n_809), .C(n_811), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_14), .B(n_147), .Y(n_205) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_15), .A2(n_203), .B(n_204), .Y(n_202) );
INVx1_ASAP7_75t_L g507 ( .A(n_16), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_17), .B(n_136), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_18), .B(n_158), .Y(n_217) );
AO21x1_ASAP7_75t_L g228 ( .A1(n_19), .A2(n_147), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g117 ( .A(n_20), .Y(n_117) );
NOR2xp33_ASAP7_75t_SL g806 ( .A(n_20), .B(n_118), .Y(n_806) );
INVx1_ASAP7_75t_L g505 ( .A(n_21), .Y(n_505) );
INVx1_ASAP7_75t_SL g491 ( .A(n_22), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_23), .B(n_148), .Y(n_469) );
NAND2x1_ASAP7_75t_L g166 ( .A(n_25), .B(n_158), .Y(n_166) );
AOI33xp33_ASAP7_75t_L g522 ( .A1(n_26), .A2(n_55), .A3(n_457), .B1(n_466), .B2(n_523), .B3(n_524), .Y(n_522) );
NAND2x1_ASAP7_75t_L g196 ( .A(n_27), .B(n_156), .Y(n_196) );
INVx1_ASAP7_75t_L g549 ( .A(n_28), .Y(n_549) );
OR2x2_ASAP7_75t_L g139 ( .A(n_29), .B(n_91), .Y(n_139) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_29), .A2(n_91), .B(n_138), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_30), .B(n_482), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_31), .B(n_156), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_32), .A2(n_33), .B1(n_785), .B2(n_786), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_32), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_33), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_34), .B(n_158), .Y(n_208) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_35), .A2(n_36), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_35), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_36), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_37), .B(n_156), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_38), .A2(n_141), .B(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g142 ( .A(n_39), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g153 ( .A(n_39), .B(n_146), .Y(n_153) );
INVx1_ASAP7_75t_L g465 ( .A(n_39), .Y(n_465) );
OR2x6_ASAP7_75t_L g115 ( .A(n_40), .B(n_116), .Y(n_115) );
INVxp67_ASAP7_75t_L g811 ( .A(n_40), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_41), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_42), .B(n_147), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_43), .B(n_482), .Y(n_529) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_44), .A2(n_89), .B1(n_121), .B2(n_122), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_44), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_44), .A2(n_171), .B1(n_210), .B2(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_45), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_46), .B(n_148), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_47), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_48), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_49), .B(n_156), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_50), .B(n_203), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_51), .B(n_148), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_52), .A2(n_141), .B(n_195), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_53), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_54), .B(n_156), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_56), .B(n_148), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_57), .Y(n_813) );
INVx1_ASAP7_75t_L g145 ( .A(n_58), .Y(n_145) );
INVx1_ASAP7_75t_L g150 ( .A(n_58), .Y(n_150) );
AND2x2_ASAP7_75t_L g534 ( .A(n_59), .B(n_136), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_60), .A2(n_78), .B1(n_463), .B2(n_482), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_61), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_62), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_63), .B(n_171), .Y(n_557) );
AOI21xp5_ASAP7_75t_SL g477 ( .A1(n_64), .A2(n_463), .B(n_478), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_65), .A2(n_141), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g501 ( .A(n_66), .Y(n_501) );
AO21x1_ASAP7_75t_L g230 ( .A1(n_67), .A2(n_141), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_68), .B(n_147), .Y(n_187) );
INVx1_ASAP7_75t_L g532 ( .A(n_69), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_70), .B(n_147), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_71), .A2(n_463), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g181 ( .A(n_72), .B(n_137), .Y(n_181) );
INVx1_ASAP7_75t_L g143 ( .A(n_73), .Y(n_143) );
INVx1_ASAP7_75t_L g152 ( .A(n_73), .Y(n_152) );
AND2x2_ASAP7_75t_L g200 ( .A(n_74), .B(n_170), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_75), .B(n_482), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_76), .B(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_77), .A2(n_780), .B1(n_781), .B2(n_782), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_77), .Y(n_780) );
AND2x2_ASAP7_75t_L g493 ( .A(n_79), .B(n_170), .Y(n_493) );
INVx1_ASAP7_75t_L g502 ( .A(n_80), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_81), .A2(n_463), .B(n_490), .Y(n_489) );
OAI22xp5_ASAP7_75t_SL g782 ( .A1(n_82), .A2(n_783), .B1(n_784), .B2(n_787), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_82), .Y(n_787) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_83), .A2(n_463), .B(n_468), .C(n_473), .Y(n_462) );
INVx1_ASAP7_75t_L g118 ( .A(n_84), .Y(n_118) );
AND2x2_ASAP7_75t_L g185 ( .A(n_85), .B(n_170), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_86), .B(n_147), .Y(n_219) );
AND2x2_ASAP7_75t_SL g475 ( .A(n_87), .B(n_170), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_88), .A2(n_463), .B1(n_520), .B2(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
AND2x2_ASAP7_75t_L g229 ( .A(n_90), .B(n_210), .Y(n_229) );
AND2x2_ASAP7_75t_L g173 ( .A(n_92), .B(n_170), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_93), .B(n_156), .Y(n_218) );
INVx1_ASAP7_75t_L g479 ( .A(n_94), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_95), .B(n_158), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_96), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_97), .A2(n_141), .B(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g526 ( .A(n_98), .B(n_170), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_99), .B(n_158), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_100), .A2(n_547), .B(n_548), .C(n_550), .Y(n_546) );
BUFx2_ASAP7_75t_L g108 ( .A(n_101), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_102), .A2(n_141), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_103), .B(n_148), .Y(n_480) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_801), .B(n_812), .Y(n_104) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_109), .B(n_440), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_108), .Y(n_800) );
OAI21x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_119), .B(n_435), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g439 ( .A(n_112), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OR2x6_ASAP7_75t_SL g775 ( .A(n_113), .B(n_114), .Y(n_775) );
AND2x6_ASAP7_75t_SL g778 ( .A(n_113), .B(n_115), .Y(n_778) );
OR2x2_ASAP7_75t_L g799 ( .A(n_113), .B(n_115), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B1(n_433), .B2(n_434), .Y(n_119) );
INVx1_ASAP7_75t_L g433 ( .A(n_120), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_123), .Y(n_434) );
XOR2x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
INVx3_ASAP7_75t_L g776 ( .A(n_127), .Y(n_776) );
OAI22xp5_ASAP7_75t_SL g790 ( .A1(n_127), .A2(n_791), .B1(n_793), .B2(n_794), .Y(n_790) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_345), .Y(n_127) );
AND4x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_257), .C(n_284), .D(n_319), .Y(n_128) );
AOI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_182), .B1(n_222), .B2(n_237), .C(n_241), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_161), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_132), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g298 ( .A(n_133), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g353 ( .A(n_133), .B(n_308), .Y(n_353) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g256 ( .A(n_134), .B(n_174), .Y(n_256) );
AND2x4_ASAP7_75t_L g292 ( .A(n_134), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g306 ( .A(n_134), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g223 ( .A(n_135), .Y(n_223) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_135), .Y(n_395) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B(n_160), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_136), .A2(n_187), .B(n_188), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_136), .Y(n_199) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_136), .A2(n_140), .B(n_160), .Y(n_269) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x4_ASAP7_75t_L g210 ( .A(n_138), .B(n_139), .Y(n_210) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
BUFx3_ASAP7_75t_L g460 ( .A(n_142), .Y(n_460) );
AND2x6_ASAP7_75t_L g156 ( .A(n_143), .B(n_149), .Y(n_156) );
INVx2_ASAP7_75t_L g467 ( .A(n_143), .Y(n_467) );
AND2x4_ASAP7_75t_L g463 ( .A(n_144), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g158 ( .A(n_145), .B(n_151), .Y(n_158) );
INVx2_ASAP7_75t_L g457 ( .A(n_145), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_146), .Y(n_458) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_153), .Y(n_147) );
INVx1_ASAP7_75t_L g503 ( .A(n_148), .Y(n_503) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx5_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_153), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
INVxp67_ASAP7_75t_L g506 ( .A(n_156), .Y(n_506) );
INVxp67_ASAP7_75t_L g508 ( .A(n_158), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_159), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_159), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_159), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_159), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_159), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_159), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_159), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_159), .A2(n_469), .B(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_159), .A2(n_472), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_159), .A2(n_472), .B(n_491), .C(n_492), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_159), .B(n_210), .Y(n_509) );
INVx1_ASAP7_75t_L g520 ( .A(n_159), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_159), .A2(n_472), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g540 ( .A1(n_159), .A2(n_472), .B(n_541), .C(n_542), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_SL g250 ( .A1(n_161), .A2(n_223), .B(n_251), .C(n_255), .Y(n_250) );
AND2x2_ASAP7_75t_L g271 ( .A(n_161), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_161), .B(n_223), .Y(n_411) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_174), .Y(n_161) );
INVx2_ASAP7_75t_L g291 ( .A(n_162), .Y(n_291) );
BUFx3_ASAP7_75t_L g307 ( .A(n_162), .Y(n_307) );
INVxp67_ASAP7_75t_L g311 ( .A(n_162), .Y(n_311) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_169), .B(n_173), .Y(n_162) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_163), .A2(n_169), .B(n_173), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_168), .Y(n_163) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_169), .A2(n_175), .B(n_181), .Y(n_174) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_169), .A2(n_175), .B(n_181), .Y(n_236) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_169), .A2(n_528), .B(n_534), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_169), .A2(n_170), .B1(n_546), .B2(n_551), .Y(n_545) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_169), .A2(n_528), .B(n_534), .Y(n_564) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_171), .B(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx4f_ASAP7_75t_L g203 ( .A(n_172), .Y(n_203) );
INVx2_ASAP7_75t_L g290 ( .A(n_174), .Y(n_290) );
AND2x2_ASAP7_75t_L g296 ( .A(n_174), .B(n_269), .Y(n_296) );
AND2x2_ASAP7_75t_L g322 ( .A(n_174), .B(n_291), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_176), .B(n_180), .Y(n_175) );
AOI211xp5_ASAP7_75t_L g319 ( .A1(n_182), .A2(n_320), .B(n_323), .C(n_333), .Y(n_319) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_183), .B(n_201), .Y(n_182) );
OAI321xp33_ASAP7_75t_L g294 ( .A1(n_183), .A2(n_242), .A3(n_295), .B1(n_297), .B2(n_298), .C(n_300), .Y(n_294) );
AND2x2_ASAP7_75t_L g415 ( .A(n_183), .B(n_390), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_183), .Y(n_418) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_192), .Y(n_183) );
INVx5_ASAP7_75t_L g240 ( .A(n_184), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_184), .B(n_254), .Y(n_253) );
NOR2x1_ASAP7_75t_SL g285 ( .A(n_184), .B(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g330 ( .A(n_184), .Y(n_330) );
AND2x2_ASAP7_75t_L g432 ( .A(n_184), .B(n_202), .Y(n_432) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
AND2x2_ASAP7_75t_L g239 ( .A(n_192), .B(n_240), .Y(n_239) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_192), .Y(n_249) );
INVx4_ASAP7_75t_L g254 ( .A(n_192), .Y(n_254) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_199), .B(n_200), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_198), .Y(n_193) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_199), .A2(n_487), .B(n_493), .Y(n_486) );
INVx1_ASAP7_75t_L g297 ( .A(n_201), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_R g400 ( .A1(n_201), .A2(n_239), .B(n_271), .C(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g420 ( .A(n_201), .B(n_245), .Y(n_420) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_211), .Y(n_201) );
INVx1_ASAP7_75t_L g238 ( .A(n_202), .Y(n_238) );
INVx2_ASAP7_75t_L g244 ( .A(n_202), .Y(n_244) );
OR2x2_ASAP7_75t_L g263 ( .A(n_202), .B(n_254), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_202), .B(n_286), .Y(n_332) );
BUFx3_ASAP7_75t_L g339 ( .A(n_202), .Y(n_339) );
INVx2_ASAP7_75t_SL g473 ( .A(n_203), .Y(n_473) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_203), .A2(n_539), .B(n_543), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_210), .Y(n_204) );
INVx1_ASAP7_75t_SL g213 ( .A(n_210), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_210), .B(n_235), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_210), .A2(n_477), .B(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g302 ( .A(n_211), .Y(n_302) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_211), .Y(n_315) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g248 ( .A(n_212), .Y(n_248) );
INVx1_ASAP7_75t_L g357 ( .A(n_212), .Y(n_357) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_220), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_213), .B(n_221), .Y(n_220) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_213), .A2(n_214), .B(n_220), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_219), .Y(n_214) );
AND2x2_ASAP7_75t_L g258 ( .A(n_222), .B(n_259), .Y(n_258) );
OAI31xp33_ASAP7_75t_L g409 ( .A1(n_222), .A2(n_410), .A3(n_412), .B(n_415), .Y(n_409) );
INVx1_ASAP7_75t_SL g427 ( .A(n_222), .Y(n_427) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
AOI21xp33_ASAP7_75t_L g241 ( .A1(n_223), .A2(n_242), .B(n_250), .Y(n_241) );
NAND2x1_ASAP7_75t_L g321 ( .A(n_223), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g350 ( .A(n_223), .Y(n_350) );
INVx2_ASAP7_75t_L g299 ( .A(n_224), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_224), .B(n_282), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_224), .B(n_281), .Y(n_391) );
NOR2xp33_ASAP7_75t_SL g399 ( .A(n_224), .B(n_350), .Y(n_399) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_236), .Y(n_224) );
AND2x2_ASAP7_75t_SL g268 ( .A(n_225), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g279 ( .A(n_225), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g308 ( .A(n_225), .B(n_290), .Y(n_308) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
BUFx2_ASAP7_75t_L g272 ( .A(n_226), .Y(n_272) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g293 ( .A(n_227), .Y(n_293) );
OAI21x1_ASAP7_75t_SL g227 ( .A1(n_228), .A2(n_230), .B(n_234), .Y(n_227) );
INVx1_ASAP7_75t_L g235 ( .A(n_229), .Y(n_235) );
INVx2_ASAP7_75t_L g280 ( .A(n_236), .Y(n_280) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_236), .Y(n_340) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx1_ASAP7_75t_L g276 ( .A(n_238), .Y(n_276) );
AND2x2_ASAP7_75t_L g355 ( .A(n_238), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g266 ( .A(n_239), .B(n_260), .Y(n_266) );
INVx2_ASAP7_75t_SL g314 ( .A(n_239), .Y(n_314) );
INVx4_ASAP7_75t_L g245 ( .A(n_240), .Y(n_245) );
AND2x2_ASAP7_75t_L g343 ( .A(n_240), .B(n_286), .Y(n_343) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_240), .B(n_356), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g378 ( .A(n_240), .B(n_254), .Y(n_378) );
INVx1_ASAP7_75t_L g384 ( .A(n_242), .Y(n_384) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_246), .Y(n_242) );
INVx1_ASAP7_75t_L g303 ( .A(n_243), .Y(n_303) );
OR2x2_ASAP7_75t_L g316 ( .A(n_243), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
OR2x2_ASAP7_75t_L g368 ( .A(n_244), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g398 ( .A(n_244), .B(n_286), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_245), .B(n_248), .Y(n_274) );
AND2x2_ASAP7_75t_L g366 ( .A(n_245), .B(n_356), .Y(n_366) );
AND2x4_ASAP7_75t_L g428 ( .A(n_245), .B(n_307), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
INVx2_ASAP7_75t_L g252 ( .A(n_247), .Y(n_252) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NOR2xp67_ASAP7_75t_SL g251 ( .A(n_252), .B(n_253), .Y(n_251) );
OAI322xp33_ASAP7_75t_SL g264 ( .A1(n_252), .A2(n_265), .A3(n_267), .B1(n_270), .B2(n_273), .C1(n_275), .C2(n_277), .Y(n_264) );
INVx1_ASAP7_75t_L g422 ( .A(n_252), .Y(n_422) );
OR2x2_ASAP7_75t_L g275 ( .A(n_253), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g301 ( .A(n_254), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_254), .B(n_302), .Y(n_317) );
INVx2_ASAP7_75t_L g344 ( .A(n_254), .Y(n_344) );
AND2x4_ASAP7_75t_L g356 ( .A(n_254), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_SL g359 ( .A(n_256), .B(n_272), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_262), .B(n_264), .Y(n_257) );
AND2x2_ASAP7_75t_L g325 ( .A(n_259), .B(n_292), .Y(n_325) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_260), .B(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
AND2x4_ASAP7_75t_SL g365 ( .A(n_261), .B(n_280), .Y(n_365) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g273 ( .A(n_263), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_266), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g401 ( .A(n_268), .B(n_365), .Y(n_401) );
NOR4xp25_ASAP7_75t_L g405 ( .A(n_268), .B(n_282), .C(n_322), .D(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g282 ( .A(n_269), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g318 ( .A(n_269), .B(n_293), .Y(n_318) );
AND2x4_ASAP7_75t_L g382 ( .A(n_269), .B(n_293), .Y(n_382) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_272), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
OR2x2_ASAP7_75t_L g371 ( .A(n_279), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g425 ( .A(n_279), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_280), .B(n_292), .Y(n_326) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AOI211xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_287), .B(n_294), .C(n_309), .Y(n_284) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_290), .B(n_293), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_291), .B(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g373 ( .A(n_291), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_292), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g388 ( .A(n_292), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B(n_304), .Y(n_300) );
AND2x4_ASAP7_75t_L g337 ( .A(n_301), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g431 ( .A(n_301), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_SL g335 ( .A(n_307), .Y(n_335) );
AND2x2_ASAP7_75t_L g394 ( .A(n_308), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g408 ( .A(n_308), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_312), .B(n_316), .C(n_318), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_310), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g386 ( .A(n_311), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g407 ( .A(n_311), .B(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
OR2x2_ASAP7_75t_L g396 ( .A(n_314), .B(n_338), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_317), .A2(n_324), .B1(n_326), .B2(n_327), .Y(n_323) );
INVx1_ASAP7_75t_SL g414 ( .A(n_318), .Y(n_414) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVxp67_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_329), .B(n_338), .Y(n_380) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_332), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B1(n_340), .B2(n_341), .Y(n_333) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI21xp5_ASAP7_75t_SL g347 ( .A1(n_338), .A2(n_348), .B(n_351), .Y(n_347) );
AND2x2_ASAP7_75t_L g376 ( .A(n_338), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND3x2_ASAP7_75t_L g342 ( .A(n_339), .B(n_343), .C(n_344), .Y(n_342) );
AND2x2_ASAP7_75t_L g404 ( .A(n_339), .B(n_361), .Y(n_404) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g389 ( .A(n_344), .B(n_390), .Y(n_389) );
NOR2xp67_ASAP7_75t_L g345 ( .A(n_346), .B(n_402), .Y(n_345) );
NAND4xp25_ASAP7_75t_L g346 ( .A(n_347), .B(n_362), .C(n_383), .D(n_400), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B1(n_358), .B2(n_360), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_354), .A2(n_368), .B1(n_388), .B2(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g369 ( .A(n_356), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_358), .A2(n_381), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx3_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B1(n_367), .B2(n_370), .C(n_374), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_379), .B1(n_380), .B2(n_381), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_377), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_377), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_389), .B2(n_391), .C(n_392), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_386), .B(n_388), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B1(n_397), .B2(n_399), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI211xp5_ASAP7_75t_SL g417 ( .A1(n_398), .A2(n_418), .B(n_419), .C(n_421), .Y(n_417) );
OAI211xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B(n_409), .C(n_416), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_423), .B1(n_426), .B2(n_428), .C(n_429), .Y(n_416) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
AOI31xp33_ASAP7_75t_L g440 ( .A1(n_435), .A2(n_441), .A3(n_788), .B(n_800), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
CKINVDCx11_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_779), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g793 ( .A(n_445), .Y(n_793) );
NAND4xp75_ASAP7_75t_L g445 ( .A(n_446), .B(n_626), .C(n_692), .D(n_755), .Y(n_445) );
NOR2x1_ASAP7_75t_L g446 ( .A(n_447), .B(n_589), .Y(n_446) );
OR3x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_559), .C(n_586), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_494), .B(n_515), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_483), .Y(n_450) );
AND2x2_ASAP7_75t_L g689 ( .A(n_451), .B(n_659), .Y(n_689) );
INVx1_ASAP7_75t_L g762 ( .A(n_451), .Y(n_762) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_474), .Y(n_451) );
INVx2_ASAP7_75t_L g514 ( .A(n_452), .Y(n_514) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_452), .Y(n_577) );
AND2x2_ASAP7_75t_L g581 ( .A(n_452), .B(n_497), .Y(n_581) );
AND2x4_ASAP7_75t_L g597 ( .A(n_452), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g601 ( .A(n_452), .Y(n_601) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_459), .C(n_461), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g482 ( .A(n_456), .B(n_460), .Y(n_482) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
OR2x6_ASAP7_75t_L g472 ( .A(n_457), .B(n_467), .Y(n_472) );
INVxp33_ASAP7_75t_L g523 ( .A(n_457), .Y(n_523) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVxp67_ASAP7_75t_L g556 ( .A(n_463), .Y(n_556) );
NOR2x1p5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_472), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_500) );
INVxp67_ASAP7_75t_L g547 ( .A(n_472), .Y(n_547) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_473), .A2(n_518), .B(n_526), .Y(n_517) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_473), .A2(n_518), .B(n_526), .Y(n_565) );
AND2x2_ASAP7_75t_L g495 ( .A(n_474), .B(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g578 ( .A(n_474), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_474), .B(n_568), .Y(n_582) );
INVx2_ASAP7_75t_L g596 ( .A(n_474), .Y(n_596) );
AND2x4_ASAP7_75t_L g600 ( .A(n_474), .B(n_601), .Y(n_600) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_474), .Y(n_635) );
OR2x2_ASAP7_75t_L g641 ( .A(n_474), .B(n_486), .Y(n_641) );
NOR2x1_ASAP7_75t_SL g670 ( .A(n_474), .B(n_497), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_474), .B(n_744), .Y(n_772) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g558 ( .A(n_482), .Y(n_558) );
AND2x2_ASAP7_75t_L g669 ( .A(n_483), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2x1_ASAP7_75t_L g703 ( .A(n_484), .B(n_496), .Y(n_703) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g511 ( .A(n_486), .Y(n_511) );
INVx2_ASAP7_75t_L g569 ( .A(n_486), .Y(n_569) );
AND2x2_ASAP7_75t_L g592 ( .A(n_486), .B(n_497), .Y(n_592) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_486), .Y(n_619) );
INVx1_ASAP7_75t_L g660 ( .A(n_486), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_510), .Y(n_494) );
AND2x2_ASAP7_75t_L g672 ( .A(n_495), .B(n_567), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_496), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g739 ( .A(n_496), .Y(n_739) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g598 ( .A(n_497), .Y(n_598) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_504), .B(n_509), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_503), .B(n_549), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B1(n_507), .B2(n_508), .Y(n_504) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_510), .A2(n_676), .B(n_680), .C(n_686), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_512), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_SL g722 ( .A(n_512), .Y(n_722) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g644 ( .A(n_514), .B(n_598), .Y(n_644) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_535), .Y(n_515) );
AOI32xp33_ASAP7_75t_L g680 ( .A1(n_516), .A2(n_664), .A3(n_681), .B1(n_682), .B2(n_684), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
INVx2_ASAP7_75t_L g606 ( .A(n_517), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_517), .B(n_538), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_519), .B(n_525), .Y(n_518) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx3_ASAP7_75t_L g618 ( .A(n_527), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_527), .B(n_544), .Y(n_649) );
AND2x2_ASAP7_75t_L g654 ( .A(n_527), .B(n_655), .Y(n_654) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_527), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
OR2x2_ASAP7_75t_L g637 ( .A(n_535), .B(n_638), .Y(n_637) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g588 ( .A(n_536), .B(n_562), .Y(n_588) );
AND2x2_ASAP7_75t_L g737 ( .A(n_536), .B(n_735), .Y(n_737) );
AND2x4_ASAP7_75t_L g536 ( .A(n_537), .B(n_544), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g574 ( .A(n_538), .Y(n_574) );
AND2x4_ASAP7_75t_L g613 ( .A(n_538), .B(n_614), .Y(n_613) );
INVxp67_ASAP7_75t_L g647 ( .A(n_538), .Y(n_647) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_538), .Y(n_655) );
AND2x2_ASAP7_75t_L g664 ( .A(n_538), .B(n_544), .Y(n_664) );
INVx1_ASAP7_75t_L g748 ( .A(n_538), .Y(n_748) );
INVx2_ASAP7_75t_L g585 ( .A(n_544), .Y(n_585) );
INVx1_ASAP7_75t_L g612 ( .A(n_544), .Y(n_612) );
INVx1_ASAP7_75t_L g679 ( .A(n_544), .Y(n_679) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_552), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI32xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_570), .A3(n_575), .B1(n_579), .B2(n_583), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_561), .B(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_566), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_562), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g663 ( .A(n_562), .B(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g688 ( .A(n_562), .Y(n_688) );
AND2x2_ASAP7_75t_L g769 ( .A(n_562), .B(n_611), .Y(n_769) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g584 ( .A(n_564), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g683 ( .A(n_564), .B(n_606), .Y(n_683) );
NOR2xp67_ASAP7_75t_L g705 ( .A(n_564), .B(n_585), .Y(n_705) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_564), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g614 ( .A(n_565), .Y(n_614) );
INVx1_ASAP7_75t_L g638 ( .A(n_565), .Y(n_638) );
AND2x2_ASAP7_75t_L g653 ( .A(n_565), .B(n_585), .Y(n_653) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g681 ( .A(n_567), .B(n_670), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_567), .B(n_600), .Y(n_751) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_568), .Y(n_720) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_569), .Y(n_702) );
INVxp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g603 ( .A(n_572), .B(n_604), .Y(n_603) );
NOR2xp67_ASAP7_75t_L g687 ( .A(n_572), .B(n_688), .Y(n_687) );
NOR2xp67_ASAP7_75t_SL g774 ( .A(n_572), .B(n_712), .Y(n_774) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g631 ( .A(n_574), .B(n_585), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_575), .B(n_641), .Y(n_699) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_SL g665 ( .A(n_576), .B(n_592), .Y(n_665) );
AND2x4_ASAP7_75t_SL g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NOR2x1_ASAP7_75t_L g624 ( .A(n_578), .B(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g730 ( .A(n_578), .B(n_601), .Y(n_730) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_578), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_579), .B(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
OR2x2_ASAP7_75t_L g701 ( .A(n_580), .B(n_702), .Y(n_701) );
NOR2x1_ASAP7_75t_L g766 ( .A(n_580), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g690 ( .A(n_581), .B(n_635), .Y(n_690) );
INVxp33_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g604 ( .A(n_584), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g764 ( .A(n_584), .B(n_646), .Y(n_764) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_607), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .B(n_602), .Y(n_590) );
AND2x2_ASAP7_75t_L g725 ( .A(n_592), .B(n_600), .Y(n_725) );
NAND2xp33_ASAP7_75t_R g593 ( .A(n_594), .B(n_599), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g767 ( .A(n_596), .Y(n_767) );
INVx4_ASAP7_75t_L g625 ( .A(n_597), .Y(n_625) );
INVx1_ASAP7_75t_L g744 ( .A(n_598), .Y(n_744) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g738 ( .A(n_600), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_SL g742 ( .A(n_600), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_603), .A2(n_668), .B1(n_772), .B2(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g632 ( .A(n_606), .B(n_618), .Y(n_632) );
AND2x2_ASAP7_75t_L g646 ( .A(n_606), .B(n_647), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_615), .B(n_620), .C(n_623), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g694 ( .A(n_610), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g622 ( .A(n_611), .Y(n_622) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g682 ( .A(n_612), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g691 ( .A(n_612), .B(n_613), .Y(n_691) );
INVx1_ASAP7_75t_L g723 ( .A(n_612), .Y(n_723) );
AND2x4_ASAP7_75t_L g704 ( .A(n_613), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g726 ( .A(n_613), .B(n_617), .Y(n_726) );
AND2x2_ASAP7_75t_L g734 ( .A(n_613), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g709 ( .A(n_617), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_617), .B(n_631), .Y(n_711) );
AND2x2_ASAP7_75t_L g714 ( .A(n_617), .B(n_664), .Y(n_714) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_618), .B(n_679), .Y(n_728) );
AND2x2_ASAP7_75t_L g656 ( .A(n_619), .B(n_644), .Y(n_656) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g752 ( .A(n_622), .B(n_632), .Y(n_752) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_624), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g636 ( .A(n_625), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_625), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_666), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_650), .Y(n_627) );
OAI222xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_633), .B1(n_637), .B2(n_639), .C1(n_642), .C2(n_645), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_635), .B(n_644), .Y(n_643) );
OR2x6_ASAP7_75t_L g715 ( .A(n_635), .B(n_685), .Y(n_715) );
NAND5xp2_ASAP7_75t_L g718 ( .A(n_635), .B(n_638), .C(n_654), .D(n_719), .E(n_721), .Y(n_718) );
NAND2x1_ASAP7_75t_L g754 ( .A(n_636), .B(n_640), .Y(n_754) );
INVx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_641), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_643), .A2(n_734), .B1(n_737), .B2(n_738), .Y(n_733) );
INVx2_ASAP7_75t_L g685 ( .A(n_644), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_644), .B(n_660), .Y(n_697) );
INVx3_ASAP7_75t_L g732 ( .A(n_645), .Y(n_732) );
NAND2x1p5_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
AND2x2_ASAP7_75t_L g677 ( .A(n_646), .B(n_678), .Y(n_677) );
BUFx2_ASAP7_75t_L g710 ( .A(n_646), .Y(n_710) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g673 ( .A(n_649), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_651), .B(n_662), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_656), .B(n_657), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g661 ( .A(n_653), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_656), .A2(n_663), .B1(n_664), .B2(n_665), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .Y(n_657) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x4_ASAP7_75t_SL g743 ( .A(n_660), .B(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_675), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B(n_673), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g712 ( .A(n_683), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_686) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_716), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_698), .C(n_706), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OA21x2_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_700), .B(n_704), .Y(n_698) );
NAND2xp33_ASAP7_75t_SL g700 ( .A(n_701), .B(n_703), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_713), .B(n_715), .Y(n_706) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_711), .C(n_712), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_710), .A2(n_750), .B1(n_752), .B2(n_753), .Y(n_749) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_740), .Y(n_716) );
NAND4xp25_ASAP7_75t_L g717 ( .A(n_718), .B(n_724), .C(n_731), .D(n_733), .Y(n_717) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g729 ( .A(n_720), .B(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVx1_ASAP7_75t_L g760 ( .A(n_723), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B1(n_727), .B2(n_729), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_729), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI21xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_745), .B(n_749), .Y(n_740) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_770), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_760), .B(n_761), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_765), .B2(n_768), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
CKINVDCx11_ASAP7_75t_R g792 ( .A(n_775), .Y(n_792) );
CKINVDCx11_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_778), .Y(n_796) );
INVx1_ASAP7_75t_L g789 ( .A(n_779), .Y(n_789) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B(n_797), .Y(n_788) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
INVx4_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
INVx3_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_803), .B(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
OR2x2_ASAP7_75t_SL g804 ( .A(n_805), .B(n_807), .Y(n_804) );
CKINVDCx16_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
endmodule