module fake_jpeg_25224_n_159 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_17),
.B(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_21),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_59),
.B1(n_53),
.B2(n_65),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_86),
.B1(n_85),
.B2(n_18),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_59),
.B1(n_53),
.B2(n_54),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_46),
.B1(n_55),
.B2(n_73),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_88),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_67),
.B1(n_48),
.B2(n_65),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_86),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_50),
.B1(n_51),
.B2(n_63),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_66),
.B1(n_64),
.B2(n_58),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_95),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_62),
.B1(n_52),
.B2(n_60),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_98),
.B1(n_103),
.B2(n_104),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_61),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_101),
.B(n_105),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

BUFx2_ASAP7_75t_SL g111 ( 
.A(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_0),
.Y(n_101)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_13),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_26),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_15),
.C(n_40),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_104),
.C(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_103),
.B1(n_94),
.B2(n_102),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_108),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_93),
.B1(n_12),
.B2(n_20),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_93),
.B1(n_42),
.B2(n_39),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_38),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_37),
.B(n_32),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_123),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_133),
.B1(n_135),
.B2(n_138),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_132),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_109),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_1),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_30),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_125),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_130),
.Y(n_147)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_146),
.B(n_2),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_29),
.B1(n_28),
.B2(n_22),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_149),
.B1(n_139),
.B2(n_143),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_134),
.B1(n_132),
.B2(n_146),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_142),
.B(n_128),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_141),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_148),
.B1(n_127),
.B2(n_140),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_154),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_5),
.B(n_6),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_5),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_7),
.Y(n_159)
);


endmodule