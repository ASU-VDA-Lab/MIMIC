module fake_jpeg_17543_n_373 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_373);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_373;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_51),
.Y(n_75)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_56),
.Y(n_80)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_18),
.B(n_13),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_23),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_60),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_27),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_96)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_17),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_94),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_39),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_73),
.A2(n_78),
.B1(n_88),
.B2(n_90),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_108),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_83),
.B(n_1),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_46),
.A2(n_27),
.B1(n_25),
.B2(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_41),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_44),
.A2(n_31),
.B1(n_35),
.B2(n_34),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_114),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_54),
.B1(n_51),
.B2(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_35),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_38),
.A2(n_33),
.B1(n_14),
.B2(n_29),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_36),
.B1(n_32),
.B2(n_30),
.Y(n_100)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_42),
.A2(n_33),
.B1(n_14),
.B2(n_16),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_110),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_48),
.B(n_28),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx6p67_ASAP7_75t_R g159 ( 
.A(n_109),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_16),
.B1(n_36),
.B2(n_20),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_52),
.B(n_20),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_20),
.C(n_47),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_55),
.A2(n_36),
.B1(n_20),
.B2(n_17),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_17),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_86),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_121),
.A2(n_71),
.B1(n_118),
.B2(n_117),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_128),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_80),
.B(n_17),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_124),
.B(n_145),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_75),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_135),
.Y(n_174)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_67),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_132),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_68),
.C(n_65),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_70),
.B1(n_101),
.B2(n_77),
.Y(n_176)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_67),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_76),
.B(n_1),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_155),
.Y(n_194)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_87),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_154),
.Y(n_180)
);

BUFx4f_ASAP7_75t_SL g152 ( 
.A(n_81),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_152),
.Y(n_170)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_87),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_17),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_158),
.Y(n_196)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_17),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_67),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_95),
.B(n_1),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_72),
.B(n_92),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_168),
.B(n_4),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_76),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_183),
.Y(n_220)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_193),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_184),
.B1(n_147),
.B2(n_143),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_101),
.B1(n_85),
.B2(n_100),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_182),
.A2(n_202),
.B1(n_210),
.B2(n_148),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_90),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_136),
.A2(n_107),
.B1(n_40),
.B2(n_112),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_2),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_185),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_120),
.B(n_3),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_191),
.Y(n_236)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

INVxp33_ASAP7_75t_SL g229 ( 
.A(n_195),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_120),
.A2(n_3),
.B(n_4),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_212),
.B(n_8),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_126),
.A2(n_118),
.B1(n_117),
.B2(n_109),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_204),
.Y(n_249)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_237)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_126),
.A2(n_104),
.B1(n_89),
.B2(n_82),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_145),
.A2(n_5),
.B(n_7),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_119),
.A2(n_71),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_161),
.B(n_142),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_197),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_248),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_127),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_222),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_130),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_221),
.A2(n_243),
.B(n_209),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_135),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_149),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_231),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_232),
.B1(n_210),
.B2(n_202),
.Y(n_264)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_200),
.A2(n_149),
.B(n_139),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_227),
.A2(n_237),
.B(n_238),
.Y(n_267)
);

OAI22x1_ASAP7_75t_L g262 ( 
.A1(n_230),
.A2(n_235),
.B1(n_211),
.B2(n_195),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_180),
.B(n_123),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_138),
.B1(n_133),
.B2(n_148),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_181),
.A2(n_182),
.B1(n_191),
.B2(n_185),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_233),
.A2(n_239),
.B1(n_247),
.B2(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_205),
.A2(n_188),
.B1(n_207),
.B2(n_190),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_81),
.B(n_10),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_181),
.A2(n_158),
.B1(n_125),
.B2(n_131),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_82),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_245),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_187),
.B(n_194),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_198),
.C(n_208),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_199),
.A2(n_159),
.B(n_81),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_242),
.A2(n_246),
.B(n_238),
.Y(n_273)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_244),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_122),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_192),
.A2(n_10),
.B(n_159),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_176),
.A2(n_159),
.B1(n_137),
.B2(n_150),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_169),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_175),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_206),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_173),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_254),
.B(n_255),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_257),
.B(n_275),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_214),
.A2(n_192),
.B(n_190),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_258),
.A2(n_262),
.B(n_273),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_259),
.B(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_278),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_179),
.B1(n_189),
.B2(n_204),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_189),
.B1(n_159),
.B2(n_170),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_170),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_211),
.C(n_177),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_280),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_220),
.B(n_172),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_272),
.C(n_279),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_193),
.Y(n_272)
);

OAI32xp33_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_150),
.A3(n_177),
.B1(n_228),
.B2(n_240),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_274),
.A2(n_277),
.B(n_263),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_231),
.B(n_215),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_229),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_249),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_228),
.B(n_236),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_221),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_227),
.C(n_217),
.Y(n_280)
);

OAI22x1_ASAP7_75t_SL g282 ( 
.A1(n_230),
.A2(n_237),
.B1(n_242),
.B2(n_226),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_245),
.B1(n_218),
.B2(n_239),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_234),
.B(n_233),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_298),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_285),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_257),
.B(n_215),
.Y(n_290)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_290),
.A2(n_301),
.B(n_288),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_299),
.B1(n_307),
.B2(n_309),
.Y(n_310)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_263),
.A2(n_218),
.B1(n_247),
.B2(n_251),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_296),
.A2(n_309),
.B1(n_291),
.B2(n_298),
.Y(n_320)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_219),
.B(n_251),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_300),
.A2(n_303),
.B(n_305),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_250),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_252),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_306),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_267),
.A2(n_283),
.B(n_276),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_253),
.B(n_249),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_274),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_279),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_317),
.C(n_318),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_264),
.B1(n_266),
.B2(n_278),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_312),
.A2(n_316),
.B1(n_323),
.B2(n_328),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_304),
.A2(n_280),
.B1(n_261),
.B2(n_270),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_313),
.A2(n_314),
.B1(n_284),
.B2(n_300),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_261),
.B1(n_268),
.B2(n_267),
.Y(n_314)
);

OAI22x1_ASAP7_75t_L g315 ( 
.A1(n_293),
.A2(n_271),
.B1(n_272),
.B2(n_249),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_290),
.B1(n_293),
.B2(n_289),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_268),
.B1(n_255),
.B2(n_254),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_256),
.C(n_223),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_223),
.Y(n_318)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

OAI322xp33_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_286),
.A3(n_288),
.B1(n_294),
.B2(n_296),
.C1(n_302),
.C2(n_315),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_295),
.C(n_292),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_328),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_303),
.C(n_305),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_331),
.Y(n_353)
);

NAND4xp25_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_340),
.C(n_317),
.D(n_311),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_321),
.A2(n_319),
.B(n_322),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_334),
.A2(n_341),
.B(n_342),
.Y(n_346)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_325),
.Y(n_336)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_337),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_321),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_338),
.B(n_339),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_324),
.B(n_286),
.Y(n_339)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_310),
.B(n_314),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_324),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_343),
.B(n_313),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_341),
.A2(n_320),
.B(n_327),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_344),
.A2(n_347),
.B1(n_332),
.B2(n_336),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_340),
.C(n_339),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_318),
.C(n_335),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_352),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_330),
.C(n_343),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_334),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_340),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_349),
.A2(n_338),
.B1(n_332),
.B2(n_333),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_357),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_356),
.A2(n_346),
.B(n_337),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g357 ( 
.A(n_351),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_353),
.C(n_346),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_354),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_363),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_362),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_364),
.B(n_348),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_367),
.Y(n_369)
);

AOI322xp5_ASAP7_75t_L g368 ( 
.A1(n_366),
.A2(n_344),
.A3(n_358),
.B1(n_345),
.B2(n_356),
.C1(n_363),
.C2(n_342),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_368),
.A2(n_365),
.B(n_353),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_370),
.A2(n_369),
.B(n_352),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_371),
.B(n_350),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_372),
.A2(n_347),
.B(n_357),
.Y(n_373)
);


endmodule