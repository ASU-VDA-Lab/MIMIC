module fake_jpeg_2060_n_623 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_623);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_623;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_10),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_11),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_58),
.B(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_63),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_64),
.B(n_81),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_68),
.Y(n_186)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g179 ( 
.A(n_69),
.Y(n_179)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_70),
.Y(n_188)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_72),
.Y(n_198)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_75),
.Y(n_214)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_78),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_80),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_19),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_87),
.Y(n_210)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_92),
.Y(n_142)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_24),
.B(n_11),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_36),
.B(n_10),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_98),
.Y(n_145)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_31),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_99),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_101),
.Y(n_222)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_103),
.B(n_107),
.Y(n_213)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_22),
.Y(n_106)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_28),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_108),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

BUFx4f_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_31),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_114),
.B(n_125),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_116),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_23),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_119),
.B(n_106),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_39),
.B(n_10),
.Y(n_120)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_44),
.B(n_12),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_128),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_44),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_28),
.Y(n_126)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_31),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_127),
.B(n_4),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_37),
.B(n_18),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_32),
.Y(n_129)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_70),
.A2(n_48),
.B1(n_41),
.B2(n_45),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_133),
.A2(n_137),
.B1(n_205),
.B2(n_207),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_57),
.B1(n_55),
.B2(n_32),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_135),
.A2(n_153),
.B1(n_167),
.B2(n_173),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_73),
.B(n_37),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_136),
.B(n_172),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_48),
.B1(n_45),
.B2(n_41),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_63),
.A2(n_57),
.B1(n_41),
.B2(n_45),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_146),
.A2(n_149),
.B1(n_155),
.B2(n_169),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_51),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_148),
.B(n_159),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_102),
.A2(n_45),
.B1(n_51),
.B2(n_50),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_69),
.A2(n_57),
.B1(n_56),
.B2(n_43),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_66),
.A2(n_20),
.B1(n_56),
.B2(n_50),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_49),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g283 ( 
.A(n_162),
.B(n_163),
.CON(n_283),
.SN(n_283)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_86),
.B(n_20),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_100),
.A2(n_55),
.B1(n_32),
.B2(n_20),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_67),
.A2(n_49),
.B1(n_46),
.B2(n_43),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_68),
.B(n_100),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_171),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_68),
.B(n_46),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_105),
.A2(n_55),
.B1(n_32),
.B2(n_27),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_113),
.B(n_55),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_176),
.B(n_178),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_87),
.B(n_113),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_72),
.A2(n_27),
.B1(n_48),
.B2(n_32),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_182),
.A2(n_200),
.B1(n_96),
.B2(n_93),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_88),
.A2(n_55),
.B1(n_27),
.B2(n_54),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_183),
.A2(n_193),
.B1(n_204),
.B2(n_216),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_75),
.B(n_13),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_184),
.B(n_199),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_91),
.A2(n_27),
.B1(n_54),
.B2(n_13),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_109),
.A2(n_27),
.B1(n_54),
.B2(n_2),
.Y(n_194)
);

AOI22x1_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_224),
.B1(n_90),
.B2(n_1),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_82),
.B(n_13),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_77),
.A2(n_54),
.B1(n_13),
.B2(n_14),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_108),
.A2(n_7),
.B1(n_17),
.B2(n_16),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_84),
.A2(n_8),
.B1(n_17),
.B2(n_16),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_85),
.A2(n_5),
.B1(n_16),
.B2(n_15),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_110),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_218),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_115),
.A2(n_5),
.B1(n_15),
.B2(n_8),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_212),
.A2(n_198),
.B1(n_187),
.B2(n_214),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_121),
.A2(n_124),
.B1(n_116),
.B2(n_118),
.Y(n_216)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_90),
.A2(n_117),
.B1(n_78),
.B2(n_80),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_142),
.B(n_0),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_227),
.B(n_243),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_141),
.B1(n_150),
.B2(n_155),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_228),
.A2(n_240),
.B1(n_285),
.B2(n_295),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_229),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_154),
.B(n_111),
.C(n_97),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_230),
.B(n_263),
.Y(n_321)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_131),
.A2(n_139),
.A3(n_138),
.B1(n_147),
.B2(n_213),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_233),
.B(n_287),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_234),
.A2(n_267),
.B1(n_231),
.B2(n_247),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_215),
.B(n_111),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_236),
.B(n_258),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_238),
.A2(n_276),
.B1(n_284),
.B2(n_300),
.Y(n_342)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_239),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_146),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_166),
.B(n_0),
.Y(n_243)
);

AO22x1_ASAP7_75t_SL g244 ( 
.A1(n_194),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_244)
);

AO22x1_ASAP7_75t_L g310 ( 
.A1(n_244),
.A2(n_234),
.B1(n_284),
.B2(n_255),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_0),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_245),
.B(n_275),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_135),
.A2(n_18),
.B(n_1),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_246),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_171),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_247),
.B(n_264),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_177),
.A2(n_1),
.B1(n_2),
.B2(n_225),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_SL g332 ( 
.A1(n_248),
.A2(n_282),
.B(n_299),
.Y(n_332)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_249),
.Y(n_335)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_251),
.Y(n_324)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_252),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_254),
.Y(n_350)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_255),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_152),
.Y(n_256)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_257),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_145),
.B(n_1),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_199),
.B(n_2),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_260),
.B(n_297),
.Y(n_341)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

INVx11_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_2),
.C(n_221),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_190),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_186),
.Y(n_265)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_143),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_134),
.Y(n_268)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_170),
.Y(n_269)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_132),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_274),
.Y(n_323)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_152),
.Y(n_272)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_175),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_202),
.B(n_194),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_224),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_281),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_224),
.B(n_173),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_278),
.B(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_161),
.Y(n_279)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_279),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_143),
.B(n_191),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_167),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_177),
.A2(n_225),
.B1(n_189),
.B2(n_161),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_182),
.A2(n_183),
.B1(n_193),
.B2(n_144),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_181),
.A2(n_187),
.B1(n_198),
.B2(n_157),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_185),
.B(n_201),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_195),
.B(n_156),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_134),
.B(n_180),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_289),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_158),
.B(n_180),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_196),
.B(n_203),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_158),
.B(n_164),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_292),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_164),
.B(n_195),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_175),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_293),
.B(n_294),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_189),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_157),
.A2(n_214),
.B1(n_188),
.B2(n_206),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_165),
.B(n_210),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_306),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_217),
.B(n_210),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_217),
.B(n_206),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_298),
.B(n_305),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_165),
.A2(n_220),
.B1(n_219),
.B2(n_151),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_130),
.A2(n_144),
.B1(n_151),
.B2(n_160),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_301),
.B(n_304),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_168),
.B(n_130),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_302),
.B(n_256),
.Y(n_351)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_160),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_303),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_168),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_141),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_215),
.Y(n_306)
);

INVx6_ASAP7_75t_SL g307 ( 
.A(n_186),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_307),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_184),
.A2(n_182),
.B1(n_146),
.B2(n_169),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_308),
.A2(n_241),
.B1(n_245),
.B2(n_243),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_310),
.A2(n_322),
.B1(n_325),
.B2(n_343),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_277),
.A2(n_231),
.B1(n_308),
.B2(n_275),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_315),
.A2(n_330),
.B1(n_346),
.B2(n_348),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_226),
.A2(n_235),
.B1(n_276),
.B2(n_237),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_226),
.A2(n_281),
.B1(n_253),
.B2(n_238),
.Y(n_330)
);

OAI32xp33_ASAP7_75t_L g333 ( 
.A1(n_241),
.A2(n_253),
.A3(n_271),
.B1(n_232),
.B2(n_233),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_333),
.B(n_351),
.Y(n_374)
);

O2A1O1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_283),
.A2(n_238),
.B(n_278),
.C(n_244),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_337),
.A2(n_269),
.B(n_272),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_267),
.A2(n_302),
.B1(n_246),
.B2(n_244),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_300),
.A2(n_274),
.B1(n_305),
.B2(n_290),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_271),
.A2(n_263),
.B1(n_244),
.B2(n_259),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_353),
.A2(n_363),
.B1(n_297),
.B2(n_251),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_258),
.B(n_260),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_361),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_260),
.B(n_227),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_232),
.A2(n_230),
.B1(n_288),
.B2(n_289),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_307),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_257),
.Y(n_371)
);

AO22x1_ASAP7_75t_SL g368 ( 
.A1(n_342),
.A2(n_293),
.B1(n_250),
.B2(n_273),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_368),
.B(n_377),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_330),
.A2(n_322),
.B1(n_326),
.B2(n_311),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_370),
.A2(n_329),
.B1(n_362),
.B2(n_352),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_270),
.C(n_236),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_373),
.C(n_399),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_306),
.C(n_291),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_323),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_382),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_292),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_356),
.Y(n_378)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_298),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_387),
.Y(n_426)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_312),
.Y(n_383)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_384),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_347),
.Y(n_385)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_357),
.B(n_264),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_386),
.B(n_391),
.Y(n_432)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_318),
.B(n_242),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_388),
.B(n_392),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_262),
.B1(n_242),
.B2(n_256),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_389),
.A2(n_394),
.B1(n_401),
.B2(n_358),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_352),
.A2(n_294),
.B1(n_297),
.B2(n_229),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_390),
.A2(n_410),
.B1(n_316),
.B2(n_365),
.Y(n_416)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_367),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_318),
.B(n_239),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_396),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_310),
.A2(n_304),
.B1(n_279),
.B2(n_301),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_344),
.A2(n_249),
.B1(n_268),
.B2(n_252),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_395),
.A2(n_397),
.B(n_406),
.Y(n_443)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_338),
.B(n_272),
.Y(n_398)
);

A2O1A1O1Ixp25_ASAP7_75t_L g424 ( 
.A1(n_398),
.A2(n_403),
.B(n_413),
.C(n_354),
.D(n_337),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_311),
.B(n_265),
.C(n_261),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_261),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_400),
.B(n_402),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_310),
.A2(n_261),
.B1(n_303),
.B2(n_325),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_323),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_338),
.B(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_404),
.A2(n_405),
.B1(n_411),
.B2(n_412),
.Y(n_430)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_344),
.B(n_346),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_363),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_341),
.C(n_358),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_319),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_408),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_361),
.B(n_319),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_409),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_340),
.B(n_359),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_366),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_313),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_353),
.B(n_359),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_416),
.A2(n_395),
.B(n_411),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_341),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_422),
.C(n_423),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_421),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_333),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_375),
.B(n_341),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_450),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_427),
.B(n_380),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_369),
.A2(n_329),
.B1(n_341),
.B2(n_316),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_428),
.A2(n_436),
.B1(n_437),
.B2(n_439),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_441),
.C(n_445),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_380),
.A2(n_332),
.B1(n_331),
.B2(n_366),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_431),
.A2(n_394),
.B1(n_377),
.B2(n_410),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_376),
.A2(n_402),
.B1(n_397),
.B2(n_378),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_372),
.B(n_350),
.C(n_317),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_438),
.C(n_440),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_369),
.A2(n_406),
.B1(n_379),
.B2(n_401),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_406),
.A2(n_331),
.B1(n_328),
.B2(n_313),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_350),
.C(n_317),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_389),
.A2(n_328),
.B1(n_334),
.B2(n_335),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_339),
.C(n_324),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_370),
.B(n_327),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_382),
.A2(n_334),
.B1(n_335),
.B2(n_327),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_444),
.A2(n_387),
.B1(n_396),
.B2(n_383),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_399),
.B(n_339),
.C(n_324),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_381),
.A2(n_347),
.B1(n_345),
.B2(n_355),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_393),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_456),
.B(n_464),
.Y(n_503)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_425),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_460),
.Y(n_504)
);

AOI32xp33_ASAP7_75t_L g461 ( 
.A1(n_414),
.A2(n_443),
.A3(n_449),
.B1(n_374),
.B2(n_415),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_461),
.B(n_462),
.Y(n_500)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_463),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_452),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_465),
.A2(n_466),
.B1(n_484),
.B2(n_485),
.Y(n_501)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_447),
.Y(n_467)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_467),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_446),
.Y(n_468)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_432),
.Y(n_469)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_443),
.A2(n_374),
.B(n_371),
.Y(n_470)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_470),
.A2(n_478),
.B(n_426),
.Y(n_492)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_471),
.Y(n_510)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_472),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_416),
.A2(n_398),
.B(n_405),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_473),
.B(n_423),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_436),
.A2(n_409),
.B1(n_368),
.B2(n_388),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_474),
.A2(n_426),
.B1(n_431),
.B2(n_427),
.Y(n_491)
);

NOR2x1_ASAP7_75t_L g475 ( 
.A(n_415),
.B(n_375),
.Y(n_475)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_475),
.Y(n_516)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_477),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_428),
.A2(n_391),
.B(n_368),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_433),
.B(n_412),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_480),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_368),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_481),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_417),
.B(n_404),
.C(n_384),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_417),
.C(n_435),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_449),
.B(n_420),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_483),
.B(n_486),
.Y(n_494)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_418),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_433),
.B(n_392),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_487),
.A2(n_488),
.B1(n_420),
.B2(n_444),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_437),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_489),
.B(n_496),
.C(n_512),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_419),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_490),
.B(n_511),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_491),
.A2(n_519),
.B1(n_464),
.B2(n_481),
.Y(n_544)
);

BUFx4f_ASAP7_75t_SL g528 ( 
.A(n_492),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_438),
.C(n_429),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_454),
.B(n_422),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_506),
.B(n_515),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_507),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_457),
.A2(n_441),
.B1(n_421),
.B2(n_440),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_508),
.A2(n_509),
.B1(n_514),
.B2(n_521),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_457),
.A2(n_439),
.B1(n_424),
.B2(n_445),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_453),
.B(n_451),
.C(n_355),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_457),
.A2(n_451),
.B1(n_385),
.B2(n_309),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_454),
.B(n_309),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_453),
.B(n_314),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_517),
.B(n_518),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_453),
.B(n_459),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_474),
.A2(n_314),
.B1(n_336),
.B2(n_479),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_465),
.A2(n_488),
.B1(n_479),
.B2(n_466),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_493),
.B(n_483),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_523),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_490),
.B(n_470),
.C(n_476),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_525),
.B(n_506),
.C(n_511),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_499),
.B(n_468),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_526),
.B(n_527),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_486),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_521),
.A2(n_520),
.B1(n_509),
.B2(n_501),
.Y(n_529)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_529),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_473),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_530),
.B(n_531),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_496),
.B(n_455),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_505),
.B(n_469),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_532),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_517),
.B(n_455),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_533),
.B(n_537),
.C(n_547),
.Y(n_554)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_495),
.Y(n_534)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_534),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_SL g535 ( 
.A(n_500),
.B(n_516),
.C(n_513),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_536),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_512),
.B(n_461),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_489),
.B(n_462),
.Y(n_537)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_540),
.Y(n_552)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_503),
.Y(n_541)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_541),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_519),
.A2(n_478),
.B(n_471),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_543),
.A2(n_507),
.B(n_492),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_544),
.A2(n_501),
.B1(n_508),
.B2(n_498),
.Y(n_553)
);

NAND2xp67_ASAP7_75t_SL g545 ( 
.A(n_492),
.B(n_477),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_545),
.A2(n_544),
.B(n_475),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_515),
.B(n_472),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_549),
.B(n_546),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_551),
.A2(n_563),
.B(n_528),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_553),
.A2(n_529),
.B1(n_542),
.B2(n_528),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_543),
.A2(n_475),
.B(n_491),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_555),
.A2(n_535),
.B(n_510),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_522),
.B(n_494),
.C(n_504),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_560),
.B(n_561),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_522),
.B(n_504),
.C(n_502),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_545),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_562),
.B(n_566),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_539),
.B(n_502),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_565),
.Y(n_578)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_528),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_546),
.B(n_480),
.C(n_456),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_567),
.B(n_531),
.C(n_533),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_569),
.B(n_572),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_570),
.A2(n_580),
.B1(n_582),
.B2(n_563),
.Y(n_593)
);

MAJx2_ASAP7_75t_L g571 ( 
.A(n_549),
.B(n_538),
.C(n_530),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_571),
.B(n_574),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_559),
.B(n_537),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_573),
.A2(n_579),
.B(n_555),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_525),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_575),
.B(n_576),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_561),
.B(n_524),
.C(n_538),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_568),
.A2(n_547),
.B1(n_514),
.B2(n_485),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_568),
.A2(n_484),
.B1(n_524),
.B2(n_497),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_554),
.B(n_458),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_460),
.C(n_463),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_584),
.B(n_551),
.C(n_553),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_586),
.B(n_587),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_581),
.B(n_564),
.C(n_554),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_577),
.Y(n_588)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_588),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_573),
.B(n_566),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_590),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_575),
.B(n_554),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_591),
.B(n_592),
.Y(n_607)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_582),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_593),
.A2(n_595),
.B1(n_580),
.B2(n_552),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_584),
.A2(n_550),
.B(n_559),
.Y(n_594)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_594),
.A2(n_550),
.B(n_558),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_578),
.A2(n_562),
.B(n_565),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_597),
.A2(n_552),
.B(n_557),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_598),
.B(n_603),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_601),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_585),
.A2(n_583),
.B(n_569),
.Y(n_601)
);

NAND2xp67_ASAP7_75t_SL g604 ( 
.A(n_597),
.B(n_557),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_604),
.B(n_606),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g606 ( 
.A1(n_595),
.A2(n_558),
.B(n_571),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_602),
.B(n_556),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_608),
.B(n_612),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_599),
.B(n_556),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_605),
.B(n_587),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_613),
.B(n_591),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_611),
.A2(n_607),
.B(n_604),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_614),
.B(n_610),
.Y(n_618)
);

NAND4xp25_ASAP7_75t_L g615 ( 
.A(n_609),
.B(n_589),
.C(n_603),
.D(n_570),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g619 ( 
.A(n_615),
.B(n_617),
.C(n_609),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_618),
.A2(n_619),
.B(n_616),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_620),
.A2(n_590),
.B1(n_593),
.B2(n_548),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_621),
.A2(n_590),
.B(n_586),
.Y(n_622)
);

NAND2x1_ASAP7_75t_L g623 ( 
.A(n_622),
.B(n_596),
.Y(n_623)
);


endmodule