module fake_jpeg_11864_n_183 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_43),
.B1(n_30),
.B2(n_16),
.Y(n_52)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_4),
.Y(n_56)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_42),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_24),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_61),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_59),
.B1(n_27),
.B2(n_31),
.Y(n_73)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_30),
.B1(n_18),
.B2(n_36),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_16),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_29),
.C(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_17),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_17),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_83),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_68),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_19),
.B(n_32),
.C(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_79),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_37),
.B1(n_40),
.B2(n_35),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_67),
.A2(n_69),
.B1(n_77),
.B2(n_16),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_40),
.B1(n_31),
.B2(n_29),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_38),
.Y(n_70)
);

XNOR2x1_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_38),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_78),
.B1(n_58),
.B2(n_56),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_27),
.B1(n_18),
.B2(n_19),
.Y(n_78)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_12),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_32),
.C(n_22),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_16),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_56),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_102),
.B(n_50),
.C(n_48),
.D(n_7),
.Y(n_122)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_46),
.B1(n_54),
.B2(n_51),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_100),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_22),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_72),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_81),
.B1(n_68),
.B2(n_63),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_66),
.B(n_64),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_114),
.B(n_121),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_81),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_118),
.B1(n_94),
.B2(n_8),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_69),
.B1(n_67),
.B2(n_77),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_115),
.B1(n_89),
.B2(n_88),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_80),
.Y(n_113)
);

NOR4xp25_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_5),
.C(n_6),
.D(n_8),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_85),
.A2(n_46),
.B(n_50),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_92),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_51),
.B1(n_75),
.B2(n_79),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_86),
.B(n_16),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_48),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_85),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_133),
.B1(n_135),
.B2(n_118),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_98),
.B(n_92),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_110),
.B1(n_122),
.B2(n_112),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_125),
.B(n_123),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_95),
.B1(n_99),
.B2(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_132),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_87),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_87),
.B1(n_90),
.B2(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_137),
.B(n_108),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_113),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_145),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_140),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_138),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_114),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_112),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_148),
.C(n_123),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_121),
.C(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_131),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_158),
.B(n_150),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_147),
.B(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_129),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_150),
.C(n_148),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_166),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_153),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_107),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_154),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_145),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_173),
.A3(n_159),
.B1(n_167),
.B2(n_163),
.C1(n_137),
.C2(n_126),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_171),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_126),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_12),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_6),
.C2(n_94),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_168),
.B(n_171),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_159),
.A3(n_142),
.B1(n_135),
.B2(n_105),
.C1(n_121),
.C2(n_14),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_180),
.B(n_9),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_94),
.B(n_9),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_10),
.Y(n_182)
);


endmodule