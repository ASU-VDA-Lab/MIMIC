module fake_netlist_6_2894_n_2311 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2311);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2311;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_2292;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_123),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_37),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_56),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_115),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_208),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_37),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_140),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_220),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_117),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_197),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_125),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_55),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_47),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_113),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_42),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_152),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_105),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_99),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_128),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_217),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_81),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_137),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_209),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_130),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_57),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_9),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_192),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_0),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_106),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_108),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_172),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_46),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_104),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_39),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_44),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_31),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_14),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_215),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_95),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_30),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_31),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_32),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_57),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_127),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_88),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_73),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_188),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_52),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_169),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_87),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_210),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_136),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_39),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_158),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_73),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_89),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_18),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_11),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_221),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_42),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_155),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_101),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_193),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_97),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_5),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_176),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_160),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_33),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_40),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_47),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_143),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_166),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_198),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_148),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_79),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_222),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_82),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_229),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_133),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_88),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_124),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_183),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_153),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_205),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_225),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_56),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_59),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_18),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_211),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_41),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_135),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_77),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_69),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_29),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_175),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_116),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_68),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_141),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_212),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_51),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_44),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_203),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_184),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_168),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_118),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_35),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_48),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_5),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_63),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_75),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_230),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_134),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_29),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_71),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_17),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_103),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_34),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_19),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_214),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_182),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_21),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_35),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_191),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g364 ( 
.A(n_204),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_21),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_146),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_7),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_3),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_84),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_139),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_159),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_151),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_12),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_20),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_22),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_164),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_219),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_16),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_119),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_82),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_180),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_66),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_224),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_11),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_46),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_156),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_122),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_86),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_201),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_14),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_51),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_207),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_171),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_189),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_67),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_77),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_170),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_17),
.Y(n_398)
);

BUFx10_ASAP7_75t_L g399 ( 
.A(n_92),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_216),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_60),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_145),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_69),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_174),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_200),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_231),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_142),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_58),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_24),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_2),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_71),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_181),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_19),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_126),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_111),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_53),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_195),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_65),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_80),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_60),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_40),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_48),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_26),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_199),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_165),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_223),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_0),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_227),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_76),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_61),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_12),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_72),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_2),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_26),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_228),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_102),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_64),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_131),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_138),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_96),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_43),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_75),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_67),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_43),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_63),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_226),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_6),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_129),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_93),
.Y(n_449)
);

INVxp33_ASAP7_75t_SL g450 ( 
.A(n_78),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_58),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_100),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_53),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_121),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_354),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_232),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_255),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_238),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_354),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_397),
.B(n_1),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_244),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_239),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_397),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_243),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_360),
.Y(n_466)
);

BUFx2_ASAP7_75t_SL g467 ( 
.A(n_265),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_381),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_354),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_354),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_354),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_354),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_245),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_354),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_246),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_403),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_434),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_385),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_252),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_354),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_393),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_265),
.B(n_1),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_385),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_256),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_385),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_258),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_263),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_394),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_404),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_263),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_261),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_263),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_263),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_267),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_428),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_268),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_237),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_335),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_335),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_269),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_237),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_364),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_271),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_263),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_276),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_277),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_288),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_430),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_290),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_282),
.B(n_3),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_364),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_385),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_430),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_291),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_293),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_295),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_298),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_302),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_430),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_303),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_310),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_430),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_312),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_313),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_317),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_320),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_322),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_451),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_253),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_451),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_451),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_451),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_323),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_324),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_262),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_262),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_336),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_283),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_338),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_283),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_344),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_342),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_344),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_343),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_282),
.B(n_4),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_371),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_334),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_345),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_351),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_334),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_352),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_418),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_356),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_418),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_359),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_363),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_253),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_280),
.B(n_4),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_285),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_366),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_294),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_371),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_372),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_423),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_376),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_377),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_270),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_383),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_386),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_362),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_500),
.B(n_294),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_463),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_455),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_478),
.B(n_387),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_465),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_541),
.B(n_546),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_505),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_459),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_R g586 ( 
.A(n_464),
.B(n_392),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_490),
.Y(n_587)
);

AND2x2_ASAP7_75t_SL g588 ( 
.A(n_461),
.B(n_242),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_490),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_504),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_493),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_473),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_455),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_493),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_462),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_475),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_548),
.B(n_362),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_479),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_495),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_486),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_489),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_500),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_494),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_497),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_551),
.B(n_280),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_499),
.B(n_387),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_484),
.B(n_285),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_506),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_567),
.B(n_234),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_488),
.B(n_318),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_508),
.B(n_318),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_456),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_456),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_510),
.B(n_379),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_460),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_567),
.B(n_234),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_495),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_496),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_512),
.Y(n_619)
);

BUFx8_ASAP7_75t_L g620 ( 
.A(n_485),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_466),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_519),
.Y(n_622)
);

CKINVDCx16_ASAP7_75t_R g623 ( 
.A(n_501),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_496),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_520),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_521),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_SL g628 ( 
.A(n_487),
.B(n_289),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_507),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_522),
.B(n_379),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_524),
.B(n_389),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_525),
.B(n_531),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_507),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_R g634 ( 
.A(n_503),
.B(n_400),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_511),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_511),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_469),
.B(n_247),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_515),
.B(n_389),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_468),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_539),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_516),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_516),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_544),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_547),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_517),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_540),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_502),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_517),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_549),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_467),
.B(n_450),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_568),
.B(n_289),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_553),
.B(n_242),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_523),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_523),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_554),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_556),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_526),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_469),
.A2(n_301),
.B(n_249),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_526),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_532),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_532),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_558),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_561),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_533),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_470),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_535),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_535),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_536),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_536),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_537),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_566),
.Y(n_672)
);

NOR2xp67_ASAP7_75t_L g673 ( 
.A(n_470),
.B(n_471),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_584),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_584),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_584),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_584),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_589),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_583),
.B(n_569),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_593),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_637),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_650),
.B(n_571),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_583),
.B(n_605),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_611),
.B(n_576),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_607),
.B(n_467),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_586),
.B(n_509),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_580),
.Y(n_687)
);

OR2x6_ASAP7_75t_L g688 ( 
.A(n_632),
.B(n_341),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_589),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_593),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_607),
.B(n_537),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_607),
.B(n_457),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_603),
.B(n_518),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_646),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_646),
.Y(n_695)
);

AND2x2_ASAP7_75t_SL g696 ( 
.A(n_588),
.B(n_482),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_603),
.B(n_527),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_603),
.B(n_528),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_580),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_614),
.B(n_529),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_630),
.B(n_530),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_645),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_658),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_642),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_631),
.B(n_538),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_615),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_603),
.B(n_542),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_609),
.B(n_341),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_645),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_616),
.B(n_429),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_607),
.B(n_610),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_657),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_610),
.B(n_458),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_610),
.B(n_540),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_605),
.B(n_651),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_651),
.B(n_540),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_642),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_606),
.B(n_560),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_602),
.B(n_429),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_610),
.B(n_577),
.Y(n_721)
);

AND2x2_ASAP7_75t_SL g722 ( 
.A(n_588),
.B(n_513),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_593),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_638),
.B(n_577),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_657),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_659),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_659),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_615),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_588),
.A2(n_550),
.B1(n_485),
.B2(n_477),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_579),
.B(n_575),
.Y(n_730)
);

INVx6_ASAP7_75t_L g731 ( 
.A(n_581),
.Y(n_731)
);

INVx4_ASAP7_75t_SL g732 ( 
.A(n_637),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_593),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_578),
.A2(n_572),
.B1(n_483),
.B2(n_476),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_612),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_642),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_652),
.B(n_564),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_638),
.A2(n_563),
.B1(n_433),
.B2(n_270),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_615),
.Y(n_739)
);

INVx4_ASAP7_75t_L g740 ( 
.A(n_642),
.Y(n_740)
);

BUFx10_ASAP7_75t_L g741 ( 
.A(n_582),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_612),
.Y(n_742)
);

OR2x6_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_563),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_612),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_638),
.B(n_543),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_592),
.B(n_564),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_638),
.B(n_471),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_646),
.B(n_472),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_597),
.B(n_543),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_581),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_581),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_666),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_596),
.B(n_564),
.Y(n_753)
);

BUFx10_ASAP7_75t_L g754 ( 
.A(n_598),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_581),
.B(n_545),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_612),
.A2(n_272),
.B1(n_284),
.B2(n_281),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_587),
.B(n_545),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_642),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_613),
.B(n_472),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_613),
.B(n_626),
.Y(n_760)
);

INVxp33_ASAP7_75t_SL g761 ( 
.A(n_634),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_590),
.B(n_534),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_600),
.B(n_481),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_666),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_658),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_642),
.Y(n_766)
);

OR2x6_ASAP7_75t_L g767 ( 
.A(n_647),
.B(n_562),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_613),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_666),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_613),
.B(n_474),
.Y(n_770)
);

AND2x6_ASAP7_75t_L g771 ( 
.A(n_626),
.B(n_249),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_587),
.B(n_552),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_626),
.A2(n_281),
.B1(n_284),
.B2(n_272),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_626),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_591),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_591),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_601),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_594),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_604),
.B(n_491),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_637),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_L g781 ( 
.A(n_637),
.B(n_364),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_594),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_661),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_661),
.Y(n_784)
);

INVx4_ASAP7_75t_SL g785 ( 
.A(n_637),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_661),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_599),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_647),
.B(n_574),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_599),
.B(n_552),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_617),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_608),
.B(n_234),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_619),
.B(n_492),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_622),
.B(n_625),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_620),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_673),
.B(n_474),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_628),
.A2(n_498),
.B1(n_300),
.B2(n_311),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_617),
.B(n_555),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_620),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_627),
.B(n_640),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_585),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_643),
.B(n_234),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_644),
.B(n_399),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_661),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_673),
.A2(n_287),
.B1(n_292),
.B2(n_286),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_618),
.B(n_573),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_649),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_618),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_655),
.B(n_382),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_656),
.B(n_236),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_661),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_670),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_637),
.A2(n_287),
.B1(n_292),
.B2(n_286),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_595),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_624),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_624),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_670),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_662),
.B(n_248),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_629),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_629),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_637),
.A2(n_308),
.B1(n_316),
.B2(n_314),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_664),
.B(n_250),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_672),
.B(n_251),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_620),
.B(n_399),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_633),
.B(n_480),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_633),
.B(n_635),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_635),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_636),
.B(n_301),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_623),
.B(n_264),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_620),
.B(n_399),
.Y(n_829)
);

BUFx10_ASAP7_75t_L g830 ( 
.A(n_636),
.Y(n_830)
);

AND3x2_ASAP7_75t_L g831 ( 
.A(n_641),
.B(n_235),
.C(n_233),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_641),
.B(n_364),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_695),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_771),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_751),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_750),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_675),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_775),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_712),
.B(n_247),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_751),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_767),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_696),
.B(n_247),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_696),
.B(n_247),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_675),
.B(n_648),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_750),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_755),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_722),
.A2(n_235),
.B1(n_254),
.B2(n_233),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_675),
.B(n_648),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_676),
.B(n_653),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_722),
.A2(n_254),
.B1(n_260),
.B2(n_257),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_749),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_676),
.B(n_653),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_679),
.B(n_390),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_676),
.B(n_654),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_683),
.B(n_654),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_716),
.B(n_623),
.Y(n_856)
);

AOI221xp5_ASAP7_75t_L g857 ( 
.A1(n_729),
.A2(n_443),
.B1(n_421),
.B2(n_416),
.C(n_380),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_692),
.B(n_259),
.Y(n_858)
);

O2A1O1Ixp5_ASAP7_75t_L g859 ( 
.A1(n_691),
.A2(n_260),
.B(n_305),
.C(n_257),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_695),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_808),
.B(n_274),
.C(n_266),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_775),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_782),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_683),
.B(n_247),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_714),
.B(n_685),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_749),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_716),
.A2(n_407),
.B1(n_412),
.B2(n_405),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_741),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_809),
.B(n_278),
.C(n_275),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_755),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_684),
.B(n_660),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_747),
.A2(n_480),
.B(n_305),
.C(n_406),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_782),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_790),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_751),
.B(n_364),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_674),
.B(n_364),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_757),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_682),
.B(n_279),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_731),
.B(n_660),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_674),
.B(n_677),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_731),
.B(n_663),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_737),
.B(n_417),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_799),
.B(n_663),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_751),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_828),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_757),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_743),
.A2(n_424),
.B1(n_440),
.B2(n_436),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_772),
.Y(n_888)
);

AND2x6_ASAP7_75t_SL g889 ( 
.A(n_817),
.B(n_308),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_731),
.B(n_665),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_731),
.B(n_665),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_719),
.B(n_721),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_715),
.B(n_667),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_721),
.B(n_296),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_745),
.B(n_667),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_821),
.B(n_668),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_SL g897 ( 
.A1(n_709),
.A2(n_273),
.B1(n_241),
.B2(n_355),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_745),
.A2(n_321),
.B1(n_306),
.B2(n_315),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_832),
.A2(n_408),
.B(n_316),
.C(n_325),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_772),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_724),
.B(n_297),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_790),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_717),
.B(n_668),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_717),
.B(n_669),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_724),
.B(n_299),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_814),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_677),
.B(n_669),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_828),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_677),
.A2(n_321),
.B1(n_306),
.B2(n_315),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_748),
.B(n_671),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_760),
.A2(n_774),
.B(n_690),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_789),
.Y(n_912)
);

NOR2x1p5_ASAP7_75t_L g913 ( 
.A(n_761),
.B(n_304),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_768),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_789),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_694),
.B(n_671),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_700),
.B(n_307),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_767),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_701),
.B(n_426),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_706),
.B(n_240),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_814),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_776),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_798),
.B(n_314),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_787),
.B(n_670),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_703),
.B(n_364),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_807),
.B(n_670),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_738),
.A2(n_406),
.B1(n_327),
.B2(n_329),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_703),
.B(n_364),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_797),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_767),
.Y(n_930)
);

A2O1A1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_774),
.A2(n_680),
.B(n_733),
.C(n_723),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_768),
.Y(n_932)
);

AO22x1_ASAP7_75t_L g933 ( 
.A1(n_822),
.A2(n_326),
.B1(n_330),
.B2(n_332),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_735),
.A2(n_327),
.B(n_425),
.C(n_439),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_797),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_742),
.A2(n_744),
.B(n_818),
.C(n_815),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_805),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_743),
.B(n_329),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_805),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_743),
.B(n_309),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_776),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_R g942 ( 
.A(n_741),
.B(n_621),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_778),
.B(n_670),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_832),
.A2(n_427),
.B(n_368),
.C(n_408),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_743),
.B(n_319),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_778),
.B(n_331),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_703),
.B(n_364),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_819),
.B(n_331),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_819),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_762),
.Y(n_950)
);

NOR2x1p5_ASAP7_75t_L g951 ( 
.A(n_761),
.B(n_328),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_826),
.B(n_339),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_796),
.B(n_337),
.C(n_333),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_709),
.A2(n_454),
.B1(n_438),
.B2(n_446),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_703),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_825),
.B(n_339),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_759),
.B(n_370),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_767),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_703),
.B(n_435),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_678),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_741),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_678),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_765),
.B(n_448),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_689),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_788),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_689),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_770),
.B(n_370),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_702),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_788),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_687),
.B(n_699),
.Y(n_970)
);

BUFx6f_ASAP7_75t_SL g971 ( 
.A(n_754),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_L g972 ( 
.A(n_771),
.B(n_449),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_687),
.B(n_699),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_705),
.B(n_707),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_765),
.B(n_452),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_705),
.B(n_402),
.Y(n_976)
);

AND2x2_ASAP7_75t_SL g977 ( 
.A(n_781),
.B(n_402),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_709),
.A2(n_711),
.B(n_688),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_702),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_707),
.B(n_414),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_752),
.B(n_414),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_765),
.B(n_415),
.Y(n_982)
);

NAND3xp33_ASAP7_75t_L g983 ( 
.A(n_734),
.B(n_348),
.C(n_346),
.Y(n_983)
);

AND2x6_ASAP7_75t_SL g984 ( 
.A(n_788),
.B(n_325),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_771),
.A2(n_415),
.B1(n_425),
.B2(n_439),
.Y(n_985)
);

AND2x2_ASAP7_75t_SL g986 ( 
.A(n_781),
.B(n_326),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_752),
.B(n_505),
.Y(n_987)
);

NOR2x1p5_ASAP7_75t_L g988 ( 
.A(n_823),
.B(n_349),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_L g989 ( 
.A(n_829),
.B(n_801),
.C(n_791),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_710),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_709),
.B(n_350),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_688),
.B(n_330),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_710),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_711),
.A2(n_688),
.B1(n_773),
.B2(n_756),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_754),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_711),
.B(n_353),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_764),
.B(n_769),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_713),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_713),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_765),
.B(n_505),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_754),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_771),
.A2(n_827),
.B1(n_764),
.B2(n_769),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_762),
.B(n_357),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_725),
.Y(n_1004)
);

INVx8_ASAP7_75t_L g1005 ( 
.A(n_971),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_865),
.B(n_830),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_842),
.A2(n_824),
.B(n_795),
.C(n_739),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_837),
.A2(n_880),
.B(n_1000),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_865),
.B(n_830),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_892),
.B(n_830),
.Y(n_1010)
);

AO21x1_ASAP7_75t_L g1011 ( 
.A1(n_842),
.A2(n_802),
.B(n_746),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_R g1012 ( 
.A(n_961),
.B(n_798),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_843),
.A2(n_728),
.B(n_739),
.C(n_688),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_922),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_892),
.B(n_777),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_880),
.A2(n_765),
.B(n_736),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_871),
.B(n_728),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_1000),
.A2(n_736),
.B(n_718),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_853),
.B(n_753),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_853),
.B(n_704),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_851),
.B(n_777),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_858),
.B(n_704),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_844),
.A2(n_736),
.B(n_718),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_848),
.A2(n_740),
.B(n_718),
.Y(n_1024)
);

AO32x1_ASAP7_75t_L g1025 ( 
.A1(n_850),
.A2(n_432),
.A3(n_332),
.B1(n_340),
.B2(n_437),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_866),
.B(n_777),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_SL g1027 ( 
.A1(n_897),
.A2(n_639),
.B1(n_409),
.B2(n_401),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_920),
.B(n_762),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_941),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_982),
.A2(n_771),
.B(n_726),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_856),
.B(n_762),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_849),
.A2(n_810),
.B(n_740),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_852),
.A2(n_810),
.B(n_740),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_858),
.B(n_704),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_917),
.B(n_758),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_885),
.B(n_908),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_846),
.B(n_793),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_847),
.A2(n_812),
.B1(n_820),
.B2(n_686),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_949),
.B(n_758),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_854),
.A2(n_816),
.B(n_810),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_870),
.B(n_730),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_982),
.A2(n_771),
.B(n_726),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_L g1043 ( 
.A(n_918),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_955),
.A2(n_816),
.B(n_780),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_955),
.A2(n_816),
.B(n_780),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1003),
.B(n_800),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_883),
.B(n_806),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_950),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_955),
.A2(n_780),
.B(n_681),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_1001),
.B(n_806),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_960),
.Y(n_1051)
);

AO22x1_ASAP7_75t_L g1052 ( 
.A1(n_989),
.A2(n_794),
.B1(n_779),
.B2(n_792),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_896),
.B(n_758),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_955),
.A2(n_780),
.B(n_681),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_907),
.A2(n_780),
.B(n_681),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_843),
.A2(n_727),
.B(n_725),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_855),
.B(n_783),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_875),
.A2(n_681),
.B(n_766),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_878),
.A2(n_693),
.B1(n_708),
.B2(n_697),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_994),
.B(n_806),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_879),
.A2(n_681),
.B(n_766),
.Y(n_1061)
);

OA22x2_ASAP7_75t_L g1062 ( 
.A1(n_978),
.A2(n_720),
.B1(n_788),
.B2(n_698),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_925),
.A2(n_727),
.B(n_783),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_838),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_857),
.B(n_763),
.C(n_720),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_932),
.Y(n_1066)
);

AO21x1_ASAP7_75t_L g1067 ( 
.A1(n_959),
.A2(n_347),
.B(n_340),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_903),
.B(n_783),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_878),
.B(n_813),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_904),
.B(n_784),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_971),
.B(n_720),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_864),
.A2(n_804),
.B(n_427),
.C(n_432),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_881),
.A2(n_766),
.B(n_811),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_890),
.A2(n_766),
.B(n_811),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_891),
.A2(n_766),
.B(n_811),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_877),
.B(n_784),
.Y(n_1076)
);

AO21x1_ASAP7_75t_L g1077 ( 
.A1(n_959),
.A2(n_347),
.B(n_368),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_886),
.B(n_784),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_888),
.B(n_786),
.Y(n_1079)
);

AOI21x1_ASAP7_75t_L g1080 ( 
.A1(n_925),
.A2(n_514),
.B(n_720),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_864),
.A2(n_437),
.B(n_441),
.C(n_444),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_961),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_L g1083 ( 
.A(n_861),
.B(n_831),
.C(n_413),
.Y(n_1083)
);

OR2x6_ASAP7_75t_SL g1084 ( 
.A(n_953),
.B(n_358),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_893),
.A2(n_910),
.B(n_895),
.Y(n_1085)
);

NOR2x1p5_ASAP7_75t_SL g1086 ( 
.A(n_834),
.B(n_514),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_900),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_833),
.B(n_732),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_911),
.A2(n_803),
.B(n_786),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_963),
.A2(n_803),
.B(n_786),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_977),
.A2(n_986),
.B1(n_915),
.B2(n_929),
.Y(n_1091)
);

INVxp67_ASAP7_75t_L g1092 ( 
.A(n_894),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_894),
.B(n_901),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_872),
.A2(n_975),
.B(n_963),
.C(n_935),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_975),
.A2(n_803),
.B(n_514),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_912),
.B(n_827),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_937),
.B(n_827),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_932),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_916),
.A2(n_947),
.B(n_928),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_962),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_928),
.A2(n_557),
.B(n_555),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_901),
.B(n_361),
.Y(n_1102)
);

INVx4_ASAP7_75t_L g1103 ( 
.A(n_835),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_939),
.B(n_827),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_986),
.A2(n_977),
.B1(n_836),
.B2(n_845),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_905),
.B(n_827),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_947),
.A2(n_785),
.B(n_732),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_914),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_905),
.B(n_365),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_876),
.A2(n_559),
.B(n_557),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_869),
.B(n_419),
.C(n_374),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_914),
.B(n_827),
.Y(n_1112)
);

AO21x1_ASAP7_75t_L g1113 ( 
.A1(n_839),
.A2(n_453),
.B(n_410),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_940),
.A2(n_410),
.B(n_441),
.C(n_444),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_876),
.A2(n_785),
.B(n_732),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_942),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_970),
.A2(n_573),
.B(n_570),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_862),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_919),
.B(n_367),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_956),
.B(n_732),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_839),
.A2(n_785),
.B(n_570),
.Y(n_1121)
);

AOI21x1_ASAP7_75t_L g1122 ( 
.A1(n_943),
.A2(n_565),
.B(n_559),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_995),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_862),
.Y(n_1124)
);

CKINVDCx10_ASAP7_75t_R g1125 ( 
.A(n_942),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_833),
.B(n_369),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_995),
.B(n_240),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_931),
.A2(n_453),
.B(n_411),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_863),
.B(n_785),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_940),
.B(n_240),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_936),
.A2(n_396),
.B(n_447),
.Y(n_1131)
);

NAND2xp33_ASAP7_75t_SL g1132 ( 
.A(n_988),
.B(n_373),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_868),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_973),
.A2(n_565),
.B(n_445),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_974),
.A2(n_431),
.B(n_422),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_938),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_997),
.A2(n_420),
.B(n_375),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_835),
.A2(n_378),
.B(n_398),
.Y(n_1138)
);

AND2x2_ASAP7_75t_SL g1139 ( 
.A(n_938),
.B(n_399),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_835),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_835),
.A2(n_395),
.B(n_391),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_863),
.B(n_873),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_964),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_840),
.A2(n_884),
.B(n_1002),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_873),
.B(n_874),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_945),
.B(n_240),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_945),
.B(n_384),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_840),
.A2(n_388),
.B(n_218),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_840),
.A2(n_213),
.B(n_206),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_991),
.B(n_6),
.Y(n_1150)
);

NOR2x1_ASAP7_75t_L g1151 ( 
.A(n_913),
.B(n_951),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_874),
.B(n_8),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_991),
.B(n_8),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_840),
.A2(n_202),
.B(n_196),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_884),
.B(n_90),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_884),
.A2(n_924),
.B(n_926),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_972),
.A2(n_187),
.B(n_186),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_902),
.B(n_9),
.Y(n_1158)
);

OAI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_996),
.A2(n_10),
.B(n_13),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_841),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_902),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_987),
.A2(n_906),
.B(n_921),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_860),
.B(n_996),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_860),
.B(n_91),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_906),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_921),
.B(n_10),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_983),
.B(n_13),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_930),
.B(n_15),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_964),
.A2(n_185),
.B(n_178),
.Y(n_1169)
);

AND2x2_ASAP7_75t_SL g1170 ( 
.A(n_938),
.B(n_132),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_958),
.B(n_15),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_966),
.A2(n_173),
.B(n_167),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_966),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_968),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_979),
.A2(n_162),
.B(n_161),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_965),
.B(n_16),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_990),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_979),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_887),
.B(n_157),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_998),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_998),
.A2(n_150),
.B(n_149),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_993),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_946),
.B(n_20),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_882),
.A2(n_147),
.B1(n_144),
.B2(n_120),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_899),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_969),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_957),
.A2(n_114),
.B(n_112),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_999),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_944),
.A2(n_867),
.B(n_927),
.C(n_967),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1004),
.A2(n_110),
.B(n_109),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_948),
.A2(n_23),
.B(n_25),
.C(n_27),
.Y(n_1191)
);

AOI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_1093),
.A2(n_954),
.B(n_923),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1136),
.B(n_923),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1093),
.B(n_992),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1016),
.A2(n_980),
.B(n_976),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1029),
.Y(n_1196)
);

AND2x6_ASAP7_75t_SL g1197 ( 
.A(n_1150),
.B(n_923),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1006),
.B(n_1009),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1092),
.B(n_992),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1102),
.A2(n_992),
.B1(n_952),
.B2(n_898),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1092),
.B(n_933),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1036),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1010),
.B(n_909),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1102),
.A2(n_859),
.B(n_934),
.C(n_985),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1140),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1019),
.B(n_889),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1085),
.A2(n_981),
.B(n_834),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1186),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1109),
.A2(n_834),
.B(n_984),
.C(n_30),
.Y(n_1209)
);

BUFx4f_ASAP7_75t_L g1210 ( 
.A(n_1005),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1109),
.B(n_834),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1067),
.A2(n_834),
.A3(n_28),
.B(n_32),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1099),
.A2(n_834),
.B(n_107),
.Y(n_1213)
);

OA21x2_ASAP7_75t_L g1214 ( 
.A1(n_1117),
.A2(n_98),
.B(n_94),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1017),
.B(n_27),
.Y(n_1215)
);

O2A1O1Ixp5_ASAP7_75t_L g1216 ( 
.A1(n_1077),
.A2(n_28),
.B(n_34),
.C(n_36),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1162),
.A2(n_1090),
.B(n_1156),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1118),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1091),
.B(n_36),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1028),
.B(n_1031),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1022),
.A2(n_38),
.B(n_41),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1091),
.B(n_38),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1063),
.A2(n_45),
.B(n_49),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1153),
.A2(n_45),
.B(n_49),
.C(n_50),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1147),
.B(n_50),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1073),
.A2(n_52),
.B(n_54),
.Y(n_1226)
);

BUFx4_ASAP7_75t_SL g1227 ( 
.A(n_1160),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1034),
.A2(n_54),
.B(n_55),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1140),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1037),
.B(n_59),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1011),
.A2(n_61),
.A3(n_62),
.B(n_64),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1037),
.B(n_62),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1065),
.B(n_65),
.Y(n_1233)
);

OAI22x1_ASAP7_75t_L g1234 ( 
.A1(n_1059),
.A2(n_1163),
.B1(n_1041),
.B2(n_1060),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1189),
.A2(n_70),
.B(n_74),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1087),
.B(n_78),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1087),
.B(n_79),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1118),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1005),
.B(n_80),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1094),
.A2(n_81),
.B(n_83),
.C(n_84),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1020),
.B(n_83),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1035),
.A2(n_85),
.B(n_86),
.Y(n_1242)
);

O2A1O1Ixp5_ASAP7_75t_L g1243 ( 
.A1(n_1106),
.A2(n_85),
.B(n_87),
.C(n_1056),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1041),
.B(n_1163),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_1140),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1046),
.Y(n_1246)
);

BUFx10_ASAP7_75t_L g1247 ( 
.A(n_1126),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1074),
.A2(n_1075),
.B(n_1089),
.Y(n_1248)
);

O2A1O1Ixp5_ASAP7_75t_L g1249 ( 
.A1(n_1183),
.A2(n_1105),
.B(n_1113),
.C(n_1166),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1114),
.A2(n_1158),
.A3(n_1152),
.B(n_1008),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1018),
.A2(n_1095),
.B(n_1101),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1144),
.A2(n_1013),
.B(n_1094),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1186),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1119),
.B(n_1130),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1014),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1023),
.A2(n_1033),
.B(n_1040),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1007),
.A2(n_1013),
.B(n_1096),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1119),
.B(n_1146),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1024),
.A2(n_1032),
.B(n_1080),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1069),
.B(n_1015),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1136),
.B(n_1048),
.Y(n_1261)
);

NAND2x1p5_ASAP7_75t_L g1262 ( 
.A(n_1103),
.B(n_1140),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1167),
.A2(n_1038),
.B(n_1159),
.C(n_1139),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1068),
.A2(n_1070),
.B(n_1057),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1064),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1127),
.B(n_1126),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1088),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1007),
.A2(n_1097),
.B(n_1104),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1182),
.B(n_1108),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1030),
.A2(n_1042),
.B(n_1145),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1139),
.A2(n_1062),
.B1(n_1167),
.B2(n_1170),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1044),
.A2(n_1045),
.B(n_1142),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1110),
.A2(n_1061),
.B(n_1039),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1088),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1058),
.A2(n_1112),
.B(n_1129),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1120),
.A2(n_1053),
.B(n_1179),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1076),
.A2(n_1078),
.B(n_1079),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1182),
.B(n_1108),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1164),
.B(n_1066),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_1048),
.Y(n_1280)
);

BUFx4f_ASAP7_75t_L g1281 ( 
.A(n_1005),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1164),
.B(n_1066),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_SL g1283 ( 
.A(n_1131),
.B(n_1128),
.C(n_1050),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1098),
.B(n_1174),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1168),
.A2(n_1072),
.B(n_1111),
.C(n_1137),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_1168),
.A3(n_1161),
.B(n_1165),
.Y(n_1286)
);

AOI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1062),
.A2(n_1047),
.B(n_1176),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1170),
.A2(n_1184),
.B1(n_1177),
.B2(n_1180),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1124),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1051),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1103),
.B(n_1098),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1124),
.A2(n_1054),
.B(n_1049),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1115),
.A2(n_1107),
.B(n_1143),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1176),
.B(n_1123),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1151),
.A2(n_1132),
.B1(n_1052),
.B2(n_1026),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1100),
.B(n_1188),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1173),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1188),
.B(n_1134),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1122),
.A2(n_1055),
.B(n_1155),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1188),
.B(n_1135),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1121),
.A2(n_1081),
.B(n_1072),
.Y(n_1301)
);

AOI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1169),
.A2(n_1175),
.B(n_1181),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_SL g1303 ( 
.A1(n_1185),
.A2(n_1190),
.B(n_1148),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1172),
.A2(n_1154),
.B(n_1149),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1187),
.A2(n_1081),
.B(n_1141),
.Y(n_1305)
);

NAND2xp33_ASAP7_75t_SL g1306 ( 
.A(n_1116),
.B(n_1021),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1188),
.B(n_1178),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1138),
.A2(n_1171),
.B(n_1086),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1185),
.A2(n_1191),
.B(n_1083),
.C(n_1071),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1043),
.B(n_1082),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1043),
.A2(n_1191),
.B(n_1178),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1173),
.A2(n_1178),
.B(n_1084),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1178),
.B(n_1173),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1173),
.A2(n_1025),
.B(n_1133),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1027),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1012),
.A2(n_1093),
.B1(n_1006),
.B2(n_1009),
.Y(n_1316)
);

NOR2x1_ASAP7_75t_L g1317 ( 
.A(n_1125),
.B(n_1025),
.Y(n_1317)
);

NAND2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1103),
.B(n_1140),
.Y(n_1318)
);

AOI21x1_ASAP7_75t_SL g1319 ( 
.A1(n_1106),
.A2(n_1183),
.B(n_1097),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1186),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1093),
.B(n_892),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1099),
.A2(n_843),
.B(n_842),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1103),
.B(n_1140),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1085),
.A2(n_955),
.B(n_1099),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1102),
.C(n_917),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_L g1326 ( 
.A(n_1093),
.B(n_1109),
.C(n_1102),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1029),
.Y(n_1327)
);

AO21x1_ASAP7_75t_L g1328 ( 
.A1(n_1093),
.A2(n_1153),
.B(n_1150),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1117),
.A2(n_1056),
.B(n_1089),
.Y(n_1329)
);

NAND3xp33_ASAP7_75t_L g1330 ( 
.A(n_1093),
.B(n_1109),
.C(n_1102),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1102),
.C(n_917),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1085),
.A2(n_955),
.B(n_1099),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1016),
.A2(n_1162),
.B(n_1090),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1093),
.B(n_892),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1016),
.A2(n_1162),
.B(n_1090),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1016),
.A2(n_1162),
.B(n_1090),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1016),
.A2(n_1162),
.B(n_1090),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1099),
.A2(n_843),
.B(n_842),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1103),
.B(n_1140),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1092),
.B(n_892),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1092),
.B(n_892),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1016),
.A2(n_1162),
.B(n_1090),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1093),
.B(n_1092),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1116),
.Y(n_1344)
);

CKINVDCx8_ASAP7_75t_R g1345 ( 
.A(n_1125),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1016),
.A2(n_1162),
.B(n_1090),
.Y(n_1346)
);

OA22x2_ASAP7_75t_L g1347 ( 
.A1(n_1059),
.A2(n_897),
.B1(n_1027),
.B2(n_1159),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1093),
.B(n_892),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1093),
.A2(n_1109),
.B(n_1102),
.C(n_917),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1092),
.B(n_892),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_SL g1351 ( 
.A1(n_1106),
.A2(n_1183),
.B(n_1097),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1103),
.B(n_1140),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1325),
.A2(n_1331),
.B(n_1349),
.C(n_1326),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1265),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_SL g1355 ( 
.A1(n_1235),
.A2(n_1233),
.B(n_1206),
.C(n_1343),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1196),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1246),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1340),
.B(n_1341),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1227),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1330),
.A2(n_1263),
.B(n_1321),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_L g1361 ( 
.A1(n_1328),
.A2(n_1243),
.B(n_1225),
.C(n_1252),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1334),
.B(n_1348),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1343),
.B(n_1350),
.Y(n_1363)
);

BUFx10_ASAP7_75t_L g1364 ( 
.A(n_1260),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_L g1365 ( 
.A(n_1297),
.B(n_1274),
.Y(n_1365)
);

AO21x1_ASAP7_75t_L g1366 ( 
.A1(n_1198),
.A2(n_1233),
.B(n_1232),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1193),
.B(n_1220),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1266),
.B(n_1206),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1267),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1252),
.A2(n_1257),
.B(n_1322),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_1253),
.Y(n_1371)
);

BUFx8_ASAP7_75t_L g1372 ( 
.A(n_1294),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1347),
.A2(n_1283),
.B1(n_1192),
.B2(n_1271),
.Y(n_1373)
);

AND2x6_ASAP7_75t_L g1374 ( 
.A(n_1297),
.B(n_1317),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1227),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1244),
.B(n_1194),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1254),
.B(n_1258),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1234),
.B(n_1316),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1203),
.B(n_1327),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1247),
.B(n_1202),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1267),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1290),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1253),
.Y(n_1383)
);

AND2x4_ASAP7_75t_SL g1384 ( 
.A(n_1274),
.B(n_1267),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1224),
.A2(n_1230),
.B(n_1240),
.C(n_1283),
.Y(n_1385)
);

CKINVDCx8_ASAP7_75t_R g1386 ( 
.A(n_1197),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1344),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1324),
.A2(n_1332),
.B(n_1211),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1255),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1218),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1202),
.B(n_1199),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1208),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1215),
.B(n_1200),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1288),
.A2(n_1282),
.B1(n_1279),
.B2(n_1284),
.Y(n_1394)
);

BUFx8_ASAP7_75t_L g1395 ( 
.A(n_1315),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1280),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1274),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1238),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1307),
.B(n_1260),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1347),
.B(n_1193),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1320),
.Y(n_1401)
);

INVx3_ASAP7_75t_SL g1402 ( 
.A(n_1239),
.Y(n_1402)
);

BUFx2_ASAP7_75t_SL g1403 ( 
.A(n_1345),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1209),
.A2(n_1201),
.B(n_1222),
.C(n_1219),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1306),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1210),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1296),
.B(n_1288),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1289),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1247),
.B(n_1261),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1269),
.B(n_1278),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1274),
.Y(n_1411)
);

AND2x2_ASAP7_75t_SL g1412 ( 
.A(n_1210),
.B(n_1281),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1338),
.A2(n_1245),
.B1(n_1261),
.B2(n_1295),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1297),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1249),
.A2(n_1285),
.B(n_1241),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1291),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1280),
.B(n_1236),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1310),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1313),
.B(n_1277),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1245),
.A2(n_1291),
.B1(n_1324),
.B2(n_1332),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1237),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1297),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1262),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1287),
.B(n_1312),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1281),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1205),
.B(n_1229),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1314),
.A2(n_1303),
.B1(n_1311),
.B2(n_1300),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1298),
.B(n_1268),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1352),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1207),
.A2(n_1276),
.B(n_1213),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1205),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1239),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1207),
.A2(n_1276),
.B(n_1213),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1229),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1270),
.B(n_1309),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1249),
.A2(n_1204),
.B(n_1301),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1262),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1239),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1256),
.A2(n_1217),
.B(n_1346),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1318),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1242),
.B(n_1228),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1308),
.B(n_1352),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1318),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1293),
.B(n_1304),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1309),
.B(n_1221),
.C(n_1228),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1292),
.B(n_1275),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1221),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1323),
.B(n_1339),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1333),
.A2(n_1335),
.B(n_1342),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1339),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1319),
.Y(n_1451)
);

AND2x2_ASAP7_75t_SL g1452 ( 
.A(n_1270),
.B(n_1329),
.Y(n_1452)
);

BUFx2_ASAP7_75t_SL g1453 ( 
.A(n_1214),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1223),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1243),
.A2(n_1305),
.B(n_1264),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1226),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1299),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1351),
.Y(n_1458)
);

INVx3_ASAP7_75t_SL g1459 ( 
.A(n_1214),
.Y(n_1459)
);

INVx3_ASAP7_75t_SL g1460 ( 
.A(n_1329),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1231),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1216),
.A2(n_1248),
.B(n_1195),
.C(n_1337),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_SL g1463 ( 
.A(n_1302),
.B(n_1250),
.Y(n_1463)
);

O2A1O1Ixp5_ASAP7_75t_SL g1464 ( 
.A1(n_1231),
.A2(n_1216),
.B(n_1212),
.C(n_1286),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1273),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1272),
.B(n_1336),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1231),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1231),
.B(n_1212),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1212),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1212),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1251),
.B(n_1259),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1246),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1193),
.B(n_1220),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1344),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1245),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1321),
.B(n_1334),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1326),
.A2(n_1330),
.B1(n_1331),
.B2(n_1325),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1246),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1325),
.A2(n_1349),
.B(n_1331),
.C(n_1093),
.Y(n_1479)
);

NAND2xp33_ASAP7_75t_L g1480 ( 
.A(n_1325),
.B(n_1331),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1246),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1326),
.A2(n_1330),
.B1(n_1331),
.B2(n_1325),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1274),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1246),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_SL g1485 ( 
.A1(n_1235),
.A2(n_1093),
.B(n_1153),
.C(n_1150),
.Y(n_1485)
);

INVx5_ASAP7_75t_L g1486 ( 
.A(n_1274),
.Y(n_1486)
);

NOR2xp67_ASAP7_75t_SL g1487 ( 
.A(n_1345),
.B(n_961),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1246),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1340),
.B(n_1341),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1253),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1321),
.B(n_1334),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1325),
.A2(n_1349),
.B(n_1331),
.Y(n_1492)
);

BUFx4f_ASAP7_75t_SL g1493 ( 
.A(n_1246),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1325),
.A2(n_1349),
.B(n_1331),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1267),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1344),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1325),
.A2(n_1349),
.B(n_1331),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1246),
.B(n_800),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1344),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1326),
.A2(n_1093),
.B1(n_1330),
.B2(n_1109),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1321),
.B(n_1334),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1325),
.A2(n_1349),
.B(n_1331),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1246),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1265),
.Y(n_1504)
);

BUFx12f_ASAP7_75t_L g1505 ( 
.A(n_1344),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1325),
.A2(n_1331),
.B(n_1349),
.C(n_1263),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1267),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1340),
.B(n_1341),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1246),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1321),
.B(n_1334),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1274),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1326),
.B(n_1330),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1265),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1325),
.A2(n_1349),
.B(n_1331),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1196),
.Y(n_1515)
);

OR2x6_ASAP7_75t_L g1516 ( 
.A(n_1279),
.B(n_1005),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1253),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1325),
.A2(n_1349),
.B(n_1331),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1265),
.Y(n_1519)
);

NAND2x1_ASAP7_75t_L g1520 ( 
.A(n_1297),
.B(n_1103),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1274),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1340),
.B(n_1341),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1321),
.B(n_1334),
.Y(n_1523)
);

BUFx12f_ASAP7_75t_L g1524 ( 
.A(n_1344),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1279),
.B(n_1005),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1253),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1227),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1469),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1377),
.B(n_1362),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1428),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1360),
.B(n_1377),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1428),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1480),
.A2(n_1514),
.B1(n_1373),
.B2(n_1482),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1479),
.A2(n_1506),
.B(n_1353),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1439),
.A2(n_1449),
.B(n_1433),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1515),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1354),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1477),
.A2(n_1494),
.B1(n_1497),
.B2(n_1492),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1488),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1504),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1505),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1513),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1519),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1382),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1389),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1472),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1500),
.A2(n_1362),
.B1(n_1491),
.B2(n_1523),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1405),
.A2(n_1368),
.B1(n_1367),
.B2(n_1473),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1442),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1441),
.Y(n_1550)
);

BUFx12f_ASAP7_75t_L g1551 ( 
.A(n_1524),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1435),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1475),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1357),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_SL g1555 ( 
.A(n_1395),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1512),
.A2(n_1492),
.B1(n_1494),
.B2(n_1497),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1485),
.A2(n_1518),
.B(n_1506),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1430),
.A2(n_1433),
.B(n_1388),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1478),
.Y(n_1559)
);

OA21x2_ASAP7_75t_L g1560 ( 
.A1(n_1455),
.A2(n_1436),
.B(n_1415),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1486),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1435),
.Y(n_1562)
);

BUFx4f_ASAP7_75t_SL g1563 ( 
.A(n_1496),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1467),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1361),
.A2(n_1430),
.B(n_1462),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1518),
.A2(n_1447),
.B1(n_1366),
.B2(n_1393),
.Y(n_1566)
);

CKINVDCx11_ASAP7_75t_R g1567 ( 
.A(n_1386),
.Y(n_1567)
);

BUFx12f_ASAP7_75t_L g1568 ( 
.A(n_1387),
.Y(n_1568)
);

AO21x1_ASAP7_75t_SL g1569 ( 
.A1(n_1393),
.A2(n_1378),
.B(n_1427),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1481),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1370),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1378),
.A2(n_1400),
.B1(n_1445),
.B2(n_1421),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1376),
.A2(n_1491),
.B1(n_1501),
.B2(n_1510),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1468),
.Y(n_1574)
);

BUFx4f_ASAP7_75t_SL g1575 ( 
.A(n_1406),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1408),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1437),
.Y(n_1577)
);

AOI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1420),
.A2(n_1471),
.B(n_1444),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1438),
.A2(n_1364),
.B1(n_1395),
.B2(n_1372),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1364),
.A2(n_1372),
.B1(n_1409),
.B2(n_1412),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1390),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1475),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1412),
.A2(n_1476),
.B1(n_1510),
.B2(n_1523),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1474),
.Y(n_1584)
);

BUFx4f_ASAP7_75t_L g1585 ( 
.A(n_1369),
.Y(n_1585)
);

BUFx2_ASAP7_75t_R g1586 ( 
.A(n_1403),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1398),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1355),
.A2(n_1385),
.B(n_1394),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_SL g1589 ( 
.A(n_1499),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1367),
.A2(n_1473),
.B1(n_1501),
.B2(n_1476),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1376),
.B(n_1399),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1484),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1383),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1363),
.A2(n_1493),
.B1(n_1418),
.B2(n_1498),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_R g1595 ( 
.A1(n_1359),
.A2(n_1527),
.B1(n_1375),
.B2(n_1396),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1493),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1385),
.A2(n_1361),
.B(n_1404),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1363),
.A2(n_1399),
.B1(n_1503),
.B2(n_1509),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1396),
.Y(n_1599)
);

BUFx4_ASAP7_75t_SL g1600 ( 
.A(n_1425),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1413),
.A2(n_1374),
.B1(n_1470),
.B2(n_1522),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1383),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1490),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1374),
.A2(n_1358),
.B1(n_1489),
.B2(n_1508),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1374),
.A2(n_1391),
.B1(n_1417),
.B2(n_1407),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1374),
.A2(n_1379),
.B1(n_1407),
.B2(n_1458),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1374),
.A2(n_1380),
.B1(n_1379),
.B2(n_1424),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1490),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1517),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1410),
.B(n_1419),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1402),
.A2(n_1432),
.B1(n_1525),
.B2(n_1516),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1404),
.A2(n_1419),
.B(n_1410),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1392),
.Y(n_1613)
);

BUFx4_ASAP7_75t_R g1614 ( 
.A(n_1429),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1517),
.B(n_1526),
.Y(n_1615)
);

AOI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1471),
.A2(n_1444),
.B(n_1446),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1402),
.A2(n_1525),
.B1(n_1516),
.B2(n_1401),
.Y(n_1617)
);

AOI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1446),
.A2(n_1466),
.B(n_1465),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_SL g1619 ( 
.A1(n_1526),
.A2(n_1525),
.B1(n_1516),
.B2(n_1461),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1371),
.Y(n_1620)
);

AO21x1_ASAP7_75t_SL g1621 ( 
.A1(n_1464),
.A2(n_1431),
.B(n_1434),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1416),
.B(n_1422),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1457),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1454),
.A2(n_1520),
.B(n_1414),
.Y(n_1624)
);

OAI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1456),
.A2(n_1451),
.B(n_1448),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1371),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1443),
.A2(n_1423),
.B1(n_1450),
.B2(n_1437),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1426),
.Y(n_1628)
);

AO21x2_ASAP7_75t_L g1629 ( 
.A1(n_1463),
.A2(n_1456),
.B(n_1466),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1369),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_SL g1631 ( 
.A(n_1451),
.B(n_1453),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1414),
.Y(n_1632)
);

OAI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1486),
.A2(n_1521),
.B1(n_1450),
.B2(n_1440),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1422),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1486),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1457),
.Y(n_1636)
);

INVx4_ASAP7_75t_L g1637 ( 
.A(n_1521),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1426),
.B(n_1423),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1451),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1451),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1452),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1452),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1460),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1365),
.A2(n_1511),
.B(n_1483),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1521),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1365),
.A2(n_1511),
.B(n_1483),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1440),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1440),
.Y(n_1648)
);

INVxp33_ASAP7_75t_L g1649 ( 
.A(n_1487),
.Y(n_1649)
);

AOI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1459),
.A2(n_1460),
.B(n_1450),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1411),
.A2(n_1397),
.B1(n_1381),
.B2(n_1495),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1411),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1397),
.B(n_1521),
.Y(n_1653)
);

BUFx8_ASAP7_75t_L g1654 ( 
.A(n_1381),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1459),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1495),
.A2(n_1330),
.B1(n_1326),
.B2(n_1093),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1507),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_1384),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1507),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1442),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1360),
.B(n_1377),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1356),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1500),
.A2(n_1093),
.B1(n_1330),
.B2(n_1326),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1356),
.Y(n_1664)
);

INVxp67_ASAP7_75t_L g1665 ( 
.A(n_1472),
.Y(n_1665)
);

OR2x6_ASAP7_75t_L g1666 ( 
.A(n_1502),
.B(n_1506),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1442),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1357),
.Y(n_1668)
);

NOR2x1_ASAP7_75t_R g1669 ( 
.A(n_1403),
.B(n_1001),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1403),
.Y(n_1670)
);

AO21x1_ASAP7_75t_L g1671 ( 
.A1(n_1480),
.A2(n_1482),
.B(n_1477),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1357),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1356),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1455),
.A2(n_1436),
.B(n_1415),
.Y(n_1674)
);

CKINVDCx11_ASAP7_75t_R g1675 ( 
.A(n_1496),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1356),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1356),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_SL g1678 ( 
.A1(n_1514),
.A2(n_1093),
.B1(n_1330),
.B2(n_1326),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1377),
.B(n_1321),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1480),
.A2(n_1330),
.B1(n_1326),
.B2(n_1093),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1356),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1500),
.A2(n_1093),
.B1(n_1330),
.B2(n_1326),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1475),
.Y(n_1683)
);

BUFx12f_ASAP7_75t_L g1684 ( 
.A(n_1505),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1480),
.A2(n_1330),
.B1(n_1326),
.B2(n_1093),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1442),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1356),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_SL g1688 ( 
.A1(n_1514),
.A2(n_1093),
.B1(n_1330),
.B2(n_1326),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1475),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1472),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1360),
.B(n_1377),
.Y(n_1691)
);

AO21x2_ASAP7_75t_L g1692 ( 
.A1(n_1597),
.A2(n_1588),
.B(n_1557),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1599),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1550),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1620),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1550),
.Y(n_1696)
);

INVx5_ASAP7_75t_L g1697 ( 
.A(n_1666),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1529),
.B(n_1573),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1658),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1528),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1602),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1591),
.B(n_1547),
.Y(n_1702)
);

NAND2xp33_ASAP7_75t_R g1703 ( 
.A(n_1670),
.B(n_1626),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1615),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1533),
.A2(n_1682),
.B1(n_1663),
.B2(n_1671),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1603),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1593),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1583),
.B(n_1678),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1574),
.B(n_1552),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1608),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1609),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1553),
.Y(n_1712)
);

BUFx3_ASAP7_75t_L g1713 ( 
.A(n_1658),
.Y(n_1713)
);

INVx6_ASAP7_75t_L g1714 ( 
.A(n_1654),
.Y(n_1714)
);

INVx2_ASAP7_75t_SL g1715 ( 
.A(n_1537),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1561),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1553),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1537),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1675),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1582),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1582),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1591),
.B(n_1679),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1589),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1535),
.A2(n_1558),
.B(n_1578),
.Y(n_1724)
);

NAND2x1p5_ASAP7_75t_L g1725 ( 
.A(n_1683),
.B(n_1650),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1683),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1574),
.B(n_1531),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1688),
.B(n_1680),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1552),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1562),
.B(n_1641),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1531),
.B(n_1661),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1562),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1564),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1564),
.Y(n_1734)
);

INVx4_ASAP7_75t_L g1735 ( 
.A(n_1561),
.Y(n_1735)
);

INVx4_ASAP7_75t_L g1736 ( 
.A(n_1561),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1654),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1539),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1616),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1661),
.B(n_1691),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1549),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1671),
.A2(n_1666),
.B1(n_1685),
.B2(n_1538),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1666),
.B(n_1534),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1641),
.B(n_1642),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1691),
.B(n_1610),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1632),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1549),
.B(n_1660),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1654),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1632),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1618),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1626),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1546),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1642),
.B(n_1610),
.Y(n_1753)
);

OA21x2_ASAP7_75t_L g1754 ( 
.A1(n_1612),
.A2(n_1571),
.B(n_1566),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1616),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1549),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1660),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1655),
.Y(n_1758)
);

OAI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1534),
.A2(n_1556),
.B(n_1656),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1660),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1572),
.B(n_1590),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1655),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1548),
.B(n_1614),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1569),
.B(n_1667),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1686),
.B(n_1643),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1559),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1540),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1560),
.B(n_1674),
.Y(n_1768)
);

INVx5_ASAP7_75t_SL g1769 ( 
.A(n_1666),
.Y(n_1769)
);

AO21x2_ASAP7_75t_L g1770 ( 
.A1(n_1625),
.A2(n_1578),
.B(n_1650),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1560),
.B(n_1674),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1570),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1613),
.Y(n_1773)
);

OAI21x1_ASAP7_75t_L g1774 ( 
.A1(n_1624),
.A2(n_1565),
.B(n_1639),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1560),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1560),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1674),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1629),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1569),
.B(n_1530),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1530),
.B(n_1532),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1690),
.Y(n_1782)
);

BUFx3_ASAP7_75t_L g1783 ( 
.A(n_1554),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_R g1784 ( 
.A1(n_1594),
.A2(n_1598),
.B(n_1595),
.Y(n_1784)
);

AO21x2_ASAP7_75t_L g1785 ( 
.A1(n_1631),
.A2(n_1640),
.B(n_1629),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1674),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1689),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1561),
.Y(n_1788)
);

OAI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1649),
.A2(n_1607),
.B(n_1606),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1532),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1565),
.B(n_1601),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1665),
.B(n_1554),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1592),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1592),
.B(n_1668),
.Y(n_1794)
);

OR2x6_ASAP7_75t_L g1795 ( 
.A(n_1565),
.B(n_1639),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1662),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1565),
.B(n_1605),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1664),
.B(n_1673),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1631),
.A2(n_1633),
.B(n_1637),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1604),
.B(n_1617),
.C(n_1611),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1544),
.Y(n_1802)
);

AO21x2_ASAP7_75t_L g1803 ( 
.A1(n_1640),
.A2(n_1636),
.B(n_1576),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_1668),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1681),
.B(n_1687),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1681),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1613),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1731),
.B(n_1621),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1731),
.B(n_1621),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1700),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1746),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1740),
.B(n_1619),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1803),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1797),
.B(n_1536),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_SL g1815 ( 
.A(n_1743),
.B(n_1635),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1697),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1740),
.B(n_1677),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1727),
.B(n_1676),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1727),
.B(n_1545),
.Y(n_1819)
);

INVxp67_ASAP7_75t_SL g1820 ( 
.A(n_1750),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1753),
.B(n_1545),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1749),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1803),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1753),
.B(n_1622),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1779),
.Y(n_1825)
);

OR2x2_ASAP7_75t_SL g1826 ( 
.A(n_1791),
.B(n_1702),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1797),
.B(n_1581),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1765),
.B(n_1622),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1747),
.B(n_1644),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1768),
.B(n_1587),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1768),
.B(n_1771),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1765),
.B(n_1638),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1771),
.B(n_1657),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1765),
.B(n_1638),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1747),
.B(n_1646),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1725),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1765),
.B(n_1652),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1747),
.B(n_1657),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1707),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1747),
.B(n_1634),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1756),
.B(n_1648),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1756),
.B(n_1647),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1757),
.B(n_1646),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1760),
.B(n_1644),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1760),
.B(n_1577),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1705),
.A2(n_1580),
.B1(n_1555),
.B2(n_1579),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1791),
.B(n_1628),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1742),
.A2(n_1586),
.B1(n_1627),
.B2(n_1630),
.Y(n_1848)
);

NOR2xp67_ASAP7_75t_L g1849 ( 
.A(n_1739),
.B(n_1577),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1744),
.B(n_1659),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1697),
.B(n_1653),
.Y(n_1851)
);

HB1xp67_ASAP7_75t_L g1852 ( 
.A(n_1741),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1697),
.B(n_1653),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1785),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1741),
.Y(n_1855)
);

BUFx2_ASAP7_75t_L g1856 ( 
.A(n_1725),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1725),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1785),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1728),
.A2(n_1595),
.B1(n_1551),
.B2(n_1684),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1708),
.A2(n_1541),
.B1(n_1551),
.B2(n_1684),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1712),
.Y(n_1861)
);

NOR2x1_ASAP7_75t_L g1862 ( 
.A(n_1692),
.B(n_1637),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1717),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1779),
.Y(n_1864)
);

OR2x6_ASAP7_75t_L g1865 ( 
.A(n_1743),
.B(n_1561),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1697),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1743),
.A2(n_1541),
.B1(n_1672),
.B2(n_1568),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1692),
.B(n_1672),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1785),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1784),
.A2(n_1630),
.B1(n_1651),
.B2(n_1670),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1743),
.A2(n_1568),
.B1(n_1567),
.B2(n_1563),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1717),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1704),
.B(n_1645),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1692),
.B(n_1596),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1697),
.B(n_1739),
.Y(n_1875)
);

AOI21xp33_ASAP7_75t_L g1876 ( 
.A1(n_1759),
.A2(n_1669),
.B(n_1635),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1839),
.B(n_1695),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1808),
.B(n_1795),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1861),
.B(n_1745),
.Y(n_1879)
);

NAND3xp33_ASAP7_75t_L g1880 ( 
.A(n_1874),
.B(n_1789),
.C(n_1801),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1874),
.B(n_1698),
.Y(n_1881)
);

OAI221xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1860),
.A2(n_1743),
.B1(n_1761),
.B2(n_1763),
.C(n_1738),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1811),
.B(n_1752),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1846),
.A2(n_1848),
.B1(n_1859),
.B2(n_1876),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_L g1885 ( 
.A(n_1868),
.B(n_1780),
.C(n_1800),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1846),
.A2(n_1697),
.B1(n_1769),
.B2(n_1714),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1822),
.B(n_1766),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1848),
.A2(n_1754),
.B1(n_1769),
.B2(n_1772),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1808),
.B(n_1795),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1871),
.A2(n_1769),
.B1(n_1714),
.B2(n_1751),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1809),
.B(n_1795),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1809),
.B(n_1795),
.Y(n_1892)
);

NAND4xp25_ASAP7_75t_L g1893 ( 
.A(n_1868),
.B(n_1722),
.C(n_1792),
.D(n_1773),
.Y(n_1893)
);

NAND3xp33_ASAP7_75t_L g1894 ( 
.A(n_1876),
.B(n_1780),
.C(n_1782),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1832),
.B(n_1834),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1819),
.B(n_1821),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1867),
.A2(n_1870),
.B1(n_1769),
.B2(n_1826),
.Y(n_1897)
);

OAI221xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1847),
.A2(n_1807),
.B1(n_1764),
.B2(n_1795),
.C(n_1799),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1866),
.B(n_1787),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1819),
.B(n_1758),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1821),
.B(n_1762),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1815),
.A2(n_1754),
.B(n_1635),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_L g1903 ( 
.A(n_1862),
.B(n_1764),
.C(n_1762),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1870),
.A2(n_1754),
.B1(n_1699),
.B2(n_1713),
.Y(n_1904)
);

OA211x2_ASAP7_75t_L g1905 ( 
.A1(n_1823),
.A2(n_1794),
.B(n_1781),
.C(n_1805),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1817),
.B(n_1710),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1817),
.B(n_1711),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1847),
.B(n_1730),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1873),
.B(n_1693),
.Y(n_1909)
);

OAI21xp33_ASAP7_75t_L g1910 ( 
.A1(n_1812),
.A2(n_1730),
.B(n_1696),
.Y(n_1910)
);

NAND4xp25_ASAP7_75t_L g1911 ( 
.A(n_1814),
.B(n_1799),
.C(n_1703),
.D(n_1802),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1843),
.B(n_1739),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1828),
.B(n_1787),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1843),
.B(n_1755),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1812),
.A2(n_1802),
.B1(n_1767),
.B2(n_1701),
.C(n_1706),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1832),
.B(n_1699),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1834),
.B(n_1713),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1828),
.B(n_1701),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1838),
.B(n_1706),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1838),
.B(n_1767),
.Y(n_1920)
);

OA21x2_ASAP7_75t_L g1921 ( 
.A1(n_1823),
.A2(n_1724),
.B(n_1774),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1810),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1844),
.B(n_1755),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1856),
.A2(n_1694),
.B1(n_1696),
.B2(n_1775),
.C(n_1790),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1824),
.B(n_1694),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1865),
.A2(n_1829),
.B1(n_1835),
.B2(n_1714),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1824),
.B(n_1790),
.Y(n_1927)
);

OAI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1836),
.A2(n_1719),
.B1(n_1804),
.B2(n_1783),
.C(n_1793),
.Y(n_1928)
);

AOI22xp33_ASAP7_75t_L g1929 ( 
.A1(n_1865),
.A2(n_1754),
.B1(n_1714),
.B2(n_1748),
.Y(n_1929)
);

OAI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1836),
.A2(n_1857),
.B1(n_1856),
.B2(n_1719),
.C(n_1783),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1866),
.B(n_1775),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1840),
.B(n_1720),
.Y(n_1932)
);

NAND4xp25_ASAP7_75t_L g1933 ( 
.A(n_1814),
.B(n_1804),
.C(n_1793),
.D(n_1733),
.Y(n_1933)
);

NOR3xp33_ASAP7_75t_L g1934 ( 
.A(n_1862),
.B(n_1736),
.C(n_1716),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1840),
.B(n_1721),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1818),
.B(n_1726),
.Y(n_1936)
);

OAI21xp5_ASAP7_75t_SL g1937 ( 
.A1(n_1866),
.A2(n_1788),
.B(n_1755),
.Y(n_1937)
);

NAND3xp33_ASAP7_75t_L g1938 ( 
.A(n_1827),
.B(n_1734),
.C(n_1733),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1818),
.B(n_1729),
.Y(n_1939)
);

OA21x2_ASAP7_75t_L g1940 ( 
.A1(n_1854),
.A2(n_1774),
.B(n_1786),
.Y(n_1940)
);

NAND3xp33_ASAP7_75t_L g1941 ( 
.A(n_1827),
.B(n_1734),
.C(n_1796),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1866),
.B(n_1775),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1837),
.B(n_1729),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1837),
.B(n_1732),
.Y(n_1944)
);

NAND3xp33_ASAP7_75t_L g1945 ( 
.A(n_1857),
.B(n_1806),
.C(n_1786),
.Y(n_1945)
);

NAND3xp33_ASAP7_75t_L g1946 ( 
.A(n_1836),
.B(n_1813),
.C(n_1830),
.Y(n_1946)
);

OAI21xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1866),
.A2(n_1788),
.B(n_1732),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1866),
.A2(n_1788),
.B(n_1709),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1829),
.B(n_1770),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1841),
.B(n_1715),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1826),
.A2(n_1748),
.B1(n_1737),
.B2(n_1723),
.Y(n_1951)
);

OAI21xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1851),
.A2(n_1853),
.B(n_1875),
.Y(n_1952)
);

NAND3xp33_ASAP7_75t_L g1953 ( 
.A(n_1813),
.B(n_1778),
.C(n_1777),
.Y(n_1953)
);

XOR2xp5_ASAP7_75t_L g1954 ( 
.A(n_1851),
.B(n_1584),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1841),
.B(n_1715),
.Y(n_1955)
);

OAI21xp5_ASAP7_75t_SL g1956 ( 
.A1(n_1851),
.A2(n_1788),
.B(n_1709),
.Y(n_1956)
);

OAI21xp33_ASAP7_75t_L g1957 ( 
.A1(n_1844),
.A2(n_1778),
.B(n_1776),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1831),
.B(n_1776),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1850),
.B(n_1770),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1842),
.B(n_1718),
.Y(n_1960)
);

NAND3xp33_ASAP7_75t_L g1961 ( 
.A(n_1830),
.B(n_1777),
.C(n_1798),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1940),
.Y(n_1962)
);

BUFx2_ASAP7_75t_L g1963 ( 
.A(n_1878),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1878),
.B(n_1835),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1922),
.Y(n_1965)
);

AND2x2_ASAP7_75t_SL g1966 ( 
.A(n_1888),
.B(n_1816),
.Y(n_1966)
);

AND2x4_ASAP7_75t_SL g1967 ( 
.A(n_1934),
.B(n_1865),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1889),
.B(n_1831),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1958),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1891),
.B(n_1892),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1940),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1949),
.B(n_1875),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1881),
.B(n_1863),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1908),
.B(n_1833),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1940),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1881),
.B(n_1863),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1912),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1958),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1912),
.Y(n_1979)
);

NAND2x1_ASAP7_75t_L g1980 ( 
.A(n_1902),
.B(n_1816),
.Y(n_1980)
);

NAND2x1_ASAP7_75t_L g1981 ( 
.A(n_1903),
.B(n_1816),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1914),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1891),
.B(n_1875),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1914),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1926),
.B(n_1923),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1923),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1931),
.B(n_1816),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1938),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1892),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1961),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1877),
.B(n_1833),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1936),
.B(n_1872),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_1899),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1959),
.B(n_1957),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1953),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1895),
.B(n_1852),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1954),
.B(n_1723),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1899),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1900),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1901),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1952),
.B(n_1855),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1921),
.Y(n_2002)
);

INVx4_ASAP7_75t_L g2003 ( 
.A(n_1921),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1896),
.B(n_1825),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1883),
.B(n_1845),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1959),
.B(n_1820),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1943),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1921),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1944),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1916),
.B(n_1917),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1887),
.B(n_1879),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1956),
.B(n_1929),
.Y(n_2012)
);

NOR2xp67_ASAP7_75t_L g2013 ( 
.A(n_1885),
.B(n_1825),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1925),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1941),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1932),
.B(n_1935),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1909),
.Y(n_2017)
);

BUFx2_ASAP7_75t_L g2018 ( 
.A(n_1946),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1929),
.B(n_1825),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1931),
.B(n_1825),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1950),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1913),
.B(n_1820),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1955),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1942),
.B(n_1864),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1960),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_1920),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_1919),
.Y(n_2027)
);

INVx2_ASAP7_75t_SL g2028 ( 
.A(n_1942),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_1990),
.B(n_1906),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_2015),
.B(n_1880),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1990),
.B(n_1907),
.Y(n_2031)
);

NOR2x1_ASAP7_75t_L g2032 ( 
.A(n_2013),
.B(n_1951),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1972),
.B(n_2001),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1972),
.B(n_1948),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1965),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1995),
.B(n_1927),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1965),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1969),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1972),
.B(n_1937),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1962),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2015),
.B(n_1893),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1966),
.A2(n_1884),
.B1(n_1897),
.B2(n_1886),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1969),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1978),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2023),
.B(n_1918),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_1995),
.B(n_1939),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2023),
.B(n_1915),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1978),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1974),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_1994),
.B(n_1898),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_2023),
.B(n_1910),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_1994),
.B(n_1945),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2023),
.B(n_1894),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1962),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1988),
.B(n_1911),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1962),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1988),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1974),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2013),
.A2(n_1884),
.B1(n_1904),
.B2(n_1882),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1979),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1979),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1972),
.B(n_1947),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1982),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1982),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1997),
.B(n_1928),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2001),
.B(n_1815),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1971),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_1968),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1963),
.B(n_1865),
.Y(n_2069)
);

INVxp67_ASAP7_75t_SL g2070 ( 
.A(n_1981),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1986),
.Y(n_2071)
);

NOR2x1p5_ASAP7_75t_SL g2072 ( 
.A(n_2002),
.B(n_2008),
.Y(n_2072)
);

AND2x4_ASAP7_75t_SL g2073 ( 
.A(n_2010),
.B(n_1865),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1986),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_1980),
.Y(n_2075)
);

NAND2x1_ASAP7_75t_SL g2076 ( 
.A(n_2012),
.B(n_1864),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2022),
.Y(n_2077)
);

NAND2x2_ASAP7_75t_L g2078 ( 
.A(n_1980),
.B(n_1737),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1971),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2022),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2006),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1971),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1967),
.B(n_1849),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1963),
.B(n_1989),
.Y(n_2084)
);

NAND2x2_ASAP7_75t_L g2085 ( 
.A(n_1981),
.B(n_1600),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2030),
.B(n_2041),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2035),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2033),
.B(n_2039),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2042),
.A2(n_1904),
.B1(n_1888),
.B2(n_1966),
.Y(n_2089)
);

NAND4xp25_ASAP7_75t_L g2090 ( 
.A(n_2055),
.B(n_1905),
.C(n_2018),
.D(n_1930),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2033),
.B(n_1964),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2037),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2057),
.B(n_2047),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2039),
.B(n_1989),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_2059),
.A2(n_1966),
.B1(n_2012),
.B2(n_1890),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_2065),
.B(n_2018),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2029),
.B(n_2031),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_2029),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2031),
.B(n_1993),
.Y(n_2099)
);

OR2x6_ASAP7_75t_L g2100 ( 
.A(n_2075),
.B(n_1987),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2058),
.B(n_2050),
.Y(n_2101)
);

INVxp67_ASAP7_75t_L g2102 ( 
.A(n_2046),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_2050),
.B(n_2052),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2074),
.Y(n_2104)
);

NAND2x1p5_ASAP7_75t_L g2105 ( 
.A(n_2075),
.B(n_1993),
.Y(n_2105)
);

NAND2xp33_ASAP7_75t_R g2106 ( 
.A(n_2052),
.B(n_1987),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2049),
.B(n_1992),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2074),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2036),
.B(n_1998),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2038),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2040),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2034),
.B(n_1964),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2034),
.B(n_1985),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2062),
.B(n_1985),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2036),
.B(n_1998),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_2084),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2046),
.B(n_2007),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2038),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2043),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2040),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2054),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2043),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2053),
.B(n_2007),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2077),
.B(n_2009),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2044),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2044),
.Y(n_2126)
);

NAND2x1p5_ASAP7_75t_L g2127 ( 
.A(n_2032),
.B(n_1987),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2062),
.B(n_2084),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2054),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2048),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2048),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_2076),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2060),
.Y(n_2133)
);

AND2x4_ASAP7_75t_SL g2134 ( 
.A(n_2083),
.B(n_1987),
.Y(n_2134)
);

NOR5xp2_ASAP7_75t_SL g2135 ( 
.A(n_2076),
.B(n_1924),
.C(n_1967),
.D(n_2028),
.E(n_1933),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_2051),
.B(n_2011),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2061),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2063),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_2083),
.B(n_2070),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2066),
.B(n_1985),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2077),
.B(n_2009),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2080),
.B(n_2017),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_SL g2143 ( 
.A(n_2096),
.B(n_2083),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2127),
.B(n_2066),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_2101),
.B(n_2080),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_2086),
.B(n_1584),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_2128),
.B(n_2069),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2104),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2108),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2127),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2110),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_2096),
.B(n_2049),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2116),
.Y(n_2153)
);

OAI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2095),
.A2(n_2085),
.B1(n_2078),
.B2(n_1967),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2128),
.B(n_2069),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2103),
.B(n_2068),
.Y(n_2156)
);

NAND3xp33_ASAP7_75t_L g2157 ( 
.A(n_2103),
.B(n_2081),
.C(n_2067),
.Y(n_2157)
);

CKINVDCx16_ASAP7_75t_R g2158 ( 
.A(n_2106),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2087),
.Y(n_2159)
);

NOR2x1_ASAP7_75t_L g2160 ( 
.A(n_2090),
.B(n_2081),
.Y(n_2160)
);

AOI222xp33_ASAP7_75t_L g2161 ( 
.A1(n_2089),
.A2(n_1973),
.B1(n_1976),
.B2(n_2019),
.C1(n_2021),
.C2(n_2025),
.Y(n_2161)
);

AND2x4_ASAP7_75t_L g2162 ( 
.A(n_2088),
.B(n_2139),
.Y(n_2162)
);

NOR2x1_ASAP7_75t_L g2163 ( 
.A(n_2093),
.B(n_2056),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2097),
.B(n_2064),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2136),
.B(n_2028),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2116),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2094),
.Y(n_2167)
);

INVx1_ASAP7_75t_SL g2168 ( 
.A(n_2139),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2092),
.Y(n_2169)
);

INVx3_ASAP7_75t_SL g2170 ( 
.A(n_2100),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2107),
.B(n_2071),
.Y(n_2171)
);

HB1xp67_ASAP7_75t_L g2172 ( 
.A(n_2094),
.Y(n_2172)
);

INVx3_ASAP7_75t_SL g2173 ( 
.A(n_2100),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2118),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2114),
.B(n_2073),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2136),
.B(n_2045),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2098),
.B(n_2021),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2111),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2119),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2114),
.B(n_2073),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_2109),
.B(n_2115),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2122),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2111),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2102),
.B(n_2025),
.Y(n_2184)
);

AOI21xp33_ASAP7_75t_L g2185 ( 
.A1(n_2160),
.A2(n_2106),
.B(n_2132),
.Y(n_2185)
);

OAI21xp33_ASAP7_75t_L g2186 ( 
.A1(n_2156),
.A2(n_2123),
.B(n_2099),
.Y(n_2186)
);

AOI221xp5_ASAP7_75t_L g2187 ( 
.A1(n_2152),
.A2(n_2142),
.B1(n_2132),
.B2(n_2117),
.C(n_2139),
.Y(n_2187)
);

NAND2x1_ASAP7_75t_L g2188 ( 
.A(n_2162),
.B(n_2100),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2168),
.B(n_2113),
.Y(n_2189)
);

OAI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2158),
.A2(n_2085),
.B1(n_2105),
.B2(n_2135),
.Y(n_2190)
);

NAND3x2_ASAP7_75t_L g2191 ( 
.A(n_2162),
.B(n_2135),
.C(n_2113),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2162),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_SL g2193 ( 
.A(n_2146),
.B(n_2105),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2153),
.Y(n_2194)
);

INVx1_ASAP7_75t_SL g2195 ( 
.A(n_2170),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2153),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2166),
.Y(n_2197)
);

AOI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_2143),
.A2(n_2134),
.B1(n_2078),
.B2(n_2140),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2167),
.B(n_2124),
.Y(n_2199)
);

OAI222xp33_ASAP7_75t_L g2200 ( 
.A1(n_2163),
.A2(n_2141),
.B1(n_2133),
.B2(n_2138),
.C1(n_2137),
.C2(n_2140),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2166),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2148),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2155),
.B(n_2112),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2172),
.B(n_2091),
.Y(n_2204)
);

O2A1O1Ixp33_ASAP7_75t_L g2205 ( 
.A1(n_2170),
.A2(n_2126),
.B(n_2131),
.C(n_2130),
.Y(n_2205)
);

OAI32xp33_ASAP7_75t_L g2206 ( 
.A1(n_2150),
.A2(n_2003),
.A3(n_2125),
.B1(n_2006),
.B2(n_1975),
.Y(n_2206)
);

AOI221xp5_ASAP7_75t_L g2207 ( 
.A1(n_2157),
.A2(n_2134),
.B1(n_2003),
.B2(n_2121),
.C(n_2120),
.Y(n_2207)
);

NAND2xp33_ASAP7_75t_SL g2208 ( 
.A(n_2173),
.B(n_1635),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2176),
.B(n_2155),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2148),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2173),
.A2(n_1985),
.B1(n_2016),
.B2(n_1984),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2149),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2149),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2165),
.B(n_1968),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2147),
.B(n_2026),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2151),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2203),
.B(n_2147),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2195),
.B(n_2147),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2192),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2188),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2194),
.Y(n_2221)
);

INVx2_ASAP7_75t_SL g2222 ( 
.A(n_2196),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2193),
.B(n_2175),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2197),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2209),
.B(n_2161),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2198),
.B(n_2175),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2189),
.B(n_2159),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2201),
.B(n_2169),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2202),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2199),
.B(n_2145),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_2186),
.B(n_2143),
.Y(n_2231)
);

AOI22xp5_ASAP7_75t_L g2232 ( 
.A1(n_2190),
.A2(n_2191),
.B1(n_2187),
.B2(n_2185),
.Y(n_2232)
);

NAND2x1_ASAP7_75t_L g2233 ( 
.A(n_2210),
.B(n_2144),
.Y(n_2233)
);

INVxp67_ASAP7_75t_L g2234 ( 
.A(n_2208),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_2204),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2205),
.B(n_2181),
.Y(n_2236)
);

INVx1_ASAP7_75t_SL g2237 ( 
.A(n_2208),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2207),
.B(n_2180),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2205),
.B(n_2181),
.Y(n_2239)
);

OR2x2_ASAP7_75t_L g2240 ( 
.A(n_2230),
.B(n_2145),
.Y(n_2240)
);

OAI21xp33_ASAP7_75t_L g2241 ( 
.A1(n_2232),
.A2(n_2190),
.B(n_2215),
.Y(n_2241)
);

NOR4xp25_ASAP7_75t_L g2242 ( 
.A(n_2236),
.B(n_2200),
.C(n_2216),
.D(n_2213),
.Y(n_2242)
);

AOI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_2239),
.A2(n_2200),
.B(n_2154),
.Y(n_2243)
);

AOI321xp33_ASAP7_75t_L g2244 ( 
.A1(n_2225),
.A2(n_2206),
.A3(n_2211),
.B1(n_2212),
.B2(n_2214),
.C(n_2144),
.Y(n_2244)
);

AOI21xp5_ASAP7_75t_L g2245 ( 
.A1(n_2231),
.A2(n_2184),
.B(n_2177),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2217),
.B(n_2180),
.Y(n_2246)
);

AOI221xp5_ASAP7_75t_L g2247 ( 
.A1(n_2235),
.A2(n_2151),
.B1(n_2182),
.B2(n_2179),
.C(n_2174),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2223),
.A2(n_2182),
.B1(n_2164),
.B2(n_2178),
.Y(n_2248)
);

AOI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_2233),
.A2(n_2218),
.B(n_2223),
.Y(n_2249)
);

AOI221x1_ASAP7_75t_L g2250 ( 
.A1(n_2221),
.A2(n_2183),
.B1(n_2178),
.B2(n_2120),
.C(n_2121),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2222),
.Y(n_2251)
);

AOI322xp5_ASAP7_75t_L g2252 ( 
.A1(n_2238),
.A2(n_2183),
.A3(n_2019),
.B1(n_2002),
.B2(n_2008),
.C1(n_1975),
.C2(n_2129),
.Y(n_2252)
);

AOI21xp5_ASAP7_75t_L g2253 ( 
.A1(n_2233),
.A2(n_2164),
.B(n_2171),
.Y(n_2253)
);

OAI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2220),
.A2(n_2171),
.B(n_2129),
.Y(n_2254)
);

AOI211xp5_ASAP7_75t_L g2255 ( 
.A1(n_2220),
.A2(n_2082),
.B(n_2079),
.C(n_2056),
.Y(n_2255)
);

NOR3xp33_ASAP7_75t_L g2256 ( 
.A(n_2241),
.B(n_2219),
.C(n_2227),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_2249),
.B(n_2226),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2240),
.Y(n_2258)
);

NOR3xp33_ASAP7_75t_L g2259 ( 
.A(n_2243),
.B(n_2219),
.C(n_2226),
.Y(n_2259)
);

NAND3xp33_ASAP7_75t_L g2260 ( 
.A(n_2242),
.B(n_2234),
.C(n_2224),
.Y(n_2260)
);

NOR2x1_ASAP7_75t_L g2261 ( 
.A(n_2251),
.B(n_2229),
.Y(n_2261)
);

NOR2x1p5_ASAP7_75t_L g2262 ( 
.A(n_2246),
.B(n_2230),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2245),
.B(n_2217),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2248),
.Y(n_2264)
);

NOR3xp33_ASAP7_75t_L g2265 ( 
.A(n_2247),
.B(n_2228),
.C(n_2222),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2254),
.Y(n_2266)
);

AO22x2_ASAP7_75t_L g2267 ( 
.A1(n_2253),
.A2(n_2229),
.B1(n_2221),
.B2(n_2237),
.Y(n_2267)
);

NAND3xp33_ASAP7_75t_L g2268 ( 
.A(n_2244),
.B(n_2252),
.C(n_2250),
.Y(n_2268)
);

AOI221xp5_ASAP7_75t_L g2269 ( 
.A1(n_2268),
.A2(n_2238),
.B1(n_2255),
.B2(n_2003),
.C(n_2079),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2259),
.B(n_2010),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2262),
.B(n_2027),
.Y(n_2271)
);

NAND3xp33_ASAP7_75t_SL g2272 ( 
.A(n_2256),
.B(n_2265),
.C(n_2257),
.Y(n_2272)
);

NAND4xp25_ASAP7_75t_L g2273 ( 
.A(n_2260),
.B(n_1575),
.C(n_2082),
.D(n_2067),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2258),
.B(n_2014),
.Y(n_2274)
);

OAI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2266),
.A2(n_2003),
.B(n_2002),
.Y(n_2275)
);

OAI211xp5_ASAP7_75t_SL g2276 ( 
.A1(n_2263),
.A2(n_1991),
.B(n_2005),
.C(n_1992),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2267),
.B(n_2014),
.Y(n_2277)
);

NOR2x2_ASAP7_75t_L g2278 ( 
.A(n_2272),
.B(n_2267),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2271),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2270),
.Y(n_2280)
);

NOR2x1_ASAP7_75t_L g2281 ( 
.A(n_2273),
.B(n_2261),
.Y(n_2281)
);

NOR2x1p5_ASAP7_75t_L g2282 ( 
.A(n_2277),
.B(n_2264),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2274),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2269),
.B(n_1970),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2276),
.A2(n_2008),
.B1(n_2024),
.B2(n_2020),
.Y(n_2285)
);

NOR2x1_ASAP7_75t_L g2286 ( 
.A(n_2275),
.B(n_1984),
.Y(n_2286)
);

OR2x2_ASAP7_75t_L g2287 ( 
.A(n_2279),
.B(n_2016),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_2281),
.B(n_2072),
.Y(n_2288)
);

NOR3xp33_ASAP7_75t_L g2289 ( 
.A(n_2280),
.B(n_1991),
.C(n_1735),
.Y(n_2289)
);

AND3x4_ASAP7_75t_L g2290 ( 
.A(n_2286),
.B(n_2278),
.C(n_2282),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2284),
.B(n_1970),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2283),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2285),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2290),
.Y(n_2294)
);

OAI22x1_ASAP7_75t_SL g2295 ( 
.A1(n_2292),
.A2(n_2000),
.B1(n_1999),
.B2(n_1984),
.Y(n_2295)
);

NOR2x1_ASAP7_75t_L g2296 ( 
.A(n_2288),
.B(n_1975),
.Y(n_2296)
);

OR2x2_ASAP7_75t_L g2297 ( 
.A(n_2287),
.B(n_1999),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2294),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2297),
.Y(n_2299)
);

AOI221xp5_ASAP7_75t_L g2300 ( 
.A1(n_2298),
.A2(n_2288),
.B1(n_2293),
.B2(n_2289),
.C(n_2295),
.Y(n_2300)
);

OR3x1_ASAP7_75t_L g2301 ( 
.A(n_2299),
.B(n_2296),
.C(n_2291),
.Y(n_2301)
);

OAI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_2300),
.A2(n_1585),
.B1(n_1984),
.B2(n_1645),
.Y(n_2302)
);

AOI21xp5_ASAP7_75t_L g2303 ( 
.A1(n_2301),
.A2(n_1585),
.B(n_2000),
.Y(n_2303)
);

AOI22x1_ASAP7_75t_L g2304 ( 
.A1(n_2303),
.A2(n_1645),
.B1(n_1735),
.B2(n_1736),
.Y(n_2304)
);

AO21x2_ASAP7_75t_L g2305 ( 
.A1(n_2302),
.A2(n_2072),
.B(n_1849),
.Y(n_2305)
);

AOI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_2304),
.A2(n_1585),
.B1(n_2024),
.B2(n_2020),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_2305),
.A2(n_2004),
.B1(n_1996),
.B2(n_1977),
.Y(n_2307)
);

OAI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_2307),
.A2(n_2305),
.B(n_1983),
.Y(n_2308)
);

AOI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2308),
.A2(n_2306),
.B1(n_2004),
.B2(n_1996),
.Y(n_2309)
);

OAI221xp5_ASAP7_75t_R g2310 ( 
.A1(n_2309),
.A2(n_1869),
.B1(n_1854),
.B2(n_1858),
.C(n_1645),
.Y(n_2310)
);

AOI211xp5_ASAP7_75t_L g2311 ( 
.A1(n_2310),
.A2(n_1645),
.B(n_1788),
.C(n_1983),
.Y(n_2311)
);


endmodule