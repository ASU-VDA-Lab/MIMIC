module real_aes_17731_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_0), .Y(n_179) );
AND2x4_ASAP7_75t_L g865 ( .A(n_1), .B(n_866), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_2), .A2(n_104), .B1(n_853), .B2(n_854), .Y(n_852) );
INVxp33_ASAP7_75t_R g853 ( .A(n_2), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_2), .B(n_876), .Y(n_875) );
BUFx3_ASAP7_75t_L g224 ( .A(n_3), .Y(n_224) );
INVx1_ASAP7_75t_L g866 ( .A(n_4), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_5), .B(n_240), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g101 ( .A1(n_6), .A2(n_102), .B1(n_816), .B2(n_817), .Y(n_101) );
INVx1_ASAP7_75t_L g816 ( .A(n_6), .Y(n_816) );
OR2x2_ASAP7_75t_L g826 ( .A(n_7), .B(n_22), .Y(n_826) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_8), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_9), .B(n_124), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_10), .B(n_124), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_11), .B(n_151), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_12), .A2(n_79), .B1(n_120), .B2(n_124), .Y(n_123) );
OAI21x1_ASAP7_75t_L g113 ( .A1(n_13), .A2(n_36), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_14), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_15), .B(n_160), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_16), .Y(n_547) );
AO32x2_ASAP7_75t_L g111 ( .A1(n_17), .A2(n_112), .A3(n_115), .B1(n_126), .B2(n_130), .Y(n_111) );
AO32x1_ASAP7_75t_L g256 ( .A1(n_17), .A2(n_112), .A3(n_115), .B1(n_126), .B2(n_130), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_18), .B(n_479), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_19), .B(n_130), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g859 ( .A(n_20), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_21), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_23), .A2(n_42), .B1(n_160), .B2(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_24), .B(n_141), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_25), .A2(n_87), .B1(n_120), .B2(n_122), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_26), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_27), .B(n_139), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_28), .A2(n_61), .B1(n_122), .B2(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_29), .B(n_124), .Y(n_580) );
INVx2_ASAP7_75t_L g821 ( .A(n_30), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_31), .B(n_125), .Y(n_489) );
BUFx3_ASAP7_75t_L g824 ( .A(n_32), .Y(n_824) );
INVx1_ASAP7_75t_L g850 ( .A(n_32), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_33), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_34), .B(n_496), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_35), .Y(n_828) );
AND2x2_ASAP7_75t_L g552 ( .A(n_37), .B(n_496), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_38), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_39), .B(n_180), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_40), .B(n_479), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_41), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_43), .B(n_566), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_44), .A2(n_74), .B1(n_139), .B2(n_180), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_45), .B(n_159), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_46), .A2(n_116), .B(n_177), .C(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_47), .A2(n_76), .B1(n_120), .B2(n_124), .Y(n_220) );
INVx1_ASAP7_75t_L g114 ( .A(n_48), .Y(n_114) );
AND2x4_ASAP7_75t_L g128 ( .A(n_49), .B(n_129), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_50), .A2(n_51), .B1(n_122), .B2(n_162), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_52), .B(n_130), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_53), .B(n_496), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_54), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_55), .B(n_122), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_56), .B(n_120), .Y(n_238) );
INVx1_ASAP7_75t_L g129 ( .A(n_57), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_58), .B(n_130), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_59), .A2(n_143), .B(n_177), .C(n_178), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g244 ( .A(n_60), .B(n_120), .C(n_243), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_62), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_63), .B(n_130), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_64), .B(n_504), .Y(n_515) );
AND2x2_ASAP7_75t_L g182 ( .A(n_65), .B(n_183), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_66), .Y(n_164) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_67), .B(n_125), .C(n_160), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_68), .A2(n_90), .B1(n_124), .B2(n_180), .Y(n_211) );
INVx2_ASAP7_75t_L g118 ( .A(n_69), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_70), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_71), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_72), .B(n_175), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_73), .B(n_124), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_75), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_77), .B(n_199), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_78), .A2(n_86), .B1(n_478), .B2(n_479), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_80), .B(n_124), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_81), .B(n_243), .Y(n_242) );
NAND2xp33_ASAP7_75t_SL g531 ( .A(n_82), .B(n_240), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_83), .B(n_195), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_84), .A2(n_97), .B1(n_122), .B2(n_162), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_85), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g466 ( .A(n_88), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_88), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_89), .B(n_151), .Y(n_150) );
NAND2xp33_ASAP7_75t_L g505 ( .A(n_91), .B(n_240), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_92), .B(n_496), .Y(n_520) );
NAND3xp33_ASAP7_75t_L g528 ( .A(n_93), .B(n_175), .C(n_240), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_94), .B(n_504), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_95), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_96), .B(n_479), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_836), .B(n_860), .C(n_868), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_100), .Y(n_99) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_818), .B(n_827), .Y(n_100) );
INVx2_ASAP7_75t_L g817 ( .A(n_102), .Y(n_817) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_463), .B1(n_467), .B2(n_468), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g854 ( .A(n_104), .Y(n_854) );
NOR2x1p5_ASAP7_75t_L g104 ( .A(n_105), .B(n_371), .Y(n_104) );
NAND4xp75_ASAP7_75t_L g105 ( .A(n_106), .B(n_268), .C(n_302), .D(n_351), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_185), .B(n_225), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_131), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g347 ( .A(n_110), .Y(n_347) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g230 ( .A(n_111), .B(n_133), .Y(n_230) );
AND2x4_ASAP7_75t_L g263 ( .A(n_111), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g284 ( .A(n_111), .Y(n_284) );
INVx4_ASAP7_75t_L g130 ( .A(n_112), .Y(n_130) );
INVx2_ASAP7_75t_SL g135 ( .A(n_112), .Y(n_135) );
BUFx3_ASAP7_75t_L g156 ( .A(n_112), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_112), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g190 ( .A(n_112), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_112), .B(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_SL g510 ( .A(n_112), .B(n_203), .Y(n_510) );
INVx1_ASAP7_75t_SL g524 ( .A(n_112), .Y(n_524) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g153 ( .A(n_113), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_119), .B1(n_123), .B2(n_125), .Y(n_115) );
O2A1O1Ixp5_ASAP7_75t_L g192 ( .A1(n_116), .A2(n_193), .B(n_194), .C(n_196), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_116), .A2(n_503), .B(n_505), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_116), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_116), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_116), .A2(n_579), .B(n_580), .Y(n_578) );
BUFx4f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g243 ( .A(n_117), .Y(n_243) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx8_ASAP7_75t_L g125 ( .A(n_118), .Y(n_125) );
INVx2_ASAP7_75t_L g144 ( .A(n_118), .Y(n_144) );
INVx1_ASAP7_75t_L g175 ( .A(n_118), .Y(n_175) );
INVx2_ASAP7_75t_SL g139 ( .A(n_120), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_120), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_121), .Y(n_122) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_121), .Y(n_124) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
INVx1_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
INVx1_ASAP7_75t_L g177 ( .A(n_121), .Y(n_177) );
INVx1_ASAP7_75t_L g180 ( .A(n_121), .Y(n_180) );
INVx1_ASAP7_75t_L g195 ( .A(n_121), .Y(n_195) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_121), .Y(n_240) );
INVx1_ASAP7_75t_L g480 ( .A(n_121), .Y(n_480) );
INVx3_ASAP7_75t_L g504 ( .A(n_121), .Y(n_504) );
INVx2_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
INVx2_ASAP7_75t_L g478 ( .A(n_122), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_122), .A2(n_489), .B(n_490), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_122), .A2(n_504), .B1(n_550), .B2(n_551), .Y(n_549) );
INVx3_ASAP7_75t_L g148 ( .A(n_124), .Y(n_148) );
INVx1_ASAP7_75t_L g494 ( .A(n_124), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_124), .A2(n_527), .B(n_528), .Y(n_526) );
INVx6_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_125), .A2(n_149), .B1(n_220), .B2(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_125), .A2(n_238), .B(n_239), .Y(n_237) );
O2A1O1Ixp5_ASAP7_75t_L g560 ( .A1(n_125), .A2(n_194), .B(n_561), .C(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_125), .A2(n_582), .B(n_583), .Y(n_581) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_126), .A2(n_137), .B(n_145), .Y(n_136) );
INVx2_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_SL g212 ( .A(n_127), .Y(n_212) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AO31x2_ASAP7_75t_L g155 ( .A1(n_128), .A2(n_156), .A3(n_157), .B(n_163), .Y(n_155) );
INVx1_ASAP7_75t_L g181 ( .A(n_128), .Y(n_181) );
BUFx10_ASAP7_75t_L g203 ( .A(n_128), .Y(n_203) );
BUFx10_ASAP7_75t_L g483 ( .A(n_128), .Y(n_483) );
INVx2_ASAP7_75t_L g218 ( .A(n_130), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_131), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_154), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_132), .B(n_298), .Y(n_375) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_132), .Y(n_402) );
OR2x2_ASAP7_75t_L g451 ( .A(n_132), .B(n_255), .Y(n_451) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g267 ( .A(n_133), .Y(n_267) );
INVx3_ASAP7_75t_L g275 ( .A(n_133), .Y(n_275) );
OR2x2_ASAP7_75t_L g283 ( .A(n_133), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g311 ( .A(n_133), .B(n_281), .Y(n_311) );
INVx1_ASAP7_75t_L g322 ( .A(n_133), .Y(n_322) );
AND2x2_ASAP7_75t_L g343 ( .A(n_133), .B(n_284), .Y(n_343) );
INVxp67_ASAP7_75t_L g367 ( .A(n_133), .Y(n_367) );
BUFx2_ASAP7_75t_L g411 ( .A(n_133), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_133), .B(n_155), .Y(n_420) );
AND2x2_ASAP7_75t_L g427 ( .A(n_133), .B(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_150), .Y(n_134) );
AOI21x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_142), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_141), .A2(n_242), .B(n_244), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_142), .A2(n_149), .B1(n_158), .B2(n_161), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_142), .A2(n_518), .B(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g482 ( .A(n_143), .Y(n_482) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g200 ( .A(n_144), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_149), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_149), .A2(n_209), .B1(n_210), .B2(n_211), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_149), .A2(n_477), .B1(n_481), .B2(n_482), .Y(n_476) );
INVx2_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
NOR2xp67_ASAP7_75t_SL g542 ( .A(n_151), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AO31x2_ASAP7_75t_L g475 ( .A1(n_152), .A2(n_476), .A3(n_483), .B(n_484), .Y(n_475) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx2_ASAP7_75t_L g235 ( .A(n_153), .Y(n_235) );
AND2x2_ASAP7_75t_L g285 ( .A(n_154), .B(n_286), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_154), .A2(n_188), .B1(n_401), .B2(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_165), .Y(n_154) );
OR2x2_ASAP7_75t_L g255 ( .A(n_155), .B(n_256), .Y(n_255) );
INVx3_ASAP7_75t_L g264 ( .A(n_155), .Y(n_264) );
AND2x2_ASAP7_75t_L g276 ( .A(n_155), .B(n_256), .Y(n_276) );
AND2x2_ASAP7_75t_L g334 ( .A(n_155), .B(n_166), .Y(n_334) );
AO31x2_ASAP7_75t_L g207 ( .A1(n_156), .A2(n_208), .A3(n_212), .B(n_213), .Y(n_207) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_160), .A2(n_162), .B1(n_172), .B2(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g201 ( .A(n_162), .Y(n_201) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
INVx1_ASAP7_75t_L g325 ( .A(n_166), .Y(n_325) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_166), .Y(n_428) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g281 ( .A(n_167), .Y(n_281) );
AOI21x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_182), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_176), .B(n_181), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_171), .B(n_174), .Y(n_170) );
AOI21x1_ASAP7_75t_L g491 ( .A1(n_174), .A2(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_SL g210 ( .A(n_175), .Y(n_210) );
INVx1_ASAP7_75t_L g508 ( .A(n_177), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_184), .B(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_184), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_205), .Y(n_186) );
AND2x2_ASAP7_75t_L g382 ( .A(n_187), .B(n_328), .Y(n_382) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI32xp33_ASAP7_75t_L g412 ( .A1(n_188), .A2(n_305), .A3(n_379), .B1(n_413), .B2(n_415), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_188), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
OR2x2_ASAP7_75t_L g232 ( .A(n_189), .B(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g251 ( .A(n_189), .B(n_207), .Y(n_251) );
BUFx2_ASAP7_75t_L g270 ( .A(n_189), .Y(n_270) );
INVx1_ASAP7_75t_L g317 ( .A(n_189), .Y(n_317) );
AND2x2_ASAP7_75t_L g350 ( .A(n_189), .B(n_329), .Y(n_350) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_204), .Y(n_189) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_190), .A2(n_191), .B(n_204), .Y(n_296) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_190), .A2(n_487), .B(n_495), .Y(n_486) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_190), .A2(n_487), .B(n_495), .Y(n_574) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_190), .A2(n_577), .B(n_584), .Y(n_576) );
OAI21x1_ASAP7_75t_L g624 ( .A1(n_190), .A2(n_577), .B(n_584), .Y(n_624) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_197), .B(n_203), .Y(n_191) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_199), .A2(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_200), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_506) );
AOI31xp67_ASAP7_75t_L g217 ( .A1(n_203), .A2(n_218), .A3(n_219), .B(n_222), .Y(n_217) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_203), .A2(n_237), .B(n_241), .Y(n_236) );
OAI21x1_ASAP7_75t_L g487 ( .A1(n_203), .A2(n_488), .B(n_491), .Y(n_487) );
OAI21x1_ASAP7_75t_L g513 ( .A1(n_203), .A2(n_514), .B(n_517), .Y(n_513) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_203), .A2(n_526), .B(n_529), .Y(n_525) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_203), .A2(n_560), .B(n_563), .Y(n_559) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_203), .A2(n_578), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g231 ( .A(n_206), .B(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g438 ( .A(n_206), .B(n_322), .Y(n_438) );
INVx1_ASAP7_75t_L g442 ( .A(n_206), .Y(n_442) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_215), .Y(n_206) );
INVx2_ASAP7_75t_L g266 ( .A(n_207), .Y(n_266) );
AND2x2_ASAP7_75t_L g290 ( .A(n_207), .B(n_249), .Y(n_290) );
AND2x2_ASAP7_75t_L g301 ( .A(n_207), .B(n_296), .Y(n_301) );
INVx1_ASAP7_75t_L g308 ( .A(n_207), .Y(n_308) );
AND2x2_ASAP7_75t_L g316 ( .A(n_207), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g329 ( .A(n_207), .Y(n_329) );
AND2x2_ASAP7_75t_L g395 ( .A(n_207), .B(n_215), .Y(n_395) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g259 ( .A(n_216), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g249 ( .A(n_217), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
OAI221xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_231), .B1(n_246), .B2(n_252), .C(n_257), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_227), .A2(n_379), .B(n_382), .Y(n_378) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
AND2x4_ASAP7_75t_L g454 ( .A(n_228), .B(n_254), .Y(n_454) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x4_ASAP7_75t_L g298 ( .A(n_229), .B(n_264), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_230), .B(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_L g363 ( .A(n_230), .Y(n_363) );
OR2x2_ASAP7_75t_L g307 ( .A(n_232), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g369 ( .A(n_232), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g440 ( .A(n_232), .Y(n_440) );
AND2x2_ASAP7_75t_L g248 ( .A(n_233), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g397 ( .A(n_233), .B(n_296), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_236), .B(n_245), .Y(n_233) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_234), .A2(n_236), .B(n_245), .Y(n_260) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_234), .A2(n_513), .B(n_520), .Y(n_512) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_234), .A2(n_559), .B(n_567), .Y(n_558) );
OAI21xp33_ASAP7_75t_SL g620 ( .A1(n_234), .A2(n_513), .B(n_520), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_234), .A2(n_559), .B(n_567), .Y(n_630) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g496 ( .A(n_235), .Y(n_496) );
INVx2_ASAP7_75t_L g566 ( .A(n_240), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g277 ( .A1(n_246), .A2(n_278), .B1(n_279), .B2(n_288), .C(n_297), .Y(n_277) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_246), .A2(n_361), .B1(n_374), .B2(n_376), .C(n_378), .Y(n_373) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
AND2x2_ASAP7_75t_L g300 ( .A(n_248), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g313 ( .A(n_249), .B(n_296), .Y(n_313) );
INVx2_ASAP7_75t_L g319 ( .A(n_249), .Y(n_319) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_252), .A2(n_384), .B1(n_389), .B2(n_393), .C(n_398), .Y(n_383) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g435 ( .A(n_255), .B(n_405), .Y(n_435) );
INVx1_ASAP7_75t_L g287 ( .A(n_256), .Y(n_287) );
INVx1_ASAP7_75t_L g324 ( .A(n_256), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_261), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g273 ( .A(n_259), .Y(n_273) );
OR2x2_ASAP7_75t_L g336 ( .A(n_259), .B(n_272), .Y(n_336) );
INVx2_ASAP7_75t_L g349 ( .A(n_259), .Y(n_349) );
INVx2_ASAP7_75t_L g294 ( .A(n_260), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx2_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
AND2x4_ASAP7_75t_L g305 ( .A(n_263), .B(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_263), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g379 ( .A(n_263), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g456 ( .A(n_263), .B(n_411), .Y(n_456) );
AND2x2_ASAP7_75t_L g280 ( .A(n_264), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
INVx1_ASAP7_75t_L g401 ( .A(n_264), .Y(n_401) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_SL g272 ( .A(n_266), .Y(n_272) );
AND2x2_ASAP7_75t_L g314 ( .A(n_266), .B(n_293), .Y(n_314) );
AND2x2_ASAP7_75t_L g388 ( .A(n_267), .B(n_342), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_274), .B(n_277), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g354 ( .A(n_270), .Y(n_354) );
AND2x2_ASAP7_75t_L g421 ( .A(n_270), .B(n_349), .Y(n_421) );
AND2x2_ASAP7_75t_L g436 ( .A(n_270), .B(n_395), .Y(n_436) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g390 ( .A(n_272), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_272), .B(n_397), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g444 ( .A1(n_272), .A2(n_346), .A3(n_414), .B1(n_445), .B2(n_446), .B3(n_447), .Y(n_444) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_275), .B(n_281), .Y(n_405) );
AND2x2_ASAP7_75t_L g433 ( .A(n_276), .B(n_381), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_282), .B(n_285), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
INVx1_ASAP7_75t_L g381 ( .A(n_281), .Y(n_381) );
OAI32xp33_ASAP7_75t_L g326 ( .A1(n_282), .A2(n_307), .A3(n_327), .B1(n_330), .B2(n_332), .Y(n_326) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g361 ( .A(n_283), .B(n_306), .Y(n_361) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
INVx2_ASAP7_75t_L g387 ( .A(n_287), .Y(n_387) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g370 ( .A(n_290), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_291), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g430 ( .A(n_291), .B(n_377), .Y(n_430) );
INVx2_ASAP7_75t_L g461 ( .A(n_291), .Y(n_461) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g376 ( .A(n_292), .B(n_377), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
AND2x2_ASAP7_75t_L g318 ( .A(n_293), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g360 ( .A(n_294), .Y(n_360) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_300), .Y(n_297) );
INVx2_ASAP7_75t_L g368 ( .A(n_298), .Y(n_368) );
AND2x2_ASAP7_75t_L g352 ( .A(n_299), .B(n_353), .Y(n_352) );
NOR3x1_ASAP7_75t_L g302 ( .A(n_303), .B(n_326), .C(n_335), .Y(n_302) );
OAI21xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_307), .B(n_309), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_306), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_308), .B(n_359), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B1(n_315), .B2(n_320), .Y(n_309) );
INVx3_ASAP7_75t_L g344 ( .A(n_311), .Y(n_344) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVxp67_ASAP7_75t_L g357 ( .A(n_313), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_313), .B(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
AND2x2_ASAP7_75t_L g458 ( .A(n_316), .B(n_349), .Y(n_458) );
AND2x2_ASAP7_75t_L g328 ( .A(n_319), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g377 ( .A(n_319), .Y(n_377) );
INVx1_ASAP7_75t_L g414 ( .A(n_319), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_319), .B(n_360), .Y(n_448) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g445 ( .A(n_323), .Y(n_445) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g331 ( .A(n_325), .Y(n_331) );
AND2x2_ASAP7_75t_L g457 ( .A(n_328), .B(n_397), .Y(n_457) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
AND2x2_ASAP7_75t_L g462 ( .A(n_334), .B(n_343), .Y(n_462) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_345), .B2(n_348), .Y(n_335) );
AOI211xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_340), .B(n_343), .C(n_344), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g419 ( .A(n_339), .B(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVxp33_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g353 ( .A(n_349), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g431 ( .A(n_350), .B(n_392), .Y(n_431) );
INVx1_ASAP7_75t_L g446 ( .A(n_350), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .C(n_362), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_361), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g392 ( .A(n_360), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B(n_366), .C(n_369), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_363), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_423), .Y(n_371) );
NOR3xp33_ASAP7_75t_SL g372 ( .A(n_373), .B(n_383), .C(n_408), .Y(n_372) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_379), .A2(n_418), .B1(n_421), .B2(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
AND2x2_ASAP7_75t_L g403 ( .A(n_386), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g426 ( .A(n_386), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g422 ( .A(n_391), .Y(n_422) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_397), .B(n_414), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .B(n_406), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_403), .A2(n_458), .B1(n_460), .B2(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI21xp33_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_412), .B(n_417), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_410), .B(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g449 ( .A(n_420), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_422), .A2(n_444), .B1(n_449), .B2(n_450), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_452), .Y(n_423) );
OAI211xp5_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_429), .B(n_432), .C(n_443), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
O2A1O1Ixp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_436), .C(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_435), .A2(n_438), .B1(n_439), .B2(n_441), .Y(n_437) );
OAI211xp5_ASAP7_75t_L g452 ( .A1(n_446), .A2(n_453), .B(n_455), .C(n_459), .Y(n_452) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx4_ASAP7_75t_L g467 ( .A(n_463), .Y(n_467) );
BUFx12f_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g834 ( .A(n_465), .B(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_704), .Y(n_468) );
NAND4xp25_ASAP7_75t_L g469 ( .A(n_470), .B(n_611), .C(n_652), .D(n_684), .Y(n_469) );
NOR2xp33_ASAP7_75t_SL g470 ( .A(n_471), .B(n_590), .Y(n_470) );
NAND3xp33_ASAP7_75t_SL g471 ( .A(n_472), .B(n_553), .C(n_570), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_497), .B1(n_533), .B2(n_537), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_473), .B(n_597), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_473), .B(n_697), .Y(n_803) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g555 ( .A(n_474), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_486), .Y(n_474) );
OR2x2_ASAP7_75t_L g536 ( .A(n_475), .B(n_486), .Y(n_536) );
INVx1_ASAP7_75t_L g600 ( .A(n_475), .Y(n_600) );
AND2x2_ASAP7_75t_L g603 ( .A(n_475), .B(n_574), .Y(n_603) );
AND2x2_ASAP7_75t_L g651 ( .A(n_475), .B(n_624), .Y(n_651) );
AND2x2_ASAP7_75t_L g659 ( .A(n_475), .B(n_633), .Y(n_659) );
OR2x2_ASAP7_75t_L g670 ( .A(n_475), .B(n_624), .Y(n_670) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_475), .Y(n_710) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_482), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g543 ( .A(n_483), .Y(n_543) );
AND2x2_ASAP7_75t_L g629 ( .A(n_486), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g658 ( .A(n_486), .B(n_557), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_497), .A2(n_629), .B(n_765), .Y(n_770) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_521), .Y(n_497) );
AND2x2_ASAP7_75t_L g537 ( .A(n_498), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g568 ( .A(n_498), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_498), .B(n_666), .Y(n_665) );
NAND2xp33_ASAP7_75t_R g700 ( .A(n_498), .B(n_666), .Y(n_700) );
INVx1_ASAP7_75t_L g734 ( .A(n_498), .Y(n_734) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_498), .Y(n_784) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_511), .Y(n_498) );
INVx1_ASAP7_75t_L g587 ( .A(n_499), .Y(n_587) );
INVx4_ASAP7_75t_L g608 ( .A(n_499), .Y(n_608) );
OR2x2_ASAP7_75t_L g691 ( .A(n_499), .B(n_616), .Y(n_691) );
BUFx2_ASAP7_75t_L g760 ( .A(n_499), .Y(n_760) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
OAI21x1_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_506), .B(n_510), .Y(n_501) );
AND2x2_ASAP7_75t_L g588 ( .A(n_511), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g675 ( .A(n_511), .Y(n_675) );
AND2x2_ASAP7_75t_L g761 ( .A(n_511), .B(n_569), .Y(n_761) );
AND2x2_ASAP7_75t_L g783 ( .A(n_511), .B(n_608), .Y(n_783) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g638 ( .A(n_512), .Y(n_638) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g586 ( .A(n_522), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g609 ( .A(n_522), .Y(n_609) );
INVx1_ASAP7_75t_L g646 ( .A(n_522), .Y(n_646) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g616 ( .A(n_523), .Y(n_616) );
AND2x2_ASAP7_75t_L g673 ( .A(n_523), .B(n_541), .Y(n_673) );
OAI21x1_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_532), .Y(n_523) );
NOR2xp33_ASAP7_75t_SL g668 ( .A(n_533), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g715 ( .A(n_535), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g731 ( .A(n_536), .B(n_597), .Y(n_731) );
INVx1_ASAP7_75t_L g739 ( .A(n_536), .Y(n_739) );
OR2x2_ASAP7_75t_L g660 ( .A(n_538), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_539), .Y(n_610) );
INVx1_ASAP7_75t_L g768 ( .A(n_539), .Y(n_768) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g569 ( .A(n_540), .Y(n_569) );
AND2x2_ASAP7_75t_L g666 ( .A(n_540), .B(n_609), .Y(n_666) );
INVx2_ASAP7_75t_L g725 ( .A(n_540), .Y(n_725) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g589 ( .A(n_541), .Y(n_589) );
AOI21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_544), .B(n_552), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_548), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_568), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g679 ( .A(n_556), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_556), .B(n_603), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_556), .B(n_669), .Y(n_775) );
AND2x2_ASAP7_75t_L g801 ( .A(n_556), .B(n_659), .Y(n_801) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_557), .Y(n_572) );
INVxp67_ASAP7_75t_SL g594 ( .A(n_557), .Y(n_594) );
AND2x2_ASAP7_75t_L g627 ( .A(n_557), .B(n_574), .Y(n_627) );
INVx1_ASAP7_75t_L g698 ( .A(n_557), .Y(n_698) );
INVx1_ASAP7_75t_L g713 ( .A(n_557), .Y(n_713) );
AND2x2_ASAP7_75t_L g765 ( .A(n_557), .B(n_718), .Y(n_765) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g636 ( .A(n_569), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g643 ( .A(n_569), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_569), .B(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g812 ( .A(n_569), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_585), .Y(n_570) );
INVx1_ASAP7_75t_L g641 ( .A(n_571), .Y(n_641) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND2x1_ASAP7_75t_L g815 ( .A(n_572), .B(n_715), .Y(n_815) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g599 ( .A(n_574), .Y(n_599) );
AND2x2_ASAP7_75t_L g664 ( .A(n_574), .B(n_630), .Y(n_664) );
INVx1_ASAP7_75t_L g678 ( .A(n_574), .Y(n_678) );
INVx3_ASAP7_75t_L g597 ( .A(n_575), .Y(n_597) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g633 ( .A(n_576), .Y(n_633) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g661 ( .A(n_586), .Y(n_661) );
AND2x2_ASAP7_75t_L g688 ( .A(n_586), .B(n_619), .Y(n_688) );
AND2x2_ASAP7_75t_L g749 ( .A(n_586), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g811 ( .A(n_586), .B(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g692 ( .A(n_588), .Y(n_692) );
AND2x2_ASAP7_75t_L g720 ( .A(n_588), .B(n_609), .Y(n_720) );
AND2x2_ASAP7_75t_L g619 ( .A(n_589), .B(n_620), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_601), .B(n_604), .Y(n_590) );
OAI22xp5_ASAP7_75t_SL g809 ( .A1(n_591), .A2(n_810), .B1(n_813), .B2(n_815), .Y(n_809) );
NAND2x1p5_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2x1_ASAP7_75t_L g794 ( .A(n_593), .B(n_595), .Y(n_794) );
BUFx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_596), .B(n_658), .Y(n_703) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g602 ( .A(n_597), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_597), .B(n_678), .Y(n_677) );
AND2x4_ASAP7_75t_L g755 ( .A(n_598), .B(n_713), .Y(n_755) );
INVx1_ASAP7_75t_L g808 ( .A(n_598), .Y(n_808) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g623 ( .A(n_600), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_610), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g618 ( .A(n_607), .Y(n_618) );
AND2x2_ASAP7_75t_L g682 ( .A(n_607), .B(n_683), .Y(n_682) );
AND3x2_ASAP7_75t_L g724 ( .A(n_607), .B(n_637), .C(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_607), .B(n_725), .Y(n_781) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g645 ( .A(n_608), .B(n_646), .Y(n_645) );
NAND2x1_ASAP7_75t_L g674 ( .A(n_608), .B(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g729 ( .A(n_608), .Y(n_729) );
AND2x2_ASAP7_75t_L g790 ( .A(n_608), .B(n_725), .Y(n_790) );
OR2x2_ASAP7_75t_L g769 ( .A(n_609), .B(n_638), .Y(n_769) );
INVx1_ASAP7_75t_L g730 ( .A(n_610), .Y(n_730) );
AOI321xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_621), .A3(n_625), .B1(n_628), .B2(n_634), .C(n_640), .Y(n_611) );
AOI211xp5_ASAP7_75t_SL g652 ( .A1(n_612), .A2(n_653), .B(n_655), .C(n_667), .Y(n_652) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g778 ( .A(n_614), .B(n_717), .C(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g793 ( .A(n_614), .Y(n_793) );
BUFx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g637 ( .A(n_616), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g787 ( .A(n_616), .B(n_751), .Y(n_787) );
INVx1_ASAP7_75t_L g639 ( .A(n_617), .Y(n_639) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
BUFx2_ASAP7_75t_L g796 ( .A(n_618), .Y(n_796) );
INVx1_ASAP7_75t_L g649 ( .A(n_619), .Y(n_649) );
AND2x2_ASAP7_75t_L g776 ( .A(n_619), .B(n_760), .Y(n_776) );
BUFx2_ASAP7_75t_L g799 ( .A(n_620), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_621), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g718 ( .A(n_624), .Y(n_718) );
OAI321xp33_ASAP7_75t_L g762 ( .A1(n_625), .A2(n_716), .A3(n_763), .B1(n_764), .B2(n_767), .C(n_770), .Y(n_762) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g687 ( .A(n_627), .B(n_631), .Y(n_687) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_629), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g751 ( .A(n_630), .Y(n_751) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_639), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g789 ( .A(n_637), .B(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g683 ( .A(n_638), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_647), .B2(n_650), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI31xp33_ASAP7_75t_L g727 ( .A1(n_643), .A2(n_679), .A3(n_728), .B(n_730), .Y(n_727) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g742 ( .A(n_645), .Y(n_742) );
OR2x2_ASAP7_75t_L g763 ( .A(n_645), .B(n_649), .Y(n_763) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx2_ASAP7_75t_L g695 ( .A(n_651), .Y(n_695) );
INVx1_ASAP7_75t_L g753 ( .A(n_651), .Y(n_753) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_660), .B1(n_662), .B2(n_665), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_L g747 ( .A(n_659), .Y(n_747) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_663), .A2(n_694), .B(n_696), .Y(n_693) );
BUFx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2x1_ASAP7_75t_L g752 ( .A(n_664), .B(n_753), .Y(n_752) );
AND2x4_ASAP7_75t_L g681 ( .A(n_666), .B(n_682), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_676), .B2(n_680), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g696 ( .A(n_670), .B(n_697), .Y(n_696) );
OR2x6_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
NOR2x1_ASAP7_75t_SL g733 ( .A(n_672), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g797 ( .A(n_672), .Y(n_797) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g702 ( .A(n_673), .B(n_683), .Y(n_702) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVx2_ASAP7_75t_L g723 ( .A(n_678), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_678), .A2(n_723), .B1(n_781), .B2(n_782), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_679), .B(n_739), .Y(n_738) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g741 ( .A(n_683), .B(n_725), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B1(n_689), .B2(n_693), .C(n_699), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_687), .B(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g807 ( .A(n_688), .Y(n_807) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g745 ( .A(n_692), .Y(n_745) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_702), .B(n_712), .Y(n_711) );
AND2x4_ASAP7_75t_L g806 ( .A(n_702), .B(n_760), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_705), .B(n_771), .Y(n_704) );
NOR4xp25_ASAP7_75t_L g705 ( .A(n_706), .B(n_726), .C(n_743), .D(n_762), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_711), .B1(n_714), .B2(n_719), .C(n_721), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_708), .A2(n_730), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_710), .B(n_713), .Y(n_779) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_719), .A2(n_744), .B1(n_748), .B2(n_752), .C(n_754), .Y(n_743) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g726 ( .A1(n_727), .A2(n_731), .B(n_732), .Y(n_726) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g814 ( .A(n_729), .B(n_741), .Y(n_814) );
INVx2_ASAP7_75t_L g756 ( .A(n_731), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .B1(n_737), .B2(n_740), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g766 ( .A(n_739), .Y(n_766) );
INVx1_ASAP7_75t_L g786 ( .A(n_739), .Y(n_786) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVxp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI21xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B(n_757), .Y(n_754) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR3x2_ASAP7_75t_L g767 ( .A(n_760), .B(n_768), .C(n_769), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
NOR4xp75_ASAP7_75t_SL g771 ( .A(n_772), .B(n_791), .C(n_804), .D(n_809), .Y(n_771) );
NAND3x1_ASAP7_75t_L g772 ( .A(n_773), .B(n_777), .C(n_788), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_780), .B1(n_784), .B2(n_785), .Y(n_777) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NOR2x1_ASAP7_75t_SL g785 ( .A(n_786), .B(n_787), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_794), .B1(n_795), .B2(n_800), .Y(n_791) );
NAND3x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .C(n_798), .Y(n_795) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_807), .B(n_808), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
BUFx12f_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
AND2x6_ASAP7_75t_SL g819 ( .A(n_820), .B(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_821), .B(n_833), .Y(n_832) );
INVx3_ASAP7_75t_L g842 ( .A(n_821), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_821), .B(n_874), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_825), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NOR2x1_ASAP7_75t_L g835 ( .A(n_824), .B(n_826), .Y(n_835) );
AND2x6_ASAP7_75t_SL g847 ( .A(n_825), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx10_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NOR2xp67_ASAP7_75t_L g837 ( .A(n_838), .B(n_843), .Y(n_837) );
INVx4_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
CKINVDCx11_ASAP7_75t_R g840 ( .A(n_841), .Y(n_840) );
BUFx6f_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_842), .B(n_872), .Y(n_871) );
OAI21xp33_ASAP7_75t_L g868 ( .A1(n_843), .A2(n_869), .B(n_875), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_851), .B(n_855), .Y(n_843) );
BUFx3_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
BUFx12f_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx4_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
CKINVDCx8_ASAP7_75t_R g858 ( .A(n_847), .Y(n_858) );
INVx5_ASAP7_75t_L g867 ( .A(n_847), .Y(n_867) );
INVx3_ASAP7_75t_L g874 ( .A(n_847), .Y(n_874) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_859), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_861), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
CKINVDCx16_ASAP7_75t_R g863 ( .A(n_864), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_867), .Y(n_864) );
INVx2_ASAP7_75t_SL g873 ( .A(n_865), .Y(n_873) );
OR2x6_ASAP7_75t_L g869 ( .A(n_870), .B(n_874), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
OR2x4_ASAP7_75t_L g878 ( .A(n_872), .B(n_879), .Y(n_878) );
BUFx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g876 ( .A(n_877), .Y(n_876) );
INVx4_ASAP7_75t_SL g877 ( .A(n_878), .Y(n_877) );
endmodule