module fake_jpeg_1434_n_474 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_474);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_474;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_50),
.A2(n_30),
.B1(n_27),
.B2(n_44),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_51),
.B(n_54),
.Y(n_124)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_52),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_55),
.B(n_60),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_15),
.B(n_14),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_20),
.B(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_27),
.Y(n_150)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_24),
.A2(n_9),
.B(n_7),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_0),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_123),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_109),
.B(n_0),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_78),
.B1(n_23),
.B2(n_41),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_66),
.A2(n_19),
.B1(n_44),
.B2(n_30),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_87),
.B1(n_62),
.B2(n_86),
.Y(n_158)
);

BUFx4f_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_42),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_66),
.B(n_32),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_59),
.B(n_32),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_150),
.Y(n_193)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_53),
.B(n_38),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_152),
.C(n_139),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_188),
.C(n_132),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_105),
.A2(n_46),
.B1(n_41),
.B2(n_29),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_179),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_78),
.B1(n_44),
.B2(n_28),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_47),
.B1(n_80),
.B2(n_81),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_173),
.B(n_142),
.Y(n_210)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_48),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_177),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_112),
.A2(n_93),
.B1(n_58),
.B2(n_57),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_180),
.B1(n_191),
.B2(n_192),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_109),
.A2(n_56),
.B1(n_82),
.B2(n_75),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_61),
.B1(n_74),
.B2(n_73),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_124),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_196),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_70),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_68),
.B1(n_101),
.B2(n_143),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_124),
.A2(n_21),
.B1(n_46),
.B2(n_28),
.Y(n_192)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_135),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_226),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_177),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_151),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_233),
.C(n_158),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_194),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_147),
.B1(n_100),
.B2(n_153),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_215),
.A2(n_183),
.B1(n_108),
.B2(n_143),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_29),
.B(n_23),
.C(n_21),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_218),
.B(n_170),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_114),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_155),
.B(n_122),
.C(n_119),
.Y(n_233)
);

OAI32xp33_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_185),
.A3(n_173),
.B1(n_177),
.B2(n_172),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_238),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_241),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_248),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_163),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_162),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_240),
.B(n_258),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_204),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_214),
.A2(n_191),
.B1(n_197),
.B2(n_198),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_250),
.B1(n_254),
.B2(n_215),
.Y(n_272)
);

AOI32xp33_ASAP7_75t_L g243 ( 
.A1(n_199),
.A2(n_130),
.A3(n_106),
.B1(n_103),
.B2(n_190),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_249),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_158),
.B(n_166),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_253),
.B(n_246),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_245),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_217),
.A2(n_158),
.B(n_189),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_246),
.A2(n_261),
.B(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_201),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_100),
.B1(n_184),
.B2(n_153),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_225),
.B1(n_227),
.B2(n_229),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_195),
.B(n_134),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_120),
.B1(n_133),
.B2(n_168),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_257),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_204),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_202),
.B(n_175),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_206),
.B(n_168),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_262),
.Y(n_286)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_203),
.B(n_170),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_249),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_264),
.B(n_268),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_205),
.B1(n_199),
.B2(n_201),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_265),
.A2(n_253),
.B1(n_241),
.B2(n_250),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_233),
.C(n_220),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_259),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_240),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_220),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_258),
.C(n_237),
.Y(n_305)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_218),
.B1(n_200),
.B2(n_211),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_278),
.B1(n_287),
.B2(n_257),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_200),
.B1(n_211),
.B2(n_209),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_260),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_283),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_200),
.B1(n_222),
.B2(n_204),
.Y(n_287)
);

OAI22x1_ASAP7_75t_SL g288 ( 
.A1(n_254),
.A2(n_242),
.B1(n_261),
.B2(n_234),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_289),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_262),
.A2(n_101),
.B1(n_107),
.B2(n_227),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_237),
.A2(n_107),
.B1(n_229),
.B2(n_230),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_212),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_292),
.B(n_305),
.C(n_313),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_293),
.A2(n_306),
.B1(n_288),
.B2(n_289),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_284),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_298),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_243),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_297),
.A2(n_308),
.B(n_314),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_303),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_268),
.A2(n_235),
.B(n_238),
.Y(n_300)
);

OAI211xp5_ASAP7_75t_L g336 ( 
.A1(n_300),
.A2(n_309),
.B(n_320),
.C(n_280),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_269),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_304),
.A2(n_317),
.B1(n_318),
.B2(n_275),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_263),
.A2(n_250),
.B1(n_251),
.B2(n_239),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_263),
.B(n_277),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_277),
.A2(n_247),
.B1(n_252),
.B2(n_255),
.Y(n_309)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_264),
.B(n_245),
.Y(n_312)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_228),
.C(n_221),
.Y(n_313)
);

A2O1A1O1Ixp25_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_212),
.B(n_219),
.C(n_228),
.D(n_86),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_267),
.B(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_319),
.Y(n_324)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_275),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_267),
.B(n_222),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_222),
.B(n_219),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_323),
.A2(n_327),
.B1(n_329),
.B2(n_331),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_311),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_342),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_278),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_328),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_311),
.A2(n_273),
.B1(n_279),
.B2(n_281),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_294),
.A2(n_306),
.B1(n_293),
.B2(n_302),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_294),
.A2(n_272),
.B1(n_290),
.B2(n_274),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_346),
.B1(n_347),
.B2(n_310),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_266),
.C(n_271),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_339),
.C(n_345),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_303),
.B(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_335),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_315),
.Y(n_337)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_280),
.Y(n_338)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_266),
.C(n_286),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_281),
.Y(n_341)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_301),
.B(n_285),
.Y(n_342)
);

FAx1_ASAP7_75t_SL g343 ( 
.A(n_308),
.B(n_305),
.CI(n_296),
.CON(n_343),
.SN(n_343)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_348),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_285),
.C(n_186),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_302),
.A2(n_291),
.B1(n_213),
.B2(n_223),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_301),
.A2(n_304),
.B1(n_296),
.B2(n_320),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_291),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_335),
.B(n_297),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_351),
.B(n_325),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_309),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_361),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_314),
.Y(n_353)
);

XNOR2x1_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_346),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_318),
.Y(n_356)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_358),
.A2(n_372),
.B1(n_373),
.B2(n_321),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_317),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_307),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_364),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_291),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_331),
.Y(n_365)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_365),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_325),
.B(n_213),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_367),
.B(n_333),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_161),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_374),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_332),
.Y(n_369)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_7),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_338),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_327),
.A2(n_45),
.B1(n_37),
.B2(n_36),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_328),
.A2(n_45),
.B1(n_37),
.B2(n_36),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_45),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_375),
.A2(n_344),
.B1(n_349),
.B2(n_342),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_377),
.A2(n_383),
.B1(n_384),
.B2(n_392),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_345),
.C(n_340),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_396),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_394),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_362),
.A2(n_344),
.B1(n_349),
.B2(n_347),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_359),
.A2(n_336),
.B(n_337),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_385),
.A2(n_360),
.B(n_373),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_324),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_391),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_321),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_355),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_343),
.Y(n_389)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_389),
.Y(n_401)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_324),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_371),
.A2(n_333),
.B1(n_341),
.B2(n_348),
.Y(n_392)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_343),
.C(n_45),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_45),
.C(n_37),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_353),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_377),
.A2(n_383),
.B1(n_358),
.B2(n_380),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_399),
.A2(n_400),
.B1(n_416),
.B2(n_31),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_393),
.A2(n_360),
.B1(n_366),
.B2(n_350),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_387),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_403),
.Y(n_417)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g418 ( 
.A1(n_404),
.A2(n_379),
.B(n_396),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_409),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_394),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_410),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_368),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_381),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_351),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_0),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_413),
.A2(n_18),
.B(n_1),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_386),
.A2(n_372),
.B1(n_374),
.B2(n_45),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_418),
.A2(n_431),
.B1(n_405),
.B2(n_413),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_378),
.Y(n_419)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_378),
.C(n_391),
.Y(n_421)
);

FAx1_ASAP7_75t_SL g435 ( 
.A(n_421),
.B(n_400),
.CI(n_407),
.CON(n_435),
.SN(n_435)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_401),
.A2(n_397),
.B(n_386),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_422),
.A2(n_2),
.B(n_3),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_403),
.A2(n_36),
.B1(n_31),
.B2(n_18),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_423),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_412),
.B(n_31),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_426),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_406),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_432),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_429),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_414),
.B(n_1),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_430),
.B(n_6),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_411),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_2),
.C(n_3),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_408),
.C(n_409),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_2),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_399),
.C(n_402),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_435),
.Y(n_456)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_437),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_416),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_438),
.B(n_446),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_5),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_440),
.A2(n_431),
.B(n_5),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_441),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_3),
.C(n_4),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_SL g453 ( 
.A(n_443),
.B(n_432),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_4),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_SL g449 ( 
.A1(n_445),
.A2(n_424),
.B(n_426),
.C(n_428),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_449),
.A2(n_455),
.B1(n_444),
.B2(n_442),
.Y(n_462)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_452),
.Y(n_458)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_453),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_434),
.A2(n_420),
.B(n_429),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_454),
.A2(n_443),
.B(n_436),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_SL g455 ( 
.A1(n_435),
.A2(n_427),
.B(n_423),
.C(n_421),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_457),
.B(n_447),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_448),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_459),
.B(n_461),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_460),
.B(n_464),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_462),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_456),
.A2(n_444),
.B(n_442),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_463),
.B(n_451),
.C(n_447),
.Y(n_466)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_466),
.Y(n_469)
);

AOI321xp33_ASAP7_75t_L g470 ( 
.A1(n_468),
.A2(n_459),
.A3(n_455),
.B1(n_458),
.B2(n_6),
.C(n_5),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_465),
.C(n_467),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_469),
.C(n_5),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_472),
.A2(n_5),
.B(n_6),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_473),
.B(n_6),
.Y(n_474)
);


endmodule