module fake_netlist_6_299_n_2079 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2079);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2079;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_1909;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_1970;
wire n_608;
wire n_630;
wire n_2059;
wire n_2073;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_1492;
wire n_987;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_2069;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_1092;
wire n_1060;
wire n_1951;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1832;
wire n_1645;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_652;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_2015;
wire n_1148;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_525),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_338),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_453),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_208),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_451),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_290),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_241),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_541),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_227),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_65),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_51),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_458),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_301),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_180),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_313),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_539),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_45),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_496),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_53),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_518),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_54),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_484),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_282),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_358),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_131),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_444),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_269),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_531),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_263),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_110),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_176),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_413),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_299),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_446),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_526),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_280),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_461),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_46),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_305),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_438),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_240),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_542),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_212),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_449),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_363),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_379),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_540),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_216),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_433),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_209),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_536),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_474),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_177),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_376),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_138),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_83),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_43),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_468),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_527),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_355),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_409),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_544),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_86),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_516),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_532),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_443),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_161),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_524),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_560),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_78),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_530),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_141),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_64),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_324),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_546),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_100),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_510),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_417),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_537),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_162),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_11),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_71),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_283),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_37),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_74),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_96),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_133),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_250),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_68),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_523),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_538),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_14),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_428),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_146),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_559),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_418),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_29),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_292),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_79),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_50),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_107),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_529),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_271),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_251),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_274),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_45),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_190),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_382),
.Y(n_672)
);

CKINVDCx16_ASAP7_75t_R g673 ( 
.A(n_151),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_316),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_535),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_383),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_320),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_462),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_400),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_32),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_351),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_70),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_362),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_59),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_181),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_148),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_92),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_235),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_256),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_163),
.Y(n_690)
);

CKINVDCx16_ASAP7_75t_R g691 ( 
.A(n_106),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_488),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_492),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_501),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_248),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_26),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_513),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_534),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_15),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_463),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_491),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_168),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_81),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_270),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_533),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_543),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_196),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_310),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_165),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_450),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_197),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_68),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_426),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_86),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_476),
.Y(n_715)
);

BUFx5_ASAP7_75t_L g716 ( 
.A(n_276),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_478),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_325),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_304),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_74),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_550),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_528),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_226),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_142),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_170),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_503),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_13),
.Y(n_727)
);

BUFx5_ASAP7_75t_L g728 ( 
.A(n_31),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_113),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_422),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_108),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_416),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_87),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_545),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_73),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_50),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_175),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_63),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_116),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_728),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_728),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_728),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_728),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_672),
.Y(n_744)
);

XOR2xp5_ASAP7_75t_L g745 ( 
.A(n_691),
.B(n_0),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_728),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_636),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_565),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_567),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_671),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_568),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_649),
.Y(n_752)
);

INVxp67_ASAP7_75t_SL g753 ( 
.A(n_582),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_634),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_637),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_646),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_650),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_574),
.B(n_0),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_578),
.Y(n_759)
);

INVxp33_ASAP7_75t_SL g760 ( 
.A(n_575),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_587),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_588),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_589),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_569),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_596),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_716),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_591),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_716),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_591),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_599),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_605),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_591),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_581),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_665),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_598),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_570),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_611),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_716),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_612),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_580),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_566),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_586),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_614),
.Y(n_783)
);

CKINVDCx14_ASAP7_75t_R g784 ( 
.A(n_580),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_583),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_716),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_619),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_571),
.Y(n_788)
);

INVxp33_ASAP7_75t_L g789 ( 
.A(n_625),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_576),
.Y(n_790)
);

INVxp33_ASAP7_75t_L g791 ( 
.A(n_626),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_577),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_632),
.Y(n_793)
);

CKINVDCx14_ASAP7_75t_R g794 ( 
.A(n_629),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_644),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_647),
.Y(n_796)
);

INVxp33_ASAP7_75t_L g797 ( 
.A(n_651),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_654),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_606),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_716),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_655),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_659),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_674),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_629),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_686),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_689),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_585),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_690),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_673),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_652),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_693),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_602),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_704),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_694),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_620),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_700),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_572),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_701),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_594),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_707),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_579),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_708),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_621),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_709),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_710),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_610),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_718),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_723),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_660),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_729),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_730),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_739),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_713),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_584),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_573),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_590),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_666),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_592),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_601),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_598),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_753),
.B(n_652),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_782),
.B(n_633),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_799),
.B(n_679),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_769),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_769),
.Y(n_845)
);

OA21x2_ASAP7_75t_L g846 ( 
.A1(n_740),
.A2(n_617),
.B(n_607),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_808),
.B(n_600),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_769),
.Y(n_848)
);

CKINVDCx6p67_ASAP7_75t_R g849 ( 
.A(n_780),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_748),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_804),
.B(n_737),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_775),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_760),
.B(n_635),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_749),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_774),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_750),
.A2(n_640),
.B1(n_645),
.B2(n_627),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_751),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_741),
.A2(n_677),
.B(n_618),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_764),
.B(n_698),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_775),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_775),
.Y(n_861)
);

BUFx12f_ASAP7_75t_L g862 ( 
.A(n_776),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_840),
.Y(n_863)
);

CKINVDCx11_ASAP7_75t_R g864 ( 
.A(n_781),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_754),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_747),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_813),
.Y(n_867)
);

OA21x2_ASAP7_75t_L g868 ( 
.A1(n_742),
.A2(n_706),
.B(n_724),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_809),
.A2(n_692),
.B1(n_717),
.B2(n_685),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_810),
.B(n_725),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_774),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_767),
.B(n_772),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_743),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_788),
.B(n_732),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_773),
.Y(n_875)
);

CKINVDCx16_ASAP7_75t_R g876 ( 
.A(n_784),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_833),
.Y(n_877)
);

OAI21x1_ASAP7_75t_L g878 ( 
.A1(n_766),
.A2(n_595),
.B(n_593),
.Y(n_878)
);

AND2x6_ASAP7_75t_L g879 ( 
.A(n_746),
.B(n_598),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_755),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_756),
.Y(n_881)
);

INVx6_ASAP7_75t_L g882 ( 
.A(n_785),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_757),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_767),
.B(n_643),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_835),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_SL g886 ( 
.A1(n_745),
.A2(n_699),
.B1(n_696),
.B2(n_653),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_838),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_L g888 ( 
.A(n_807),
.B(n_648),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_790),
.B(n_658),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_772),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_839),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_768),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_SL g893 ( 
.A1(n_794),
.A2(n_661),
.B1(n_663),
.B2(n_656),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_778),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_744),
.A2(n_726),
.B1(n_670),
.B2(n_680),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_786),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_792),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_752),
.A2(n_682),
.B1(n_684),
.B2(n_664),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_800),
.Y(n_899)
);

BUFx8_ASAP7_75t_SL g900 ( 
.A(n_817),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_821),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_834),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_752),
.A2(n_703),
.B1(n_712),
.B2(n_687),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_759),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_761),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_762),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_785),
.B(n_812),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_763),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_765),
.A2(n_603),
.B(n_597),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_823),
.Y(n_910)
);

BUFx8_ASAP7_75t_SL g911 ( 
.A(n_837),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_770),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_771),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_812),
.A2(n_720),
.B1(n_727),
.B2(n_714),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_836),
.B(n_702),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_777),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_832),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_815),
.B(n_688),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_815),
.B(n_705),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_779),
.B(n_711),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_758),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_831),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_783),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_819),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_787),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_793),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_855),
.B(n_789),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_867),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_894),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_863),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_863),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_844),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_925),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_845),
.Y(n_934)
);

XOR2xp5_ASAP7_75t_L g935 ( 
.A(n_886),
.B(n_826),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_871),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_845),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_882),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_900),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_848),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_925),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_907),
.B(n_791),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_926),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_926),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_894),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_852),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_860),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_876),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_848),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_896),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_896),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_861),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_872),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_912),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_921),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_861),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_872),
.Y(n_957)
);

AND2x6_ASAP7_75t_L g958 ( 
.A(n_918),
.B(n_615),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_884),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_865),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_884),
.B(n_797),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_906),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_912),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_916),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_916),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_865),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_877),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_873),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_908),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_917),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_922),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_890),
.B(n_795),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_923),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_885),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_846),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_875),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_889),
.B(n_796),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_887),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_891),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_846),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_858),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_880),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_890),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_858),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_881),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_910),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_899),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_882),
.B(n_811),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_899),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_904),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_841),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_905),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_913),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_868),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_883),
.Y(n_995)
);

AND2x6_ASAP7_75t_L g996 ( 
.A(n_847),
.B(n_615),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_868),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_878),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_859),
.B(n_798),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_842),
.B(n_801),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_853),
.B(n_818),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_892),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_892),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_892),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_920),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_851),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_851),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_870),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_879),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_870),
.Y(n_1010)
);

INVx6_ASAP7_75t_L g1011 ( 
.A(n_866),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_842),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_843),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_879),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_847),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_843),
.B(n_802),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_879),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_919),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_909),
.Y(n_1019)
);

CKINVDCx16_ASAP7_75t_R g1020 ( 
.A(n_948),
.Y(n_1020)
);

AND3x2_ASAP7_75t_L g1021 ( 
.A(n_936),
.B(n_924),
.C(n_805),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_960),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_960),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_1018),
.B(n_850),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_959),
.B(n_895),
.Y(n_1025)
);

INVx5_ASAP7_75t_L g1026 ( 
.A(n_1011),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_L g1027 ( 
.A(n_1011),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_987),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_960),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_966),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_957),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_966),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_957),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_934),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_936),
.B(n_924),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_1005),
.B(n_897),
.Y(n_1036)
);

OR2x6_ASAP7_75t_L g1037 ( 
.A(n_927),
.B(n_862),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_L g1038 ( 
.A(n_976),
.B(n_893),
.C(n_856),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_957),
.B(n_854),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_966),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_953),
.B(n_874),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_953),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_967),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_954),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_962),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_963),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_964),
.Y(n_1047)
);

INVx5_ASAP7_75t_L g1048 ( 
.A(n_934),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_997),
.B(n_902),
.Y(n_1049)
);

INVxp67_ASAP7_75t_SL g1050 ( 
.A(n_975),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_965),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_977),
.B(n_915),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_959),
.B(n_854),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_983),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_961),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_986),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_942),
.B(n_876),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1012),
.B(n_857),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_971),
.Y(n_1059)
);

AND3x2_ASAP7_75t_L g1060 ( 
.A(n_976),
.B(n_806),
.C(n_803),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_938),
.B(n_866),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_982),
.Y(n_1062)
);

BUFx8_ASAP7_75t_SL g1063 ( 
.A(n_939),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_999),
.B(n_857),
.Y(n_1064)
);

BUFx4f_ASAP7_75t_L g1065 ( 
.A(n_967),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_989),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_1013),
.B(n_866),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_L g1068 ( 
.A(n_975),
.B(n_980),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_934),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_974),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1001),
.B(n_901),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_978),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_937),
.Y(n_1073)
);

AND3x2_ASAP7_75t_L g1074 ( 
.A(n_991),
.B(n_816),
.C(n_814),
.Y(n_1074)
);

OAI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1015),
.A2(n_869),
.B1(n_829),
.B2(n_849),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_979),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_967),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_991),
.B(n_914),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_988),
.B(n_604),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_973),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1006),
.B(n_888),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_985),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_928),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_975),
.B(n_820),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_980),
.B(n_822),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_972),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_937),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_972),
.A2(n_825),
.B1(n_827),
.B2(n_824),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1007),
.Y(n_1089)
);

NOR2x1p5_ASAP7_75t_L g1090 ( 
.A(n_1000),
.B(n_731),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_937),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_980),
.B(n_828),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_935),
.Y(n_1093)
);

INVx4_ASAP7_75t_L g1094 ( 
.A(n_940),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_955),
.B(n_898),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_969),
.Y(n_1096)
);

BUFx8_ASAP7_75t_SL g1097 ( 
.A(n_992),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_969),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_970),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1016),
.B(n_903),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_970),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_SL g1102 ( 
.A(n_1009),
.B(n_733),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_940),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_981),
.B(n_830),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1008),
.Y(n_1105)
);

BUFx8_ASAP7_75t_SL g1106 ( 
.A(n_995),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1010),
.B(n_911),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_935),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_929),
.Y(n_1109)
);

CKINVDCx14_ASAP7_75t_R g1110 ( 
.A(n_958),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_940),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_990),
.B(n_719),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_932),
.Y(n_1113)
);

INVxp33_ASAP7_75t_L g1114 ( 
.A(n_930),
.Y(n_1114)
);

AO22x1_ASAP7_75t_L g1115 ( 
.A1(n_996),
.A2(n_736),
.B1(n_738),
.B2(n_735),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_931),
.B(n_721),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1009),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_1009),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1036),
.B(n_993),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1042),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1052),
.B(n_981),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_1056),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1100),
.A2(n_996),
.B1(n_998),
.B2(n_958),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1024),
.B(n_864),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_L g1125 ( 
.A(n_1071),
.B(n_968),
.C(n_941),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_1056),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_1077),
.B(n_933),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1033),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1089),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1055),
.B(n_943),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1064),
.B(n_929),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1025),
.B(n_949),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1041),
.B(n_981),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_1034),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_1068),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1066),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1025),
.B(n_952),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1045),
.Y(n_1138)
);

AND2x6_ASAP7_75t_L g1139 ( 
.A(n_1081),
.B(n_1019),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_L g1140 ( 
.A(n_1078),
.B(n_944),
.C(n_951),
.Y(n_1140)
);

NAND2xp33_ASAP7_75t_L g1141 ( 
.A(n_1049),
.B(n_984),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1062),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1050),
.B(n_1054),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_1088),
.A2(n_956),
.B(n_950),
.Y(n_1144)
);

BUFx8_ASAP7_75t_L g1145 ( 
.A(n_1057),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_1117),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1084),
.A2(n_1017),
.B(n_946),
.C(n_947),
.Y(n_1147)
);

INVx8_ASAP7_75t_L g1148 ( 
.A(n_1026),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1072),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1105),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1044),
.A2(n_996),
.B1(n_998),
.B2(n_958),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1085),
.B(n_984),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_1074),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1046),
.Y(n_1154)
);

NAND2x1_ASAP7_75t_L g1155 ( 
.A(n_1118),
.B(n_984),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1047),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1051),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1038),
.B(n_950),
.C(n_945),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1092),
.B(n_994),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1104),
.B(n_1058),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1065),
.B(n_945),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1031),
.B(n_994),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1061),
.B(n_1014),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1053),
.B(n_1014),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1086),
.A2(n_1028),
.B(n_1082),
.C(n_1080),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1117),
.B(n_994),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1114),
.B(n_998),
.Y(n_1167)
);

INVxp67_ASAP7_75t_L g1168 ( 
.A(n_1035),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1109),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1053),
.B(n_1014),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1096),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1059),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1070),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1049),
.B(n_1019),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1049),
.B(n_1004),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_1034),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1076),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1113),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1035),
.B(n_688),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1075),
.B(n_1002),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1098),
.B(n_1003),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1020),
.B(n_1039),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1043),
.B(n_608),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1099),
.B(n_609),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1101),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1083),
.B(n_109),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1090),
.A2(n_615),
.B1(n_715),
.B2(n_616),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1022),
.B(n_613),
.Y(n_1188)
);

AO22x2_ASAP7_75t_L g1189 ( 
.A1(n_1067),
.A2(n_9),
.B1(n_17),
.B2(n_1),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1023),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1029),
.B(n_622),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1095),
.A2(n_715),
.B1(n_624),
.B2(n_628),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1027),
.B(n_623),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1095),
.A2(n_631),
.B1(n_638),
.B2(n_630),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1030),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1079),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1132),
.B(n_1107),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1138),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1126),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1122),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1154),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1152),
.A2(n_1159),
.B(n_1133),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1156),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1148),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1163),
.B(n_1091),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1124),
.B(n_1108),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1157),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1137),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1129),
.B(n_1037),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1164),
.B(n_1032),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1196),
.A2(n_1112),
.B1(n_1116),
.B2(n_1110),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1150),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1142),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1146),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1121),
.A2(n_1040),
.B1(n_1111),
.B2(n_1094),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_1169),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1160),
.B(n_1115),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1135),
.B(n_1069),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1148),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1146),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1149),
.Y(n_1221)
);

NAND2x1_ASAP7_75t_L g1222 ( 
.A(n_1139),
.B(n_1069),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1170),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1119),
.B(n_1093),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1182),
.B(n_1021),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1172),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1136),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1143),
.B(n_1073),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1173),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1165),
.A2(n_1102),
.B(n_1073),
.C(n_1087),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1177),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1145),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1186),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1186),
.B(n_1026),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1167),
.B(n_1087),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1178),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1125),
.B(n_1103),
.Y(n_1237)
);

O2A1O1Ixp5_ASAP7_75t_L g1238 ( 
.A1(n_1131),
.A2(n_1060),
.B(n_1103),
.C(n_641),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1120),
.B(n_1048),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1192),
.B(n_1048),
.Y(n_1240)
);

BUFx4f_ASAP7_75t_L g1241 ( 
.A(n_1153),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1128),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1130),
.B(n_639),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1185),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1171),
.B(n_642),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1171),
.B(n_657),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1181),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1162),
.B(n_662),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1134),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1145),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1127),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1123),
.B(n_667),
.Y(n_1252)
);

NOR3xp33_ASAP7_75t_SL g1253 ( 
.A(n_1158),
.B(n_669),
.C(n_668),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1190),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_SL g1255 ( 
.A(n_1168),
.B(n_1063),
.Y(n_1255)
);

NOR3xp33_ASAP7_75t_SL g1256 ( 
.A(n_1194),
.B(n_676),
.C(n_675),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1195),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1144),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1180),
.B(n_1127),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1166),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1179),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1139),
.B(n_678),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1176),
.B(n_1037),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_SL g1264 ( 
.A(n_1187),
.B(n_683),
.C(n_681),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1175),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1139),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1140),
.B(n_1097),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1141),
.A2(n_715),
.B(n_697),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1161),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1147),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_L g1271 ( 
.A(n_1193),
.B(n_695),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1188),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1191),
.B(n_1151),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1232),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1204),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1229),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1199),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1201),
.Y(n_1278)
);

INVx5_ASAP7_75t_L g1279 ( 
.A(n_1214),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1203),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1222),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1207),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1212),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1200),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1263),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1226),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1224),
.A2(n_1183),
.B1(n_1184),
.B2(n_1139),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1231),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1263),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1197),
.B(n_1174),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1208),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1223),
.B(n_1189),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1236),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1210),
.B(n_1155),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1272),
.B(n_1106),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1247),
.B(n_1189),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1223),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1227),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1223),
.B(n_722),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1217),
.A2(n_734),
.B(n_3),
.C(n_1),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1265),
.B(n_2),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1210),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1259),
.A2(n_1273),
.B(n_1258),
.C(n_1202),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1233),
.B(n_2),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1205),
.Y(n_1305)
);

INVx4_ASAP7_75t_L g1306 ( 
.A(n_1214),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1233),
.B(n_3),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_1256),
.B(n_4),
.C(n_5),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1233),
.B(n_4),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1214),
.B(n_5),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1205),
.B(n_6),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1228),
.B(n_6),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1198),
.Y(n_1313)
);

AND3x1_ASAP7_75t_SL g1314 ( 
.A(n_1244),
.B(n_7),
.C(n_8),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1218),
.B(n_7),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1219),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1206),
.B(n_8),
.Y(n_1317)
);

INVx6_ASAP7_75t_L g1318 ( 
.A(n_1250),
.Y(n_1318)
);

XNOR2xp5_ASAP7_75t_L g1319 ( 
.A(n_1211),
.B(n_111),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1213),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1251),
.B(n_9),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1221),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1266),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1269),
.B(n_10),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1242),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1254),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1234),
.B(n_112),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1257),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1260),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1264),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1239),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1220),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1216),
.B(n_12),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1237),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1235),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1245),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_R g1337 ( 
.A(n_1255),
.B(n_114),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1248),
.B(n_13),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1225),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1241),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1246),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1209),
.B(n_16),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1243),
.B(n_17),
.Y(n_1343)
);

INVx4_ASAP7_75t_L g1344 ( 
.A(n_1261),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1270),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1249),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1240),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1230),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_R g1349 ( 
.A(n_1267),
.B(n_115),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1238),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1252),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1278),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1317),
.A2(n_1253),
.B(n_1271),
.C(n_1268),
.Y(n_1353)
);

A2O1A1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1338),
.A2(n_1262),
.B(n_1215),
.C(n_20),
.Y(n_1354)
);

INVx8_ASAP7_75t_L g1355 ( 
.A(n_1279),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1340),
.Y(n_1356)
);

AOI211x1_ASAP7_75t_L g1357 ( 
.A1(n_1296),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1303),
.A2(n_118),
.B(n_117),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1336),
.B(n_18),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1348),
.A2(n_120),
.B(n_119),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1341),
.A2(n_564),
.B(n_122),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1292),
.B(n_19),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1350),
.A2(n_123),
.B(n_121),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1351),
.B(n_21),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1280),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1345),
.A2(n_125),
.B(n_124),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1281),
.A2(n_127),
.B(n_126),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1300),
.A2(n_129),
.A3(n_130),
.B(n_128),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1331),
.B(n_21),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1305),
.B(n_22),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1347),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1290),
.A2(n_23),
.B(n_24),
.Y(n_1372)
);

CKINVDCx11_ASAP7_75t_R g1373 ( 
.A(n_1340),
.Y(n_1373)
);

NOR2x1_ASAP7_75t_SL g1374 ( 
.A(n_1279),
.B(n_132),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1282),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1291),
.B(n_25),
.Y(n_1376)
);

A2O1A1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1287),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1283),
.Y(n_1378)
);

BUFx12f_ASAP7_75t_L g1379 ( 
.A(n_1340),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1281),
.A2(n_1323),
.B(n_1334),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1312),
.A2(n_27),
.B(n_28),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1284),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1318),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1343),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1323),
.A2(n_135),
.B(n_134),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1302),
.B(n_30),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1313),
.A2(n_137),
.B(n_136),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1279),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1301),
.A2(n_140),
.B(n_139),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1277),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1286),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1276),
.B(n_31),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1313),
.A2(n_144),
.B(n_143),
.Y(n_1393)
);

NAND3xp33_ASAP7_75t_L g1394 ( 
.A(n_1330),
.B(n_32),
.C(n_33),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1315),
.A2(n_147),
.B(n_145),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1274),
.Y(n_1396)
);

AO21x1_ASAP7_75t_L g1397 ( 
.A1(n_1335),
.A2(n_33),
.B(n_34),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1297),
.B(n_34),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1295),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1327),
.B(n_35),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1288),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1326),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1306),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1299),
.B(n_36),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1318),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1298),
.B(n_38),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1325),
.A2(n_150),
.B(n_149),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1332),
.A2(n_563),
.B(n_153),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1319),
.B(n_1327),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1329),
.A2(n_154),
.B(n_152),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1293),
.A2(n_156),
.B(n_155),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1342),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1320),
.A2(n_158),
.B(n_157),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1308),
.A2(n_39),
.B(n_40),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1332),
.A2(n_160),
.B(n_159),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1321),
.A2(n_41),
.B(n_42),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_SL g1417 ( 
.A1(n_1304),
.A2(n_41),
.B(n_42),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1322),
.A2(n_1328),
.B(n_1309),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1306),
.B(n_164),
.Y(n_1419)
);

AOI211x1_ASAP7_75t_L g1420 ( 
.A1(n_1324),
.A2(n_46),
.B(n_43),
.C(n_44),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1285),
.B(n_44),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1289),
.B(n_47),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1349),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1339),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1310),
.A2(n_562),
.B(n_167),
.Y(n_1425)
);

OAI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1333),
.A2(n_48),
.B(n_49),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1311),
.B(n_1307),
.Y(n_1427)
);

BUFx5_ASAP7_75t_L g1428 ( 
.A(n_1294),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1294),
.A2(n_561),
.B(n_169),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1346),
.B(n_51),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1316),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1344),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1432)
);

AOI21xp33_ASAP7_75t_L g1433 ( 
.A1(n_1344),
.A2(n_52),
.B(n_55),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1314),
.A2(n_171),
.B(n_166),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1337),
.A2(n_173),
.B(n_172),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1275),
.B(n_55),
.Y(n_1436)
);

INVx4_ASAP7_75t_L g1437 ( 
.A(n_1279),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1348),
.A2(n_178),
.B(n_174),
.Y(n_1438)
);

O2A1O1Ixp5_ASAP7_75t_L g1439 ( 
.A1(n_1350),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1351),
.B(n_56),
.Y(n_1440)
);

AOI211x1_ASAP7_75t_L g1441 ( 
.A1(n_1296),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1348),
.A2(n_182),
.B(n_179),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1285),
.B(n_183),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1303),
.A2(n_558),
.B(n_185),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1351),
.B(n_184),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1405),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1427),
.B(n_60),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1409),
.B(n_186),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1362),
.B(n_187),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1352),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1363),
.A2(n_189),
.B(n_188),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_SL g1452 ( 
.A(n_1437),
.B(n_1388),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1390),
.B(n_191),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1396),
.Y(n_1454)
);

BUFx4_ASAP7_75t_SL g1455 ( 
.A(n_1423),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_SL g1456 ( 
.A(n_1388),
.B(n_192),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1373),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1402),
.B(n_193),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1365),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1382),
.B(n_194),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1358),
.A2(n_198),
.B(n_195),
.Y(n_1461)
);

NAND2xp33_ASAP7_75t_L g1462 ( 
.A(n_1426),
.B(n_1424),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1356),
.Y(n_1463)
);

OR2x6_ASAP7_75t_SL g1464 ( 
.A(n_1399),
.B(n_60),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1375),
.B(n_61),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1378),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1391),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1356),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1445),
.B(n_1400),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1359),
.B(n_61),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1404),
.B(n_199),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1355),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1401),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1379),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1369),
.B(n_1398),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1418),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1355),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1406),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1394),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1416),
.A2(n_66),
.B1(n_62),
.B2(n_65),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1431),
.B(n_200),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1392),
.Y(n_1482)
);

INVx5_ASAP7_75t_L g1483 ( 
.A(n_1383),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1372),
.B(n_201),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1444),
.A2(n_203),
.B(n_202),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1368),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1364),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1443),
.B(n_204),
.Y(n_1488)
);

NAND2x1p5_ASAP7_75t_L g1489 ( 
.A(n_1403),
.B(n_205),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1428),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1397),
.Y(n_1491)
);

NAND2x1p5_ASAP7_75t_L g1492 ( 
.A(n_1435),
.B(n_206),
.Y(n_1492)
);

AOI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1380),
.A2(n_210),
.B(n_207),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1377),
.B(n_66),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1353),
.A2(n_213),
.B(n_211),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1370),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1428),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1354),
.A2(n_215),
.B(n_214),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1414),
.B(n_67),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1428),
.Y(n_1500)
);

BUFx10_ASAP7_75t_L g1501 ( 
.A(n_1440),
.Y(n_1501)
);

AOI21xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1436),
.A2(n_67),
.B(n_69),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1428),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_SL g1504 ( 
.A1(n_1395),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1420),
.B(n_1357),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1421),
.B(n_217),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_SL g1507 ( 
.A1(n_1361),
.A2(n_75),
.B(n_72),
.C(n_73),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1386),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1384),
.A2(n_76),
.B1(n_72),
.B2(n_75),
.C(n_77),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1430),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1366),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1368),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1422),
.B(n_218),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1376),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1441),
.B(n_1412),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1389),
.A2(n_220),
.B(n_219),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1419),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_SL g1518 ( 
.A1(n_1374),
.A2(n_222),
.B(n_221),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1408),
.A2(n_224),
.B(n_223),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1434),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1432),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1425),
.B(n_225),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1433),
.B(n_228),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1371),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1417),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1439),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1385),
.B(n_229),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1387),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1410),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1381),
.B(n_1429),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1367),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1415),
.B(n_79),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1393),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1411),
.A2(n_231),
.B(n_230),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1407),
.A2(n_233),
.B(n_232),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1360),
.A2(n_236),
.B(n_234),
.Y(n_1536)
);

BUFx8_ASAP7_75t_L g1537 ( 
.A(n_1413),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1438),
.Y(n_1538)
);

CKINVDCx16_ASAP7_75t_R g1539 ( 
.A(n_1442),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1378),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1390),
.B(n_237),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1427),
.B(n_80),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1521),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1461),
.A2(n_239),
.B(n_238),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1485),
.A2(n_243),
.B(n_242),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1478),
.B(n_82),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1483),
.B(n_83),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1459),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1467),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1497),
.B(n_244),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1496),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1462),
.A2(n_87),
.B(n_84),
.C(n_85),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1456),
.A2(n_246),
.B(n_245),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1507),
.A2(n_88),
.B(n_84),
.C(n_85),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1473),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1495),
.A2(n_249),
.B(n_247),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1466),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1482),
.B(n_88),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1540),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1450),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1491),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1475),
.B(n_89),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1498),
.A2(n_253),
.B(n_252),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1517),
.B(n_254),
.Y(n_1564)
);

O2A1O1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1499),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1504),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1476),
.Y(n_1567)
);

AND2x6_ASAP7_75t_L g1568 ( 
.A(n_1525),
.B(n_1527),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1503),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1514),
.B(n_93),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1510),
.B(n_93),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1508),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1486),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1446),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1519),
.A2(n_257),
.B(n_255),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1449),
.B(n_94),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1487),
.B(n_94),
.Y(n_1577)
);

O2A1O1Ixp5_ASAP7_75t_L g1578 ( 
.A1(n_1516),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1486),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1469),
.A2(n_1480),
.B(n_1509),
.C(n_1479),
.Y(n_1580)
);

INVx4_ASAP7_75t_L g1581 ( 
.A(n_1483),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1490),
.B(n_258),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1512),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1453),
.B(n_95),
.Y(n_1584)
);

NOR2xp67_ASAP7_75t_L g1585 ( 
.A(n_1472),
.B(n_1477),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1465),
.B(n_97),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1541),
.B(n_98),
.Y(n_1587)
);

O2A1O1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1502),
.A2(n_1494),
.B(n_1532),
.C(n_1530),
.Y(n_1588)
);

BUFx10_ASAP7_75t_L g1589 ( 
.A(n_1457),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1463),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1447),
.B(n_98),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1512),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1526),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1471),
.B(n_99),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1448),
.B(n_1454),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1533),
.A2(n_99),
.B(n_100),
.Y(n_1596)
);

NOR2xp67_ASAP7_75t_L g1597 ( 
.A(n_1500),
.B(n_101),
.Y(n_1597)
);

A2O1A1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1494),
.A2(n_1523),
.B(n_1524),
.C(n_1484),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1474),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1542),
.B(n_101),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1515),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1464),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1534),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1511),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1529),
.Y(n_1605)
);

NOR2xp67_ASAP7_75t_L g1606 ( 
.A(n_1470),
.B(n_105),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1501),
.B(n_108),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1489),
.A2(n_259),
.B(n_260),
.Y(n_1608)
);

AOI21x1_ASAP7_75t_SL g1609 ( 
.A1(n_1505),
.A2(n_261),
.B(n_262),
.Y(n_1609)
);

A2O1A1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1535),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1460),
.B(n_267),
.Y(n_1611)
);

NAND2x1p5_ASAP7_75t_L g1612 ( 
.A(n_1488),
.B(n_268),
.Y(n_1612)
);

BUFx12f_ASAP7_75t_L g1613 ( 
.A(n_1474),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_R g1614 ( 
.A(n_1463),
.B(n_272),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1536),
.A2(n_273),
.B(n_275),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1481),
.B(n_1458),
.Y(n_1616)
);

O2A1O1Ixp5_ASAP7_75t_L g1617 ( 
.A1(n_1520),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1452),
.B(n_281),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1529),
.Y(n_1619)
);

AOI221x1_ASAP7_75t_SL g1620 ( 
.A1(n_1506),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.C(n_287),
.Y(n_1620)
);

CKINVDCx6p67_ASAP7_75t_R g1621 ( 
.A(n_1468),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_SL g1622 ( 
.A(n_1513),
.B(n_288),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1468),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1528),
.B(n_289),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1539),
.B(n_1492),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1531),
.Y(n_1626)
);

A2O1A1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1522),
.A2(n_1451),
.B(n_1538),
.C(n_1531),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_L g1628 ( 
.A(n_1518),
.B(n_291),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1493),
.B(n_293),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1455),
.B(n_557),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1537),
.A2(n_294),
.B(n_295),
.Y(n_1631)
);

A2O1A1Ixp33_ASAP7_75t_SL g1632 ( 
.A1(n_1491),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1475),
.B(n_556),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1497),
.B(n_300),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1461),
.A2(n_302),
.B(n_303),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1521),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1475),
.B(n_309),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1475),
.B(n_555),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1478),
.B(n_311),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1497),
.B(n_312),
.Y(n_1640)
);

AOI221x1_ASAP7_75t_L g1641 ( 
.A1(n_1502),
.A2(n_314),
.B1(n_315),
.B2(n_317),
.C(n_318),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1446),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1496),
.B(n_319),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1467),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1461),
.A2(n_321),
.B(n_322),
.Y(n_1645)
);

A2O1A1Ixp33_ASAP7_75t_SL g1646 ( 
.A1(n_1491),
.A2(n_327),
.B(n_323),
.C(n_326),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1466),
.B(n_328),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1496),
.B(n_329),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1475),
.B(n_330),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1459),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1467),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1475),
.B(n_554),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1466),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_L g1654 ( 
.A(n_1462),
.B(n_331),
.C(n_332),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1478),
.B(n_333),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1478),
.B(n_334),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1593),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1551),
.B(n_335),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1653),
.B(n_1572),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1569),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1549),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1581),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1557),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1555),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1609),
.A2(n_336),
.B(n_337),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1559),
.Y(n_1666)
);

INVx8_ASAP7_75t_L g1667 ( 
.A(n_1613),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1644),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1589),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1567),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1651),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1561),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1548),
.B(n_339),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1574),
.B(n_340),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1650),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1604),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1560),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1573),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1580),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1642),
.B(n_344),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1617),
.A2(n_345),
.B(n_346),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1621),
.Y(n_1682)
);

AOI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1626),
.A2(n_553),
.B(n_347),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1568),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1579),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1605),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1583),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1625),
.B(n_348),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1592),
.B(n_349),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1588),
.A2(n_350),
.B(n_352),
.Y(n_1690)
);

AND2x4_ASAP7_75t_SL g1691 ( 
.A(n_1624),
.B(n_552),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1619),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1596),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1596),
.Y(n_1694)
);

AO21x1_ASAP7_75t_L g1695 ( 
.A1(n_1552),
.A2(n_353),
.B(n_354),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1568),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1643),
.Y(n_1697)
);

AO21x2_ASAP7_75t_L g1698 ( 
.A1(n_1627),
.A2(n_1646),
.B(n_1632),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1558),
.B(n_356),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1648),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1647),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1546),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1615),
.A2(n_357),
.B(n_359),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1571),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1629),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_SL g1706 ( 
.A1(n_1602),
.A2(n_364),
.B1(n_360),
.B2(n_361),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1568),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1647),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1616),
.B(n_365),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_1599),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1590),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1623),
.Y(n_1712)
);

OA21x2_ASAP7_75t_L g1713 ( 
.A1(n_1578),
.A2(n_551),
.B(n_366),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1586),
.Y(n_1714)
);

AOI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1585),
.A2(n_549),
.B(n_367),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1630),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1577),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1618),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1570),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1618),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1639),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1655),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1562),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1591),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1656),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1582),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1600),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1630),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1633),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1550),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1634),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1657),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1705),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1684),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1672),
.B(n_1598),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1663),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1705),
.B(n_1606),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1659),
.B(n_1595),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1679),
.A2(n_1543),
.B1(n_1622),
.B2(n_1607),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1692),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1667),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1677),
.B(n_1565),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1714),
.B(n_1576),
.Y(n_1743)
);

AO31x2_ASAP7_75t_L g1744 ( 
.A1(n_1693),
.A2(n_1641),
.A3(n_1603),
.B(n_1610),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1696),
.B(n_1637),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1670),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1692),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_1667),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1662),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1670),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1667),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1661),
.Y(n_1752)
);

AOI21x1_ASAP7_75t_L g1753 ( 
.A1(n_1694),
.A2(n_1597),
.B(n_1547),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1711),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1663),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1664),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1682),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1666),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1668),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1675),
.B(n_1620),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1710),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1671),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1697),
.B(n_1638),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1660),
.Y(n_1764)
);

NAND2xp33_ASAP7_75t_R g1765 ( 
.A(n_1669),
.B(n_1614),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1700),
.B(n_1649),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1678),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1685),
.B(n_1566),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1728),
.B(n_1652),
.Y(n_1769)
);

INVxp67_ASAP7_75t_SL g1770 ( 
.A(n_1686),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1662),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1687),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1676),
.B(n_1594),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1702),
.B(n_1631),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1704),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1679),
.A2(n_1563),
.B1(n_1654),
.B2(n_1636),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1723),
.B(n_1584),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1717),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1721),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1712),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1721),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1722),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1724),
.B(n_1554),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1722),
.Y(n_1784)
);

OAI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1707),
.A2(n_1718),
.B1(n_1720),
.B2(n_1716),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1725),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1719),
.B(n_1587),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1725),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1682),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1729),
.B(n_1640),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1729),
.B(n_1611),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1695),
.A2(n_1556),
.B1(n_1628),
.B2(n_1575),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1783),
.A2(n_1710),
.B1(n_1716),
.B2(n_1713),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1734),
.B(n_1707),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1741),
.B(n_1669),
.Y(n_1795)
);

BUFx3_ASAP7_75t_L g1796 ( 
.A(n_1761),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1782),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1749),
.B(n_1718),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1732),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1775),
.B(n_1727),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1752),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1771),
.B(n_1720),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1747),
.Y(n_1803)
);

INVxp67_ASAP7_75t_SL g1804 ( 
.A(n_1742),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1775),
.B(n_1713),
.Y(n_1805)
);

INVx4_ASAP7_75t_L g1806 ( 
.A(n_1757),
.Y(n_1806)
);

BUFx3_ASAP7_75t_L g1807 ( 
.A(n_1748),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1733),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1780),
.B(n_1701),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1756),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1757),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1758),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1778),
.B(n_1708),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1735),
.B(n_1698),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1763),
.B(n_1766),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1769),
.B(n_1726),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1759),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1784),
.Y(n_1818)
);

INVxp67_ASAP7_75t_L g1819 ( 
.A(n_1735),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1740),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1740),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1757),
.Y(n_1822)
);

INVx4_ASAP7_75t_L g1823 ( 
.A(n_1789),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1779),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1772),
.B(n_1698),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1781),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1737),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1788),
.Y(n_1828)
);

OAI21xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1739),
.A2(n_1776),
.B(n_1792),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1827),
.B(n_1773),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1829),
.A2(n_1739),
.B1(n_1774),
.B2(n_1760),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1799),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1798),
.B(n_1745),
.Y(n_1833)
);

INVxp67_ASAP7_75t_SL g1834 ( 
.A(n_1808),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1806),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1802),
.B(n_1738),
.Y(n_1836)
);

CKINVDCx20_ASAP7_75t_R g1837 ( 
.A(n_1796),
.Y(n_1837)
);

NOR2xp67_ASAP7_75t_L g1838 ( 
.A(n_1819),
.B(n_1786),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1794),
.B(n_1733),
.Y(n_1839)
);

OR2x6_ASAP7_75t_SL g1840 ( 
.A(n_1814),
.B(n_1783),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1801),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1807),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1806),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_L g1844 ( 
.A(n_1823),
.B(n_1774),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1822),
.B(n_1751),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1811),
.B(n_1754),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1820),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1820),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1823),
.B(n_1767),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1821),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1815),
.B(n_1743),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1821),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1825),
.B(n_1742),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1816),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1810),
.Y(n_1855)
);

AND2x4_ASAP7_75t_SL g1856 ( 
.A(n_1795),
.B(n_1789),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1812),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1797),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1804),
.B(n_1768),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1809),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1804),
.B(n_1768),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1818),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1809),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1824),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1845),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1832),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1845),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1831),
.A2(n_1814),
.B1(n_1793),
.B2(n_1819),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1859),
.B(n_1861),
.C(n_1793),
.Y(n_1869)
);

OAI21x1_ASAP7_75t_L g1870 ( 
.A1(n_1844),
.A2(n_1825),
.B(n_1805),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1838),
.Y(n_1871)
);

OAI211xp5_ASAP7_75t_L g1872 ( 
.A1(n_1853),
.A2(n_1601),
.B(n_1706),
.C(n_1805),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1860),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1832),
.Y(n_1874)
);

OA21x2_ASAP7_75t_L g1875 ( 
.A1(n_1847),
.A2(n_1800),
.B(n_1803),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1834),
.B(n_1813),
.Y(n_1876)
);

OAI321xp33_ASAP7_75t_L g1877 ( 
.A1(n_1848),
.A2(n_1785),
.A3(n_1753),
.B1(n_1760),
.B2(n_1800),
.C(n_1813),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1860),
.Y(n_1878)
);

INVx5_ASAP7_75t_L g1879 ( 
.A(n_1835),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1841),
.Y(n_1880)
);

NAND4xp25_ASAP7_75t_L g1881 ( 
.A(n_1842),
.B(n_1706),
.C(n_1765),
.D(n_1699),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1847),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_SL g1883 ( 
.A1(n_1856),
.A2(n_1690),
.B1(n_1789),
.B2(n_1688),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1839),
.B(n_1803),
.Y(n_1884)
);

AOI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1850),
.A2(n_1817),
.B1(n_1699),
.B2(n_1770),
.C(n_1787),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1833),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1840),
.A2(n_1777),
.B1(n_1730),
.B2(n_1689),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1884),
.B(n_1843),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1868),
.B(n_1849),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1871),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1879),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1879),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1866),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1876),
.B(n_1886),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1879),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1865),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1872),
.A2(n_1863),
.B1(n_1849),
.B2(n_1837),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_SL g1898 ( 
.A(n_1867),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1873),
.B(n_1830),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1874),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1878),
.B(n_1836),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1890),
.B(n_1880),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1893),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1894),
.B(n_1869),
.Y(n_1904)
);

NAND2x1p5_ASAP7_75t_L g1905 ( 
.A(n_1892),
.B(n_1682),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1893),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1891),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1900),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1895),
.Y(n_1909)
);

INVx3_ASAP7_75t_SL g1910 ( 
.A(n_1898),
.Y(n_1910)
);

INVxp67_ASAP7_75t_L g1911 ( 
.A(n_1889),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1899),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1888),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1901),
.B(n_1887),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1910),
.B(n_1897),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1914),
.B(n_1896),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1907),
.B(n_1882),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1913),
.B(n_1905),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1909),
.B(n_1882),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1904),
.B(n_1850),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1902),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1903),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1911),
.B(n_1912),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1908),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1908),
.B(n_1885),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1916),
.B(n_1906),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1915),
.B(n_1852),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1924),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1918),
.B(n_1852),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1924),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1917),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1919),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1921),
.B(n_1855),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1920),
.B(n_1846),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1922),
.Y(n_1935)
);

NAND2x1p5_ASAP7_75t_L g1936 ( 
.A(n_1923),
.B(n_1658),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1934),
.A2(n_1925),
.B1(n_1881),
.B2(n_1875),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1927),
.B(n_1877),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1930),
.Y(n_1939)
);

OAI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1928),
.A2(n_1875),
.B1(n_1857),
.B2(n_1862),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1926),
.Y(n_1941)
);

NAND3xp33_ASAP7_75t_L g1942 ( 
.A(n_1932),
.B(n_1883),
.C(n_1858),
.Y(n_1942)
);

AOI31xp33_ASAP7_75t_L g1943 ( 
.A1(n_1931),
.A2(n_1680),
.A3(n_1674),
.B(n_1612),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1929),
.B(n_1933),
.Y(n_1944)
);

AOI322xp5_ASAP7_75t_L g1945 ( 
.A1(n_1935),
.A2(n_1846),
.A3(n_1854),
.B1(n_1870),
.B2(n_1864),
.C1(n_1851),
.C2(n_1689),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1936),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1939),
.B(n_1826),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1941),
.B(n_1828),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1944),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_1762),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_1946),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1937),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1938),
.B(n_1736),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1940),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1945),
.B(n_1755),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1943),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1939),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1940),
.B(n_1691),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1941),
.B(n_1764),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1939),
.B(n_1746),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1951),
.A2(n_1709),
.B1(n_1691),
.B2(n_1731),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1957),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1956),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1952),
.B(n_1791),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1954),
.Y(n_1965)
);

INVxp67_ASAP7_75t_L g1966 ( 
.A(n_1949),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1959),
.B(n_1958),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1955),
.A2(n_1553),
.B(n_1703),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1948),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1950),
.Y(n_1970)
);

O2A1O1Ixp33_ASAP7_75t_SL g1971 ( 
.A1(n_1947),
.A2(n_1564),
.B(n_1673),
.C(n_1545),
.Y(n_1971)
);

INVx1_ASAP7_75t_SL g1972 ( 
.A(n_1960),
.Y(n_1972)
);

OAI211xp5_ASAP7_75t_SL g1973 ( 
.A1(n_1963),
.A2(n_1953),
.B(n_1608),
.C(n_1635),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1967),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1969),
.Y(n_1975)
);

OAI21xp33_ASAP7_75t_L g1976 ( 
.A1(n_1965),
.A2(n_1673),
.B(n_1790),
.Y(n_1976)
);

NOR2x1_ASAP7_75t_L g1977 ( 
.A(n_1962),
.B(n_1544),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1966),
.B(n_1750),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1970),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1964),
.B(n_1730),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_SL g1981 ( 
.A(n_1972),
.B(n_1645),
.C(n_1715),
.Y(n_1981)
);

NAND4xp25_ASAP7_75t_L g1982 ( 
.A(n_1974),
.B(n_1968),
.C(n_1961),
.D(n_1971),
.Y(n_1982)
);

A2O1A1Ixp33_ASAP7_75t_L g1983 ( 
.A1(n_1975),
.A2(n_1681),
.B(n_1665),
.C(n_1726),
.Y(n_1983)
);

XOR2x2_ASAP7_75t_L g1984 ( 
.A(n_1977),
.B(n_1980),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1979),
.B(n_1683),
.Y(n_1985)
);

AND3x2_ASAP7_75t_L g1986 ( 
.A(n_1978),
.B(n_368),
.C(n_369),
.Y(n_1986)
);

AND2x2_ASAP7_75t_SL g1987 ( 
.A(n_1973),
.B(n_1744),
.Y(n_1987)
);

OAI211xp5_ASAP7_75t_L g1988 ( 
.A1(n_1976),
.A2(n_1744),
.B(n_371),
.C(n_372),
.Y(n_1988)
);

NOR3xp33_ASAP7_75t_L g1989 ( 
.A(n_1981),
.B(n_370),
.C(n_373),
.Y(n_1989)
);

NOR2x1_ASAP7_75t_L g1990 ( 
.A(n_1979),
.B(n_374),
.Y(n_1990)
);

NAND4xp25_ASAP7_75t_L g1991 ( 
.A(n_1974),
.B(n_375),
.C(n_377),
.D(n_378),
.Y(n_1991)
);

NOR2x1_ASAP7_75t_L g1992 ( 
.A(n_1979),
.B(n_380),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1975),
.A2(n_1744),
.B1(n_384),
.B2(n_385),
.C(n_386),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1974),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1994),
.A2(n_381),
.B1(n_387),
.B2(n_388),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1990),
.B(n_1992),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1984),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1982),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1987),
.B(n_389),
.Y(n_1999)
);

NAND3xp33_ASAP7_75t_L g2000 ( 
.A(n_1986),
.B(n_390),
.C(n_391),
.Y(n_2000)
);

NAND3xp33_ASAP7_75t_L g2001 ( 
.A(n_1989),
.B(n_392),
.C(n_393),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1988),
.A2(n_394),
.B(n_395),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1985),
.A2(n_396),
.B(n_397),
.Y(n_2003)
);

AOI222xp33_ASAP7_75t_L g2004 ( 
.A1(n_1993),
.A2(n_398),
.B1(n_399),
.B2(n_401),
.C1(n_402),
.C2(n_403),
.Y(n_2004)
);

OAI31xp33_ASAP7_75t_L g2005 ( 
.A1(n_1991),
.A2(n_1983),
.A3(n_405),
.B(n_406),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1984),
.A2(n_404),
.B(n_407),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1994),
.B(n_408),
.Y(n_2007)
);

NAND3xp33_ASAP7_75t_L g2008 ( 
.A(n_1994),
.B(n_410),
.C(n_411),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1994),
.A2(n_412),
.B(n_414),
.Y(n_2009)
);

OAI211xp5_ASAP7_75t_L g2010 ( 
.A1(n_1994),
.A2(n_415),
.B(n_419),
.C(n_420),
.Y(n_2010)
);

NOR2x1_ASAP7_75t_L g2011 ( 
.A(n_2008),
.B(n_421),
.Y(n_2011)
);

AND4x1_ASAP7_75t_L g2012 ( 
.A(n_2006),
.B(n_423),
.C(n_424),
.D(n_425),
.Y(n_2012)
);

NOR3xp33_ASAP7_75t_SL g2013 ( 
.A(n_1997),
.B(n_427),
.C(n_429),
.Y(n_2013)
);

NOR2x1p5_ASAP7_75t_L g2014 ( 
.A(n_1996),
.B(n_430),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1999),
.Y(n_2015)
);

NOR2xp67_ASAP7_75t_L g2016 ( 
.A(n_2000),
.B(n_548),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2007),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1998),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2001),
.Y(n_2019)
);

NAND3xp33_ASAP7_75t_L g2020 ( 
.A(n_2004),
.B(n_2003),
.C(n_2005),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_2002),
.B(n_431),
.Y(n_2021)
);

NAND4xp75_ASAP7_75t_L g2022 ( 
.A(n_2009),
.B(n_1995),
.C(n_2010),
.D(n_435),
.Y(n_2022)
);

NOR2x1_ASAP7_75t_L g2023 ( 
.A(n_2008),
.B(n_432),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1997),
.B(n_434),
.Y(n_2024)
);

XNOR2xp5_ASAP7_75t_L g2025 ( 
.A(n_1997),
.B(n_436),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_2007),
.B(n_437),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_2007),
.B(n_439),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1996),
.B(n_440),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1996),
.Y(n_2029)
);

NAND3xp33_ASAP7_75t_L g2030 ( 
.A(n_1997),
.B(n_441),
.C(n_442),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_2014),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_2016),
.B(n_445),
.Y(n_2032)
);

NOR2x1_ASAP7_75t_L g2033 ( 
.A(n_2030),
.B(n_447),
.Y(n_2033)
);

AOI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_2018),
.A2(n_448),
.B1(n_452),
.B2(n_454),
.Y(n_2034)
);

AOI21xp33_ASAP7_75t_SL g2035 ( 
.A1(n_2025),
.A2(n_2021),
.B(n_2029),
.Y(n_2035)
);

OAI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_2013),
.A2(n_2020),
.B1(n_2015),
.B2(n_2012),
.C(n_2028),
.Y(n_2036)
);

OAI21xp33_ASAP7_75t_SL g2037 ( 
.A1(n_2022),
.A2(n_455),
.B(n_456),
.Y(n_2037)
);

NAND4xp75_ASAP7_75t_L g2038 ( 
.A(n_2024),
.B(n_2023),
.C(n_2011),
.D(n_2017),
.Y(n_2038)
);

NOR2x1_ASAP7_75t_L g2039 ( 
.A(n_2026),
.B(n_457),
.Y(n_2039)
);

NAND4xp75_ASAP7_75t_L g2040 ( 
.A(n_2019),
.B(n_2027),
.C(n_460),
.D(n_464),
.Y(n_2040)
);

OAI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_2018),
.A2(n_459),
.B1(n_465),
.B2(n_466),
.C(n_467),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_R g2042 ( 
.A(n_2025),
.B(n_469),
.Y(n_2042)
);

AND3x4_ASAP7_75t_L g2043 ( 
.A(n_2033),
.B(n_470),
.C(n_471),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_2031),
.B(n_547),
.Y(n_2044)
);

XNOR2x1_ASAP7_75t_L g2045 ( 
.A(n_2038),
.B(n_472),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_2032),
.B(n_473),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2039),
.Y(n_2047)
);

NOR2xp67_ASAP7_75t_L g2048 ( 
.A(n_2037),
.B(n_475),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2032),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2036),
.A2(n_477),
.B1(n_479),
.B2(n_480),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2045),
.Y(n_2051)
);

XNOR2xp5_ASAP7_75t_L g2052 ( 
.A(n_2043),
.B(n_2040),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_2048),
.Y(n_2053)
);

AND3x1_ASAP7_75t_L g2054 ( 
.A(n_2049),
.B(n_2034),
.C(n_2042),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2053),
.Y(n_2055)
);

NAND4xp75_ASAP7_75t_L g2056 ( 
.A(n_2054),
.B(n_2047),
.C(n_2046),
.D(n_2050),
.Y(n_2056)
);

OAI322xp33_ASAP7_75t_L g2057 ( 
.A1(n_2055),
.A2(n_2051),
.A3(n_2035),
.B1(n_2052),
.B2(n_2041),
.C1(n_2044),
.C2(n_487),
.Y(n_2057)
);

NAND4xp25_ASAP7_75t_SL g2058 ( 
.A(n_2056),
.B(n_481),
.C(n_482),
.D(n_483),
.Y(n_2058)
);

CKINVDCx20_ASAP7_75t_R g2059 ( 
.A(n_2057),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2058),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_2060),
.Y(n_2061)
);

AOI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_2059),
.A2(n_485),
.B1(n_486),
.B2(n_489),
.C(n_490),
.Y(n_2062)
);

OAI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_2061),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_2063)
);

HB1xp67_ASAP7_75t_L g2064 ( 
.A(n_2062),
.Y(n_2064)
);

NOR2xp67_ASAP7_75t_L g2065 ( 
.A(n_2064),
.B(n_497),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2063),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.Y(n_2066)
);

AOI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_2065),
.A2(n_502),
.B1(n_504),
.B2(n_505),
.Y(n_2067)
);

NAND3xp33_ASAP7_75t_L g2068 ( 
.A(n_2066),
.B(n_506),
.C(n_507),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2065),
.A2(n_508),
.B(n_509),
.Y(n_2069)
);

OAI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_2065),
.A2(n_511),
.B1(n_512),
.B2(n_514),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_2067),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2069),
.B(n_515),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_2070),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2068),
.Y(n_2074)
);

OR2x6_ASAP7_75t_L g2075 ( 
.A(n_2074),
.B(n_517),
.Y(n_2075)
);

OR2x6_ASAP7_75t_L g2076 ( 
.A(n_2071),
.B(n_519),
.Y(n_2076)
);

OR2x6_ASAP7_75t_L g2077 ( 
.A(n_2073),
.B(n_520),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2077),
.A2(n_2072),
.B(n_2076),
.Y(n_2078)
);

AOI211xp5_ASAP7_75t_L g2079 ( 
.A1(n_2078),
.A2(n_2075),
.B(n_521),
.C(n_522),
.Y(n_2079)
);


endmodule