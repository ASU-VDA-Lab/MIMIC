module real_jpeg_12437_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.B(n_20),
.C(n_26),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_2),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_48)
);

NAND2x1_ASAP7_75t_SL g70 ( 
.A(n_2),
.B(n_47),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_2),
.B(n_34),
.C(n_57),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_72),
.B(n_74),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_41),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_41),
.Y(n_68)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_76),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_75),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_65),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_16),
.B(n_65),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_42),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_29),
.Y(n_17)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_19),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_46)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_19),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B(n_23),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_22),
.B(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_22),
.B(n_30),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_23),
.A2(n_24),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_24),
.B(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B(n_38),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_30),
.A2(n_38),
.B(n_93),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_31),
.B(n_40),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_31),
.A2(n_39),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_33),
.B(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_48),
.B(n_49),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2x1_ASAP7_75t_R g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B1(n_60),
.B2(n_62),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_59),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_68),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.C(n_71),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_74),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_89),
.B(n_107),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_86),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_97),
.B(n_106),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_95),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_101),
.B(n_105),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);


endmodule