module fake_jpeg_2705_n_179 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_42),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_1),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_76),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_55),
.B(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_79),
.Y(n_96)
);

AOI22x1_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_57),
.B1(n_51),
.B2(n_53),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_55),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_80),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_67),
.B1(n_56),
.B2(n_62),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_89),
.B1(n_90),
.B2(n_98),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_67),
.B1(n_63),
.B2(n_58),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_56),
.B1(n_58),
.B2(n_57),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_97),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_49),
.B1(n_45),
.B2(n_51),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_80),
.B1(n_50),
.B2(n_51),
.Y(n_105)
);

OR2x4_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_45),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_51),
.B1(n_50),
.B2(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_53),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_108),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_113),
.B1(n_115),
.B2(n_119),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_82),
.B1(n_47),
.B2(n_54),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_2),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_118),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_54),
.B1(n_4),
.B2(n_5),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_40),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_95),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_39),
.C(n_38),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_9),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_6),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_137),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_92),
.B1(n_88),
.B2(n_85),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_131),
.B1(n_135),
.B2(n_17),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_7),
.B(n_8),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_18),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_36),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_33),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_31),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_134),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVxp33_ASAP7_75t_SL g145 ( 
.A(n_133),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_16),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_17),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_117),
.C(n_106),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.C(n_150),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_109),
.B1(n_119),
.B2(n_19),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_25),
.C(n_29),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_133),
.B1(n_121),
.B2(n_123),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_30),
.C(n_18),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

BUFx4f_ASAP7_75t_SL g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_155),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_20),
.C(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_20),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_159),
.Y(n_165)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_130),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_162),
.A2(n_147),
.B1(n_144),
.B2(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_168),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_146),
.C(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_124),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_163),
.B1(n_156),
.B2(n_158),
.Y(n_170)
);

OAI31xp33_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_151),
.A3(n_167),
.B(n_152),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_169),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_170),
.C(n_164),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_164),
.B(n_126),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_127),
.Y(n_179)
);


endmodule