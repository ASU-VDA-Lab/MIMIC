module fake_jpeg_10370_n_57 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_57);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_57;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g26 ( 
.A(n_6),
.B(n_4),
.CON(n_26),
.SN(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_0),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_12),
.Y(n_47)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_10),
.Y(n_44)
);

AO22x1_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_31),
.B1(n_27),
.B2(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_24),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_44),
.B(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_13),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_47),
.B1(n_45),
.B2(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_41),
.C(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_46),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_14),
.C(n_16),
.Y(n_56)
);

AOI221xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.C(n_21),
.Y(n_57)
);


endmodule