module fake_ibex_858_n_374 (n_85, n_84, n_64, n_3, n_73, n_65, n_95, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_97, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_92, n_96, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_374);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_95;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_97;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_92;
input n_96;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_374;

wire n_151;
wire n_171;
wire n_103;
wire n_204;
wire n_274;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_193;
wire n_108;
wire n_350;
wire n_165;
wire n_255;
wire n_175;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_239;
wire n_134;
wire n_371;
wire n_357;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_176;
wire n_216;
wire n_166;
wire n_163;
wire n_114;
wire n_236;
wire n_189;
wire n_317;
wire n_280;
wire n_340;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_113;
wire n_117;
wire n_265;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_210;
wire n_348;
wire n_220;
wire n_287;
wire n_243;
wire n_228;
wire n_147;
wire n_251;
wire n_373;
wire n_244;
wire n_343;
wire n_310;
wire n_323;
wire n_143;
wire n_106;
wire n_224;
wire n_183;
wire n_333;
wire n_110;
wire n_306;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_109;
wire n_127;
wire n_121;
wire n_325;
wire n_301;
wire n_296;
wire n_120;
wire n_168;
wire n_155;
wire n_315;
wire n_122;
wire n_116;
wire n_370;
wire n_289;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_235;
wire n_136;
wire n_261;
wire n_367;
wire n_221;
wire n_355;
wire n_281;
wire n_102;
wire n_99;
wire n_269;
wire n_156;
wire n_126;
wire n_356;
wire n_104;
wire n_141;
wire n_222;
wire n_186;
wire n_349;
wire n_295;
wire n_331;
wire n_230;
wire n_185;
wire n_352;
wire n_290;
wire n_174;
wire n_157;
wire n_219;
wire n_246;
wire n_146;
wire n_207;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_139;
wire n_275;
wire n_98;
wire n_129;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_347;
wire n_335;
wire n_263;
wire n_353;
wire n_359;
wire n_262;
wire n_299;
wire n_137;
wire n_338;
wire n_173;
wire n_363;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_257;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_365;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_329;
wire n_188;
wire n_200;
wire n_199;
wire n_308;
wire n_135;
wire n_283;
wire n_366;
wire n_111;
wire n_322;
wire n_227;
wire n_115;
wire n_248;
wire n_101;
wire n_190;
wire n_138;
wire n_238;
wire n_214;
wire n_332;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_225;
wire n_360;
wire n_272;
wire n_223;
wire n_320;
wire n_285;
wire n_247;
wire n_288;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_148;
wire n_342;
wire n_233;
wire n_118;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_178;
wire n_303;
wire n_362;
wire n_162;
wire n_240;
wire n_282;
wire n_266;
wire n_294;
wire n_112;
wire n_284;
wire n_172;
wire n_250;
wire n_313;
wire n_345;
wire n_119;
wire n_361;
wire n_319;
wire n_195;
wire n_212;
wire n_311;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_302;
wire n_344;
wire n_297;
wire n_252;
wire n_107;
wire n_149;
wire n_254;
wire n_213;
wire n_271;
wire n_241;
wire n_292;
wire n_364;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_160;
wire n_184;
wire n_232;

INVx2_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_9),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVxp33_ASAP7_75t_SL g105 ( 
.A(n_46),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

INVxp33_ASAP7_75t_SL g107 ( 
.A(n_51),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_16),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_5),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVxp33_ASAP7_75t_SL g112 ( 
.A(n_2),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_7),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_69),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_49),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_25),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_34),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_41),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_20),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_11),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_48),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_22),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_24),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_21),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_4),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_44),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_66),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_52),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_6),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_26),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_84),
.Y(n_150)
);

INVxp33_ASAP7_75t_SL g151 ( 
.A(n_12),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_79),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_42),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_82),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_17),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_55),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_27),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_45),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_60),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_67),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_32),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_37),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_36),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_31),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_39),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_97),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_75),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_38),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g177 ( 
.A(n_3),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_95),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_18),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_14),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_53),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_59),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_35),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_103),
.B(n_30),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_148),
.Y(n_204)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_136),
.B(n_0),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_146),
.A2(n_0),
.B1(n_1),
.B2(n_13),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_137),
.B(n_1),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_120),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_112),
.A2(n_177),
.B1(n_163),
.B2(n_173),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_126),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_154),
.B(n_28),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_122),
.B(n_47),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_117),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_165),
.A2(n_65),
.B1(n_81),
.B2(n_91),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_149),
.B(n_157),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_100),
.B(n_161),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_140),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_141),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_142),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_162),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_143),
.B(n_166),
.Y(n_241)
);

BUFx8_ASAP7_75t_L g242 ( 
.A(n_144),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_147),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_155),
.A2(n_168),
.B1(n_186),
.B2(n_185),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_159),
.B(n_167),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_200),
.A2(n_105),
.B1(n_107),
.B2(n_151),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_201),
.A2(n_171),
.B(n_183),
.C(n_182),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_200),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_152),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

AO22x2_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_110),
.B1(n_170),
.B2(n_187),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_125),
.B1(n_130),
.B2(n_174),
.Y(n_264)
);

AO22x2_ASAP7_75t_L g265 ( 
.A1(n_189),
.A2(n_180),
.B1(n_179),
.B2(n_110),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_206),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_230),
.Y(n_272)
);

NAND2x1p5_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_164),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_217),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_134),
.B1(n_138),
.B2(n_150),
.Y(n_276)
);

AO22x2_ASAP7_75t_L g277 ( 
.A1(n_191),
.A2(n_158),
.B1(n_175),
.B2(n_176),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_192),
.B(n_178),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_237),
.B1(n_238),
.B2(n_234),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_235),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_194),
.B(n_209),
.Y(n_282)
);

OR2x6_ASAP7_75t_L g283 ( 
.A(n_231),
.B(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_224),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_215),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

AO22x2_ASAP7_75t_L g291 ( 
.A1(n_196),
.A2(n_247),
.B1(n_239),
.B2(n_243),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_190),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_202),
.B(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_211),
.Y(n_295)
);

AO22x2_ASAP7_75t_L g296 ( 
.A1(n_214),
.A2(n_229),
.B1(n_245),
.B2(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_190),
.Y(n_297)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_195),
.Y(n_299)
);

BUFx8_ASAP7_75t_L g300 ( 
.A(n_197),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_197),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_197),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_226),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_250),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_195),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_198),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_198),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_266),
.A2(n_236),
.B1(n_240),
.B2(n_272),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_278),
.B(n_236),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_259),
.B(n_240),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_253),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_256),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_273),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_269),
.B(n_279),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_283),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_260),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_297),
.A2(n_252),
.B(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_251),
.B(n_262),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_262),
.B(n_290),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_283),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_317),
.B1(n_292),
.B2(n_319),
.Y(n_326)
);

NAND2x1p5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_280),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_271),
.B(n_286),
.C(n_285),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_296),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_262),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_314),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_249),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_276),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_264),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_314),
.B(n_300),
.Y(n_339)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_265),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_277),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_257),
.Y(n_343)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_331),
.A2(n_303),
.B(n_301),
.C(n_304),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_338),
.A2(n_321),
.B1(n_270),
.B2(n_284),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_334),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_263),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_329),
.Y(n_348)
);

NOR2x1_ASAP7_75t_SL g349 ( 
.A(n_326),
.B(n_335),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_288),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_311),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_344),
.A2(n_332),
.B(n_341),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_348),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_325),
.Y(n_355)
);

OR2x6_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_340),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_343),
.A2(n_330),
.B(n_310),
.C(n_334),
.Y(n_357)
);

NAND4xp25_ASAP7_75t_L g358 ( 
.A(n_351),
.B(n_339),
.C(n_309),
.D(n_306),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_354),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_350),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_358),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_356),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_359),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_362),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_360),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_363),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_366),
.B(n_361),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_367),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_368),
.A2(n_365),
.B1(n_339),
.B2(n_357),
.Y(n_369)
);

AOI211xp5_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_353),
.B(n_345),
.C(n_346),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_370),
.B(n_352),
.Y(n_371)
);

OR3x1_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_349),
.C(n_299),
.Y(n_372)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_372),
.Y(n_373)
);

AOI221xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_347),
.B1(n_281),
.B2(n_333),
.C(n_327),
.Y(n_374)
);


endmodule