module fake_jpeg_27881_n_194 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_194);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_26),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_23),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_56),
.Y(n_63)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_20),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_30),
.B1(n_33),
.B2(n_16),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_30),
.B1(n_17),
.B2(n_24),
.Y(n_70)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_65),
.B(n_69),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_48),
.B1(n_59),
.B2(n_61),
.Y(n_97)
);

AOI32xp33_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_32),
.A3(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_19),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_27),
.B1(n_20),
.B2(n_24),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_80),
.B(n_21),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_18),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_84),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_34),
.Y(n_80)
);

OA22x2_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_83),
.Y(n_87)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_38),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_55),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_91),
.B(n_97),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_57),
.B(n_56),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_103),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_55),
.C(n_37),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_104),
.C(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_21),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_19),
.C(n_26),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_76),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_84),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_113),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_79),
.B(n_80),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_64),
.B1(n_83),
.B2(n_88),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_120),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_123),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_85),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_81),
.B1(n_48),
.B2(n_61),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_98),
.B1(n_93),
.B2(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_127),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_64),
.Y(n_123)
);

AO22x1_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_81),
.B1(n_61),
.B2(n_35),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_86),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_99),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_136),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_96),
.B(n_92),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_139),
.B(n_115),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_143),
.B1(n_140),
.B2(n_138),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_12),
.A3(n_11),
.B1(n_10),
.B2(n_9),
.C1(n_8),
.C2(n_6),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_141),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_88),
.B(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_89),
.C(n_67),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_62),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_109),
.B1(n_124),
.B2(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_19),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_0),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_138),
.A2(n_121),
.B1(n_109),
.B2(n_115),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_150),
.B1(n_154),
.B2(n_135),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_141),
.Y(n_161)
);

FAx1_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_124),
.CI(n_116),
.CON(n_149),
.SN(n_149)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_151),
.B(n_158),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_117),
.B(n_108),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_159),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_26),
.B1(n_72),
.B2(n_2),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_11),
.B1(n_9),
.B2(n_4),
.C(n_5),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_1),
.Y(n_169)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_1),
.B(n_4),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_130),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_6),
.B(n_7),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_130),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_169),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_145),
.C(n_133),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_145),
.C(n_133),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_146),
.C(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_149),
.C(n_152),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_166),
.C(n_162),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_165),
.A2(n_159),
.B(n_148),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_5),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_182),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_170),
.B(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_187),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_183),
.Y(n_187)
);

OAI221xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_164),
.B1(n_179),
.B2(n_180),
.C(n_171),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_6),
.CI(n_7),
.CON(n_189),
.SN(n_189)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_187),
.B(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_190),
.Y(n_194)
);


endmodule