module fake_jpeg_1846_n_178 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_65),
.Y(n_74)
);

NAND2x1_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_0),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_63),
.Y(n_75)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_63),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_53),
.B1(n_46),
.B2(n_47),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_46),
.B1(n_53),
.B2(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_78),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_54),
.B1(n_57),
.B2(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_49),
.B1(n_59),
.B2(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_9),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_48),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_62),
.B1(n_59),
.B2(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_59),
.B1(n_65),
.B2(n_3),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_73),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_2),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_9),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_102),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_72),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_111),
.C(n_13),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_70),
.B1(n_73),
.B2(n_6),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_105),
.B(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_104),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_5),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_8),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_22),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_23),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_10),
.B(n_11),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_10),
.B(n_12),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_81),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_34),
.C(n_33),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_81),
.B(n_11),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_105),
.B(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_24),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_128),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_19),
.B(n_115),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_29),
.B1(n_38),
.B2(n_37),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_130),
.A2(n_20),
.B1(n_36),
.B2(n_35),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_130),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_144),
.B1(n_145),
.B2(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_143),
.Y(n_151)
);

XNOR2x2_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_13),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_117),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_43),
.Y(n_139)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_138),
.A3(n_141),
.B1(n_144),
.B2(n_147),
.C1(n_149),
.C2(n_140),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_120),
.C(n_129),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_31),
.B(n_30),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_148),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_154),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_155),
.A2(n_158),
.B(n_159),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_116),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_139),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_142),
.B(n_149),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_152),
.Y(n_168)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_168),
.A2(n_169),
.B1(n_162),
.B2(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_165),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_170),
.C(n_161),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_171),
.B(n_158),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_171),
.CI(n_151),
.CON(n_177),
.SN(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_176),
.Y(n_178)
);


endmodule