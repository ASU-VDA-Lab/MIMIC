module real_jpeg_7211_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_1),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_1),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_1),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_2),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_2),
.Y(n_190)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_2),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_3),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_3),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_3),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_3),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_3),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_3),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_4),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_4),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_4),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_4),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_5),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_5),
.B(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_5),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_5),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_5),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_5),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_5),
.B(n_407),
.Y(n_406)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_7),
.Y(n_147)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_7),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_7),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_7),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_7),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_8),
.B(n_151),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_8),
.B(n_26),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_8),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_8),
.B(n_67),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_8),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_8),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_8),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_8),
.B(n_441),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_9),
.Y(n_149)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_11),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_11),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_11),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_11),
.B(n_443),
.Y(n_442)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_12),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_12),
.Y(n_292)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_12),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_81),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_13),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_13),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_13),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_13),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_13),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_14),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_14),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_14),
.B(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_14),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_14),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_14),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_14),
.B(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_15),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_15),
.Y(n_277)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_15),
.Y(n_427)
);

BUFx5_ASAP7_75t_L g441 ( 
.A(n_15),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_162),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_161),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_20),
.B(n_102),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_47),
.B2(n_48),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.C(n_46),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_24),
.A2(n_25),
.B1(n_46),
.B2(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_27),
.B(n_223),
.Y(n_222)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_30),
.B(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.C(n_42),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_31),
.A2(n_37),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_31),
.Y(n_141)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_35),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_35),
.Y(n_262)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_36),
.Y(n_181)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_37),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_37),
.A2(n_140),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_37),
.B(n_145),
.C(n_188),
.Y(n_326)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_40),
.Y(n_247)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_41),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_42),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_42),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_46),
.A2(n_88),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_46),
.B(n_346),
.C(n_363),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_46),
.A2(n_88),
.B1(n_150),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_72),
.B2(n_73),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_54),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.C(n_64),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_90),
.C(n_95),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_64),
.B1(n_65),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_56),
.A2(n_95),
.B1(n_96),
.B2(n_101),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_56),
.A2(n_101),
.B1(n_226),
.B2(n_234),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_56),
.B(n_119),
.C(n_227),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_57),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_58),
.Y(n_383)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_59),
.Y(n_275)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_59),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_65),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_64),
.A2(n_65),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_65),
.B(n_201),
.C(n_206),
.Y(n_289)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_68),
.Y(n_231)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_78),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_97),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_83),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_76),
.A2(n_77),
.B1(n_271),
.B2(n_278),
.Y(n_270)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_77),
.B(n_348),
.C(n_349),
.Y(n_347)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_83),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_130),
.C(n_136),
.Y(n_156)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.C(n_99),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_85),
.A2(n_86),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_88),
.B(n_144),
.C(n_150),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_89),
.B(n_99),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_90),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_94),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_96),
.B1(n_113),
.B2(n_117),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_95),
.A2(n_96),
.B1(n_188),
.B2(n_282),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_96),
.B(n_107),
.C(n_113),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_96),
.B(n_183),
.C(n_188),
.Y(n_182)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_97),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_98),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_152),
.C(n_158),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_103),
.B(n_152),
.CI(n_158),
.CON(n_485),
.SN(n_485)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_137),
.C(n_143),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_104),
.A2(n_105),
.B1(n_488),
.B2(n_489),
.Y(n_487)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_118),
.C(n_127),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_106),
.B(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_145),
.C(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_113),
.B(n_307),
.C(n_311),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_113),
.A2(n_117),
.B1(n_145),
.B2(n_283),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_113),
.A2(n_117),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_118),
.B(n_127),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_123),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_119),
.A2(n_227),
.B1(n_232),
.B2(n_233),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_119),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_119),
.A2(n_232),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_121),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_122),
.B(n_123),
.Y(n_328)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_132),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_132),
.B(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_132),
.B(n_257),
.C(n_259),
.Y(n_269)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_137),
.B(n_143),
.Y(n_488)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_144),
.B(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_145),
.A2(n_188),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_145),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_145),
.A2(n_283),
.B1(n_393),
.B2(n_394),
.Y(n_411)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_148),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_148),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_150),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_153),
.A2(n_154),
.B1(n_491),
.B2(n_492),
.Y(n_490)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_156),
.B(n_157),
.Y(n_492)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_483),
.B(n_497),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_352),
.B(n_368),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_320),
.B(n_351),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_297),
.B(n_319),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_166),
.B(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_264),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_167),
.B(n_264),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_224),
.C(n_252),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_168),
.B(n_318),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_168),
.Y(n_500)
);

FAx1_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_198),
.CI(n_208),
.CON(n_168),
.SN(n_168)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_169),
.B(n_198),
.C(n_208),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_182),
.C(n_191),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_170),
.B(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_172),
.B(n_175),
.C(n_179),
.Y(n_263)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_182),
.A2(n_191),
.B1(n_192),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_182),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_183),
.B(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_188),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx8_ASAP7_75t_L g378 ( 
.A(n_190),
.Y(n_378)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_313)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_201),
.A2(n_207),
.B1(n_240),
.B2(n_241),
.Y(n_401)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_210),
.B(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_209),
.B(n_215),
.C(n_222),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_213),
.B(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_219),
.Y(n_417)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_220),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_223),
.B(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_223),
.B(n_399),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_223),
.B(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_224),
.B(n_252),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.C(n_237),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_225),
.A2(n_235),
.B1(n_236),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_227),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_237),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.C(n_248),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_238),
.A2(n_239),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_243),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_471)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_255),
.C(n_263),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_265),
.B(n_267),
.C(n_296),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_284),
.B1(n_295),
.B2(n_296),
.Y(n_266)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_279),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_269),
.B(n_270),
.C(n_279),
.Y(n_337)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_276),
.Y(n_349)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_283),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_293),
.C(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_317),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_298),
.B(n_317),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_303),
.C(n_314),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_299),
.A2(n_300),
.B1(n_476),
.B2(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_303),
.B(n_314),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.C(n_313),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_304),
.B(n_463),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_306),
.B(n_313),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_307),
.A2(n_308),
.B1(n_311),
.B2(n_312),
.Y(n_390)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_321),
.B(n_352),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_322),
.B(n_323),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_353),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_323),
.B(n_353),
.Y(n_482)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_336),
.CI(n_350),
.CON(n_323),
.SN(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_330),
.B2(n_331),
.Y(n_325)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_331),
.C(n_332),
.Y(n_360)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_339),
.C(n_341),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

INVx8_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_354),
.B(n_356),
.C(n_358),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_361),
.B2(n_367),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_359),
.B(n_362),
.C(n_364),
.Y(n_493)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_361),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

OAI31xp33_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_479),
.A3(n_480),
.B(n_482),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_473),
.B(n_478),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_458),
.B(n_472),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_412),
.B(n_457),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_402),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_373),
.B(n_402),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_391),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_388),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_375),
.B(n_388),
.C(n_391),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.C(n_384),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_377),
.B1(n_379),
.B2(n_380),
.Y(n_404)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_384),
.B(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_397),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_392),
.B(n_467),
.C(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_401),
.Y(n_397)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_398),
.Y(n_467)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_405),
.C(n_411),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_403),
.B(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_405),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_405),
.A2(n_411),
.B1(n_449),
.B2(n_455),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_406),
.Y(n_447)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_451),
.B(n_456),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_437),
.B(n_450),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_422),
.B(n_436),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_433),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_433),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_428),
.B(n_432),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_428),
.Y(n_432)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_432),
.A2(n_439),
.B1(n_444),
.B2(n_445),
.Y(n_438)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_446),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_446),
.Y(n_450)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_439),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_442),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_440),
.A2(n_442),
.B(n_444),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_448),
.B(n_449),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_453),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_460),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_462),
.B1(n_464),
.B2(n_465),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_466),
.C(n_469),
.Y(n_474)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_474),
.B(n_475),
.Y(n_478)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_476),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_494),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_484),
.A2(n_498),
.B(n_499),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_486),
.Y(n_499)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_485),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_490),
.C(n_493),
.Y(n_486)
);

FAx1_ASAP7_75t_SL g496 ( 
.A(n_487),
.B(n_490),
.CI(n_493),
.CON(n_496),
.SN(n_496)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_488),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_496),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g501 ( 
.A(n_496),
.Y(n_501)
);


endmodule