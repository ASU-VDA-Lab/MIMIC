module fake_netlist_5_1548_n_1495 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1495);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1495;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_370;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_1319;
wire n_561;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_157),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_88),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_290),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_241),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_231),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_31),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_46),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_0),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_270),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_342),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_117),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_341),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_17),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_53),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_208),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_345),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_144),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_87),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_124),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_330),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_77),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_332),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_103),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_359),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_174),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_322),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_129),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_179),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_257),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_141),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_236),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_221),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_259),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_52),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_152),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_293),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_357),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_266),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_323),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_143),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_277),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_67),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_73),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_244),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_38),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_8),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_235),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_265),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_227),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_201),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_297),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_107),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_81),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_4),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_263),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_312),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_100),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_313),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_249),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_62),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_28),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_302),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_106),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_147),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_238),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_316),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_348),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_108),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_296),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_123),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_43),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_203),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_146),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_264),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_127),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_226),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_258),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_58),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_156),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_267),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_306),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_50),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_169),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_134),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_331),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_168),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_254),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_155),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_149),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_138),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_262),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_343),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_56),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_75),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_337),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_109),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_111),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_274),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_354),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_298),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_280),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_98),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_177),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_275),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_202),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_171),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_130),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_287),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_92),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_172),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_185),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_248),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_308),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_45),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_333),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_349),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_19),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_338),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_242),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_10),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_46),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_0),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_87),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_116),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_200),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_145),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_347),
.Y(n_490)
);

BUFx10_ASAP7_75t_L g491 ( 
.A(n_289),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_12),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_170),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_269),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_340),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_113),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_50),
.Y(n_497)
);

BUFx5_ASAP7_75t_L g498 ( 
.A(n_163),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_5),
.Y(n_499)
);

BUFx5_ASAP7_75t_L g500 ( 
.A(n_324),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_10),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_247),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_222),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_22),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_178),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_11),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_176),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_303),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_310),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_60),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_304),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_166),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_355),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_44),
.Y(n_514)
);

CKINVDCx14_ASAP7_75t_R g515 ( 
.A(n_81),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_276),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_328),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_164),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_180),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_126),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_228),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_230),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_22),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_77),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_1),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_283),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_15),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_90),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_311),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_210),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_307),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_317),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_102),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_115),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_60),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_84),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_105),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_99),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_40),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_294),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_17),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_209),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_29),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_272),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_216),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_318),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g547 ( 
.A(n_159),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_346),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_232),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_173),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_161),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_55),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_295),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_84),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_195),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_89),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_28),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_260),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_24),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_158),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_88),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_214),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_37),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_184),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_175),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_5),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_59),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_186),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_233),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_135),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_71),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_75),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_339),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_142),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_212),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_191),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_55),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_309),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_151),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_160),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_91),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_181),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_80),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_204),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_120),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_321),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_70),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_292),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_15),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_268),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_253),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_278),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_69),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_36),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_300),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_206),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_234),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_515),
.B(n_1),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_372),
.B(n_2),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_375),
.B(n_2),
.Y(n_600)
);

BUFx12f_ASAP7_75t_L g601 ( 
.A(n_468),
.Y(n_601)
);

NOR2x1_ASAP7_75t_L g602 ( 
.A(n_511),
.B(n_93),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_372),
.Y(n_603)
);

BUFx12f_ASAP7_75t_L g604 ( 
.A(n_468),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_374),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_375),
.B(n_421),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_491),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_511),
.B(n_3),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_387),
.B(n_462),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_421),
.B(n_431),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_431),
.B(n_3),
.Y(n_611)
);

BUFx8_ASAP7_75t_SL g612 ( 
.A(n_557),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_528),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_508),
.B(n_4),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_394),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_374),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_491),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_372),
.B(n_6),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_508),
.B(n_6),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_372),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_360),
.Y(n_621)
);

BUFx12f_ASAP7_75t_L g622 ( 
.A(n_550),
.Y(n_622)
);

BUFx12f_ASAP7_75t_L g623 ( 
.A(n_550),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_519),
.B(n_7),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_524),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_570),
.B(n_7),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_568),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_524),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_374),
.Y(n_629)
);

BUFx12f_ASAP7_75t_L g630 ( 
.A(n_568),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_513),
.B(n_8),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_524),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_528),
.B(n_9),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_547),
.B(n_9),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_374),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_378),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_362),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_404),
.B(n_11),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_393),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_394),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_393),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_378),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_581),
.B(n_12),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_579),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_545),
.B(n_13),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_552),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_366),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_361),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_378),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_378),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_408),
.Y(n_652)
);

BUFx12f_ASAP7_75t_L g653 ( 
.A(n_579),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_445),
.B(n_13),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_367),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_513),
.B(n_14),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_569),
.B(n_16),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_405),
.B(n_16),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_588),
.B(n_18),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_393),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_363),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_373),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_393),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_365),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_559),
.B(n_18),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_484),
.B(n_19),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_380),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_408),
.Y(n_668)
);

BUFx12f_ASAP7_75t_L g669 ( 
.A(n_377),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_559),
.B(n_20),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_567),
.B(n_20),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_402),
.Y(n_672)
);

BUFx12f_ASAP7_75t_L g673 ( 
.A(n_406),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_408),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_408),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_415),
.Y(n_676)
);

BUFx8_ASAP7_75t_SL g677 ( 
.A(n_403),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_567),
.B(n_21),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_368),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_525),
.B(n_21),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_370),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_461),
.B(n_23),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_371),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_393),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_464),
.B(n_23),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_364),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_414),
.B(n_24),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_422),
.B(n_25),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_433),
.B(n_25),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_383),
.B(n_26),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_384),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_423),
.B(n_26),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_399),
.B(n_27),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_393),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_390),
.B(n_27),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_395),
.B(n_29),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_410),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_376),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_498),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_411),
.B(n_30),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_485),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_499),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_413),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_501),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_379),
.Y(n_705)
);

INVx5_ASAP7_75t_L g706 ( 
.A(n_498),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_416),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_504),
.B(n_30),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_456),
.B(n_31),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_510),
.B(n_32),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_477),
.B(n_32),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_417),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_426),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_437),
.B(n_33),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_498),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_381),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_438),
.Y(n_717)
);

NOR2x1_ASAP7_75t_L g718 ( 
.A(n_442),
.B(n_94),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_514),
.B(n_33),
.Y(n_719)
);

INVx5_ASAP7_75t_L g720 ( 
.A(n_498),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_535),
.B(n_34),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_539),
.B(n_34),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_556),
.B(n_35),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_439),
.B(n_35),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_498),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_480),
.B(n_36),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_540),
.B(n_37),
.Y(n_727)
);

BUFx12f_ASAP7_75t_L g728 ( 
.A(n_483),
.Y(n_728)
);

INVxp33_ASAP7_75t_SL g729 ( 
.A(n_486),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_382),
.Y(n_730)
);

INVx5_ASAP7_75t_L g731 ( 
.A(n_498),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_443),
.B(n_38),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_385),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_444),
.Y(n_734)
);

INVx5_ASAP7_75t_L g735 ( 
.A(n_500),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_606),
.Y(n_736)
);

BUFx10_ASAP7_75t_L g737 ( 
.A(n_645),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_SL g738 ( 
.A1(n_644),
.A2(n_497),
.B1(n_506),
.B2(n_492),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_644),
.A2(n_527),
.B1(n_536),
.B2(n_523),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_625),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_649),
.B(n_664),
.Y(n_741)
);

AO22x2_ASAP7_75t_L g742 ( 
.A1(n_608),
.A2(n_577),
.B1(n_594),
.B2(n_563),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_634),
.A2(n_401),
.B1(n_427),
.B2(n_369),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_598),
.B(n_447),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_SL g745 ( 
.A1(n_624),
.A2(n_543),
.B1(n_554),
.B2(n_541),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_SL g746 ( 
.A(n_626),
.B(n_441),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_638),
.A2(n_561),
.B1(n_572),
.B2(n_566),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_603),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_620),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_676),
.B(n_386),
.Y(n_750)
);

NAND3x1_ASAP7_75t_L g751 ( 
.A(n_654),
.B(n_693),
.C(n_690),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_613),
.B(n_583),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_654),
.A2(n_474),
.B1(n_475),
.B2(n_454),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_632),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_661),
.B(n_388),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_609),
.A2(n_512),
.B1(n_558),
.B2(n_553),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_679),
.B(n_389),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_690),
.A2(n_585),
.B1(n_573),
.B2(n_589),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_693),
.A2(n_593),
.B1(n_571),
.B2(n_587),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_639),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_700),
.A2(n_457),
.B1(n_392),
.B2(n_396),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_698),
.B(n_705),
.Y(n_762)
);

AO22x2_ASAP7_75t_L g763 ( 
.A1(n_608),
.A2(n_458),
.B1(n_463),
.B2(n_449),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_607),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_646),
.A2(n_469),
.B1(n_470),
.B2(n_466),
.Y(n_765)
);

AO22x1_ASAP7_75t_L g766 ( 
.A1(n_631),
.A2(n_597),
.B1(n_479),
.B2(n_481),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_SL g767 ( 
.A1(n_646),
.A2(n_482),
.B1(n_487),
.B2(n_473),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_631),
.B(n_488),
.Y(n_768)
);

OAI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_659),
.A2(n_494),
.B1(n_495),
.B2(n_490),
.Y(n_769)
);

AO22x2_ASAP7_75t_L g770 ( 
.A1(n_657),
.A2(n_507),
.B1(n_534),
.B2(n_502),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_625),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_700),
.A2(n_397),
.B1(n_398),
.B2(n_391),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_659),
.A2(n_562),
.B1(n_574),
.B2(n_549),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_621),
.B(n_637),
.Y(n_774)
);

CKINVDCx6p67_ASAP7_75t_R g775 ( 
.A(n_601),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_628),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_657),
.A2(n_582),
.B1(n_578),
.B2(n_41),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_724),
.A2(n_407),
.B1(n_409),
.B2(n_400),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_669),
.B(n_39),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_628),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_681),
.B(n_412),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_729),
.B(n_418),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_724),
.A2(n_420),
.B1(n_424),
.B2(n_419),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_727),
.A2(n_428),
.B1(n_429),
.B2(n_425),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_716),
.B(n_430),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_730),
.B(n_683),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_683),
.B(n_432),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_600),
.A2(n_435),
.B1(n_436),
.B2(n_434),
.Y(n_788)
);

AO22x2_ASAP7_75t_L g789 ( 
.A1(n_656),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_616),
.Y(n_790)
);

AO22x2_ASAP7_75t_L g791 ( 
.A1(n_682),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_727),
.A2(n_446),
.B1(n_448),
.B2(n_440),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_617),
.B(n_450),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_615),
.Y(n_794)
);

OR2x6_ASAP7_75t_L g795 ( 
.A(n_673),
.B(n_42),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_733),
.B(n_627),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_728),
.A2(n_452),
.B1(n_453),
.B2(n_451),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_600),
.A2(n_459),
.B1(n_460),
.B2(n_455),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_633),
.B(n_465),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_677),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_616),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_615),
.B(n_467),
.Y(n_802)
);

AO22x2_ASAP7_75t_L g803 ( 
.A1(n_682),
.A2(n_48),
.B1(n_45),
.B2(n_47),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_611),
.A2(n_472),
.B1(n_476),
.B2(n_471),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_680),
.A2(n_489),
.B1(n_493),
.B2(n_478),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_SL g806 ( 
.A1(n_611),
.A2(n_503),
.B1(n_505),
.B2(n_496),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_641),
.B(n_509),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_614),
.A2(n_517),
.B1(n_518),
.B2(n_516),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_641),
.B(n_520),
.Y(n_809)
);

OA22x2_ASAP7_75t_L g810 ( 
.A1(n_672),
.A2(n_521),
.B1(n_526),
.B2(n_522),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_616),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_688),
.B(n_529),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_689),
.A2(n_711),
.B1(n_726),
.B2(n_709),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_612),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_658),
.B(n_530),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_666),
.B(n_531),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_648),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_L g818 ( 
.A1(n_614),
.A2(n_533),
.B1(n_537),
.B2(n_532),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_605),
.B(n_538),
.Y(n_819)
);

AO22x2_ASAP7_75t_L g820 ( 
.A1(n_685),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_635),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_604),
.B(n_49),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_622),
.A2(n_542),
.B1(n_546),
.B2(n_544),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_635),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_619),
.A2(n_551),
.B1(n_555),
.B2(n_548),
.Y(n_825)
);

OA22x2_ASAP7_75t_L g826 ( 
.A1(n_672),
.A2(n_560),
.B1(n_565),
.B2(n_564),
.Y(n_826)
);

BUFx10_ASAP7_75t_L g827 ( 
.A(n_695),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_623),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_756),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_817),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_790),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_736),
.B(n_630),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_801),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_762),
.B(n_768),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_741),
.B(n_802),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_811),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_807),
.B(n_647),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_768),
.B(n_640),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_737),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_809),
.B(n_799),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_821),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_824),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_783),
.B(n_653),
.Y(n_843)
);

XNOR2x2_ASAP7_75t_L g844 ( 
.A(n_789),
.B(n_665),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_740),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_780),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_775),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_771),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_776),
.Y(n_849)
);

XNOR2xp5_ASAP7_75t_L g850 ( 
.A(n_753),
.B(n_695),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_782),
.B(n_696),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_744),
.B(n_642),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_749),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_786),
.B(n_696),
.Y(n_854)
);

AND2x6_ASAP7_75t_L g855 ( 
.A(n_813),
.B(n_602),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_794),
.B(n_714),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_796),
.B(n_647),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_754),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_787),
.B(n_605),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_748),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_760),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_764),
.B(n_702),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_800),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_827),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_752),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_759),
.B(n_714),
.Y(n_866)
);

AND2x6_ASAP7_75t_L g867 ( 
.A(n_774),
.B(n_732),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_827),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_828),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_743),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_819),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_742),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_742),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_765),
.A2(n_610),
.B(n_606),
.Y(n_874)
);

XOR2xp5_ASAP7_75t_L g875 ( 
.A(n_758),
.B(n_575),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_816),
.Y(n_876)
);

XOR2x2_ASAP7_75t_L g877 ( 
.A(n_751),
.B(n_687),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_755),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_757),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_763),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_763),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_770),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_789),
.B(n_687),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_770),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_772),
.B(n_732),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_750),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_810),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_826),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_812),
.Y(n_889)
);

XOR2x2_ASAP7_75t_L g890 ( 
.A(n_761),
.B(n_692),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_815),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_746),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_815),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_764),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_781),
.Y(n_895)
);

XOR2x2_ASAP7_75t_L g896 ( 
.A(n_738),
.B(n_692),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_785),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_766),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_778),
.B(n_610),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_767),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_769),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_791),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_791),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_779),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_793),
.B(n_655),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_803),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_779),
.B(n_662),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_803),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_820),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_737),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_820),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_777),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_777),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_784),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_792),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_739),
.B(n_686),
.Y(n_916)
);

AND2x2_ASAP7_75t_SL g917 ( 
.A(n_797),
.B(n_685),
.Y(n_917)
);

XOR2xp5_ASAP7_75t_L g918 ( 
.A(n_814),
.B(n_576),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_745),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_747),
.B(n_599),
.Y(n_920)
);

XNOR2x1_ASAP7_75t_L g921 ( 
.A(n_795),
.B(n_708),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_805),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_773),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_853),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_862),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_835),
.B(n_702),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_840),
.B(n_667),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_899),
.B(n_788),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_894),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_867),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_851),
.B(n_806),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_898),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_837),
.B(n_701),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_854),
.B(n_798),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_852),
.A2(n_808),
.B(n_804),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_858),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_852),
.B(n_818),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_834),
.B(n_718),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_883),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_830),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_867),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_834),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_838),
.A2(n_874),
.B(n_885),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_867),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_891),
.B(n_704),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_867),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_876),
.B(n_599),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_864),
.Y(n_948)
);

INVxp33_ASAP7_75t_L g949 ( 
.A(n_857),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_886),
.B(n_618),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_893),
.B(n_795),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_887),
.B(n_888),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_889),
.B(n_618),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_871),
.B(n_665),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_838),
.B(n_825),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_848),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_856),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_860),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_849),
.Y(n_959)
);

AND2x2_ASAP7_75t_SL g960 ( 
.A(n_917),
.B(n_670),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_868),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_861),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_900),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_916),
.B(n_670),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_845),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_897),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_846),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_874),
.B(n_671),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_914),
.B(n_823),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_856),
.B(n_671),
.Y(n_970)
);

AND2x2_ASAP7_75t_SL g971 ( 
.A(n_920),
.B(n_678),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_895),
.B(n_678),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_841),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_901),
.A2(n_663),
.B(n_660),
.Y(n_974)
);

AND2x6_ASAP7_75t_L g975 ( 
.A(n_912),
.B(n_708),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_855),
.B(n_915),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_832),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_878),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_831),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_905),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_855),
.B(n_879),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_905),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_923),
.B(n_710),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_865),
.B(n_710),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_865),
.B(n_719),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_863),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_883),
.B(n_719),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_833),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_836),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_883),
.B(n_721),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_913),
.B(n_866),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_922),
.B(n_721),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_841),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_920),
.B(n_691),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_919),
.B(n_691),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_872),
.B(n_722),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_873),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_882),
.B(n_884),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_870),
.B(n_822),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_842),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_859),
.B(n_697),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_859),
.B(n_697),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_880),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_881),
.B(n_697),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_890),
.B(n_703),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_839),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_902),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_896),
.B(n_703),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_875),
.B(n_822),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_903),
.B(n_703),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_906),
.B(n_707),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_910),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_908),
.B(n_722),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_907),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_909),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_850),
.B(n_580),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_911),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_843),
.B(n_707),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_907),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_877),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_844),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_984),
.B(n_921),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_952),
.B(n_957),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_940),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_964),
.B(n_892),
.Y(n_1025)
);

HB1xp67_ASAP7_75t_L g1026 ( 
.A(n_991),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_964),
.B(n_684),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_984),
.B(n_904),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_968),
.B(n_694),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_930),
.B(n_904),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_986),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_1014),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_1003),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_952),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_985),
.B(n_904),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_SL g1036 ( 
.A(n_971),
.B(n_847),
.Y(n_1036)
);

NAND2x1p5_ASAP7_75t_L g1037 ( 
.A(n_930),
.B(n_635),
.Y(n_1037)
);

AO21x2_ASAP7_75t_L g1038 ( 
.A1(n_943),
.A2(n_723),
.B(n_715),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_1003),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_952),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_986),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_959),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_939),
.B(n_723),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_924),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_SL g1045 ( 
.A(n_971),
.B(n_829),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_966),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_930),
.B(n_869),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_959),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_968),
.B(n_699),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_977),
.B(n_584),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_936),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_1005),
.B(n_918),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_957),
.B(n_95),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_983),
.B(n_928),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_983),
.B(n_707),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_936),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_980),
.B(n_982),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_958),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_939),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_966),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_992),
.B(n_712),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_929),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_985),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_962),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_992),
.B(n_972),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_980),
.B(n_982),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_1014),
.B(n_96),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_972),
.B(n_586),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1000),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1007),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1007),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_1014),
.Y(n_1072)
);

CKINVDCx12_ASAP7_75t_R g1073 ( 
.A(n_999),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1015),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_1014),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_954),
.B(n_712),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_942),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_1006),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_954),
.B(n_712),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_934),
.B(n_713),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_927),
.B(n_713),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_927),
.B(n_713),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1000),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_949),
.B(n_590),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_1008),
.B(n_717),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_942),
.B(n_97),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_926),
.B(n_717),
.Y(n_1087)
);

BUFx5_ASAP7_75t_L g1088 ( 
.A(n_944),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_976),
.B(n_717),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_951),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1015),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_937),
.B(n_734),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_926),
.B(n_734),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_1006),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_945),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1017),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_937),
.B(n_734),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1070),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_1032),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1032),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_1062),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1071),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1062),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1077),
.Y(n_1104)
);

BUFx4_ASAP7_75t_SL g1105 ( 
.A(n_1031),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1074),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_1041),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1077),
.Y(n_1108)
);

BUFx5_ASAP7_75t_L g1109 ( 
.A(n_1086),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1023),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1094),
.Y(n_1111)
);

INVx5_ASAP7_75t_L g1112 ( 
.A(n_1032),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1091),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_1072),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1065),
.B(n_970),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_1046),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1096),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_1072),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_1028),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1072),
.Y(n_1120)
);

BUFx2_ASAP7_75t_SL g1121 ( 
.A(n_1078),
.Y(n_1121)
);

BUFx2_ASAP7_75t_SL g1122 ( 
.A(n_1060),
.Y(n_1122)
);

AND2x2_ASAP7_75t_SL g1123 ( 
.A(n_1086),
.B(n_960),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1090),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1034),
.B(n_942),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_1059),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1075),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1022),
.B(n_970),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1075),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1040),
.B(n_942),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1054),
.A2(n_1021),
.B1(n_935),
.B2(n_1020),
.Y(n_1131)
);

INVx3_ASAP7_75t_SL g1132 ( 
.A(n_1043),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1075),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_1065),
.Y(n_1134)
);

BUFx4_ASAP7_75t_SL g1135 ( 
.A(n_1043),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1044),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_1043),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1030),
.B(n_1021),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1024),
.Y(n_1139)
);

CKINVDCx16_ASAP7_75t_R g1140 ( 
.A(n_1047),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1025),
.B(n_1020),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1058),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1064),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1051),
.Y(n_1144)
);

INVx5_ASAP7_75t_L g1145 ( 
.A(n_1033),
.Y(n_1145)
);

INVx8_ASAP7_75t_L g1146 ( 
.A(n_1067),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1054),
.B(n_931),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1067),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1025),
.A2(n_969),
.B1(n_960),
.B2(n_1016),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1033),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1035),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1039),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1063),
.B(n_925),
.Y(n_1153)
);

BUFx12f_ASAP7_75t_L g1154 ( 
.A(n_1085),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1026),
.Y(n_1155)
);

NAND2x1p5_ASAP7_75t_L g1156 ( 
.A(n_1039),
.B(n_941),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1042),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1048),
.Y(n_1158)
);

CKINVDCx16_ASAP7_75t_R g1159 ( 
.A(n_1047),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1056),
.Y(n_1160)
);

INVx3_ASAP7_75t_SL g1161 ( 
.A(n_1052),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1069),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1061),
.B(n_933),
.Y(n_1163)
);

INVx8_ASAP7_75t_L g1164 ( 
.A(n_1112),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1141),
.A2(n_1045),
.B1(n_1128),
.B2(n_1123),
.Y(n_1165)
);

CKINVDCx6p67_ASAP7_75t_R g1166 ( 
.A(n_1107),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1102),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1102),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1107),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1134),
.B(n_1147),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_SL g1171 ( 
.A1(n_1140),
.A2(n_1036),
.B1(n_1159),
.B2(n_1009),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1139),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1134),
.B(n_1027),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1112),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_SL g1175 ( 
.A1(n_1149),
.A2(n_990),
.B(n_987),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1111),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_1103),
.Y(n_1177)
);

CKINVDCx8_ASAP7_75t_R g1178 ( 
.A(n_1121),
.Y(n_1178)
);

CKINVDCx14_ASAP7_75t_R g1179 ( 
.A(n_1126),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1106),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1123),
.A2(n_1131),
.B1(n_1119),
.B2(n_1148),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1131),
.A2(n_990),
.B(n_987),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1148),
.A2(n_978),
.B1(n_963),
.B2(n_1023),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1142),
.Y(n_1184)
);

CKINVDCx6p67_ASAP7_75t_R g1185 ( 
.A(n_1124),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1115),
.A2(n_1036),
.B1(n_991),
.B2(n_1095),
.Y(n_1186)
);

CKINVDCx14_ASAP7_75t_R g1187 ( 
.A(n_1124),
.Y(n_1187)
);

OAI21xp33_ASAP7_75t_L g1188 ( 
.A1(n_1153),
.A2(n_1068),
.B(n_1061),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1146),
.A2(n_978),
.B1(n_1057),
.B2(n_975),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1106),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1146),
.A2(n_1018),
.B1(n_948),
.B2(n_961),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1116),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1146),
.A2(n_948),
.B1(n_961),
.B2(n_951),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_1161),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1138),
.A2(n_1055),
.B1(n_1079),
.B2(n_1076),
.Y(n_1195)
);

BUFx8_ASAP7_75t_L g1196 ( 
.A(n_1155),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1154),
.A2(n_1057),
.B1(n_975),
.B2(n_1084),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1154),
.A2(n_1109),
.B1(n_1153),
.B2(n_1151),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1151),
.A2(n_1081),
.B1(n_1082),
.B2(n_1055),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1143),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1109),
.A2(n_951),
.B1(n_999),
.B2(n_981),
.Y(n_1201)
);

BUFx8_ASAP7_75t_SL g1202 ( 
.A(n_1137),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1098),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1103),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1138),
.A2(n_1076),
.B1(n_1079),
.B2(n_1027),
.Y(n_1205)
);

INVx6_ASAP7_75t_L g1206 ( 
.A(n_1116),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1109),
.A2(n_975),
.B1(n_949),
.B2(n_1053),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1163),
.B(n_933),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1109),
.B(n_947),
.Y(n_1209)
);

BUFx10_ASAP7_75t_L g1210 ( 
.A(n_1101),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1109),
.A2(n_975),
.B1(n_1053),
.B2(n_932),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1161),
.A2(n_1012),
.B1(n_1066),
.B2(n_994),
.Y(n_1212)
);

INVx6_ASAP7_75t_L g1213 ( 
.A(n_1105),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1105),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1113),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1104),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1117),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1136),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1099),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1167),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1172),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1168),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1204),
.B(n_1177),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1188),
.A2(n_953),
.B1(n_947),
.B2(n_950),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1180),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1170),
.B(n_1109),
.Y(n_1226)
);

CKINVDCx11_ASAP7_75t_R g1227 ( 
.A(n_1178),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1184),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1200),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_L g1230 ( 
.A(n_1165),
.B(n_1050),
.C(n_953),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1188),
.A2(n_950),
.B1(n_1080),
.B2(n_995),
.Y(n_1231)
);

BUFx12f_ASAP7_75t_L g1232 ( 
.A(n_1194),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1179),
.B(n_1132),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1201),
.A2(n_1093),
.B1(n_1087),
.B2(n_1110),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1181),
.A2(n_1110),
.B1(n_945),
.B2(n_955),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1213),
.A2(n_1214),
.B1(n_1209),
.B2(n_1208),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1164),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1171),
.B(n_996),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1164),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1190),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1164),
.Y(n_1241)
);

OAI222xp33_ASAP7_75t_L g1242 ( 
.A1(n_1186),
.A2(n_1138),
.B1(n_1080),
.B2(n_1158),
.C1(n_1157),
.C2(n_1160),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1198),
.A2(n_1030),
.B1(n_1130),
.B2(n_1125),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1203),
.Y(n_1244)
);

AOI222xp33_ASAP7_75t_L g1245 ( 
.A1(n_1182),
.A2(n_945),
.B1(n_975),
.B2(n_996),
.C1(n_1013),
.C2(n_1019),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1213),
.A2(n_1092),
.B1(n_1097),
.B2(n_975),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1214),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1215),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1217),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1186),
.A2(n_1130),
.B1(n_1125),
.B2(n_1010),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1193),
.A2(n_1130),
.B1(n_1125),
.B2(n_1011),
.Y(n_1251)
);

INVx5_ASAP7_75t_SL g1252 ( 
.A(n_1166),
.Y(n_1252)
);

OAI21xp33_ASAP7_75t_L g1253 ( 
.A1(n_1183),
.A2(n_1097),
.B(n_1092),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1199),
.A2(n_1038),
.B1(n_1162),
.B2(n_1083),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1210),
.B(n_1013),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1199),
.A2(n_1038),
.B1(n_1144),
.B2(n_1049),
.Y(n_1256)
);

OAI21xp33_ASAP7_75t_L g1257 ( 
.A1(n_1182),
.A2(n_1004),
.B(n_989),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1211),
.A2(n_1122),
.B1(n_938),
.B2(n_946),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1195),
.A2(n_1144),
.B1(n_1029),
.B2(n_1049),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1196),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1195),
.A2(n_1029),
.B1(n_1089),
.B2(n_988),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1169),
.B(n_1129),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1174),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1205),
.A2(n_1089),
.B1(n_974),
.B2(n_500),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1192),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1205),
.A2(n_1089),
.B1(n_500),
.B2(n_956),
.Y(n_1266)
);

BUFx12f_ASAP7_75t_L g1267 ( 
.A(n_1196),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1210),
.B(n_997),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1206),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1218),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1173),
.B(n_998),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1173),
.A2(n_500),
.B1(n_956),
.B2(n_979),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1191),
.A2(n_500),
.B1(n_956),
.B2(n_965),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1176),
.A2(n_944),
.B1(n_946),
.B2(n_1135),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1206),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1212),
.A2(n_1197),
.B1(n_1207),
.B2(n_1189),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1175),
.A2(n_938),
.B1(n_1108),
.B2(n_1104),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1238),
.A2(n_500),
.B1(n_1202),
.B2(n_1187),
.Y(n_1278)
);

OAI211xp5_ASAP7_75t_L g1279 ( 
.A1(n_1224),
.A2(n_1236),
.B(n_1175),
.C(n_1245),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1271),
.B(n_1216),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1236),
.A2(n_1073),
.B1(n_1185),
.B2(n_967),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1224),
.A2(n_956),
.B1(n_1017),
.B2(n_941),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1274),
.A2(n_1219),
.B1(n_1216),
.B2(n_1108),
.Y(n_1283)
);

AOI222xp33_ASAP7_75t_L g1284 ( 
.A1(n_1235),
.A2(n_591),
.B1(n_592),
.B2(n_595),
.C1(n_596),
.C2(n_998),
.Y(n_1284)
);

AOI221xp5_ASAP7_75t_L g1285 ( 
.A1(n_1257),
.A2(n_1231),
.B1(n_1242),
.B2(n_1250),
.C(n_1264),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1276),
.A2(n_941),
.B1(n_993),
.B2(n_1150),
.Y(n_1286)
);

OAI221xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1276),
.A2(n_1135),
.B1(n_1001),
.B2(n_1002),
.C(n_1129),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1226),
.B(n_1114),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1223),
.B(n_1127),
.Y(n_1289)
);

OAI222xp33_ASAP7_75t_L g1290 ( 
.A1(n_1246),
.A2(n_1273),
.B1(n_1258),
.B2(n_1251),
.C1(n_1234),
.C2(n_1243),
.Y(n_1290)
);

AO22x1_ASAP7_75t_L g1291 ( 
.A1(n_1233),
.A2(n_1174),
.B1(n_1133),
.B2(n_1118),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1253),
.A2(n_1152),
.B1(n_1150),
.B2(n_1099),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1246),
.A2(n_1152),
.B1(n_1118),
.B2(n_973),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1220),
.B(n_1100),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1277),
.A2(n_1247),
.B1(n_1255),
.B2(n_1265),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1267),
.A2(n_1088),
.B1(n_973),
.B2(n_1100),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1221),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1222),
.B(n_1225),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1252),
.A2(n_1100),
.B1(n_1120),
.B2(n_1088),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1260),
.A2(n_973),
.B1(n_1120),
.B2(n_1100),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1240),
.B(n_1120),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1261),
.A2(n_1145),
.B1(n_1156),
.B2(n_1037),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1268),
.A2(n_1088),
.B1(n_1145),
.B2(n_1156),
.Y(n_1303)
);

NAND3xp33_ASAP7_75t_SL g1304 ( 
.A(n_1261),
.B(n_1037),
.C(n_668),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1262),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1269),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1254),
.A2(n_1088),
.B1(n_1145),
.B2(n_706),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1254),
.A2(n_1145),
.B(n_651),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1256),
.A2(n_1264),
.B(n_1266),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1256),
.A2(n_1088),
.B1(n_706),
.B2(n_725),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1270),
.B(n_51),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1252),
.A2(n_706),
.B1(n_725),
.B2(n_720),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1227),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1244),
.B(n_1248),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1249),
.Y(n_1316)
);

AOI222xp33_ASAP7_75t_L g1317 ( 
.A1(n_1232),
.A2(n_731),
.B1(n_725),
.B2(n_720),
.C1(n_735),
.C2(n_56),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1266),
.A2(n_731),
.B1(n_735),
.B2(n_675),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1272),
.A2(n_675),
.B1(n_674),
.B2(n_651),
.C(n_643),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1259),
.A2(n_1272),
.B1(n_1252),
.B2(n_1275),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1275),
.A2(n_735),
.B1(n_650),
.B2(n_605),
.Y(n_1321)
);

OAI222xp33_ASAP7_75t_L g1322 ( 
.A1(n_1259),
.A2(n_735),
.B1(n_52),
.B2(n_53),
.C1(n_54),
.C2(n_57),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1239),
.A2(n_650),
.B1(n_636),
.B2(n_652),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1239),
.A2(n_650),
.B1(n_636),
.B2(n_652),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1237),
.A2(n_675),
.B1(n_674),
.B2(n_643),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1237),
.A2(n_1241),
.B1(n_1263),
.B2(n_652),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1230),
.A2(n_636),
.B1(n_629),
.B2(n_59),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1230),
.A2(n_51),
.B1(n_57),
.B2(n_61),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1230),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1220),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1280),
.B(n_63),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1317),
.B(n_629),
.C(n_64),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1328),
.A2(n_64),
.B(n_65),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1287),
.A2(n_629),
.B1(n_66),
.B2(n_67),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1305),
.B(n_65),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1298),
.B(n_66),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1316),
.B(n_68),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1312),
.B(n_68),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1315),
.B(n_69),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1279),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1297),
.B(n_72),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1328),
.B(n_1329),
.C(n_1327),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1329),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_1343)
);

AOI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1322),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.C(n_79),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1278),
.A2(n_1290),
.B(n_1281),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1297),
.B(n_78),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1288),
.B(n_1330),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1309),
.B(n_79),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1285),
.B(n_101),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1289),
.B(n_80),
.Y(n_1350)
);

AND4x1_ASAP7_75t_L g1351 ( 
.A(n_1278),
.B(n_82),
.C(n_83),
.D(n_85),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1295),
.B(n_83),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1311),
.B(n_86),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1301),
.B(n_358),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1309),
.B(n_104),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_SL g1356 ( 
.A1(n_1320),
.A2(n_110),
.B(n_112),
.Y(n_1356)
);

NAND3xp33_ASAP7_75t_L g1357 ( 
.A(n_1284),
.B(n_114),
.C(n_118),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1320),
.A2(n_119),
.B(n_121),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1308),
.B(n_122),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1294),
.B(n_125),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1306),
.B(n_353),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1283),
.B(n_128),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1286),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1300),
.A2(n_1282),
.B1(n_1313),
.B2(n_1293),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1292),
.B(n_136),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1282),
.B(n_1291),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_SL g1367 ( 
.A(n_1314),
.B(n_137),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1326),
.B(n_139),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1308),
.B(n_352),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1303),
.B(n_140),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1307),
.B(n_350),
.Y(n_1371)
);

NAND4xp25_ASAP7_75t_L g1372 ( 
.A(n_1296),
.B(n_148),
.C(n_150),
.D(n_153),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1310),
.B(n_154),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1299),
.B(n_162),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1302),
.B(n_165),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1318),
.B(n_167),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1347),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1332),
.B(n_1357),
.C(n_1349),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1349),
.B(n_1325),
.C(n_1319),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1348),
.B(n_1304),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1331),
.B(n_1323),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1348),
.B(n_182),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1351),
.B(n_1324),
.C(n_1321),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1342),
.A2(n_183),
.B1(n_187),
.B2(n_188),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1341),
.B(n_189),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1350),
.B(n_190),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1346),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1338),
.B(n_192),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1340),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1337),
.B(n_197),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1337),
.B(n_198),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_L g1392 ( 
.A(n_1345),
.B(n_199),
.C(n_205),
.Y(n_1392)
);

AOI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1333),
.A2(n_207),
.B1(n_211),
.B2(n_213),
.C(n_215),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1343),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1355),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1335),
.B(n_220),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1343),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1355),
.B(n_229),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1336),
.B(n_237),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1339),
.B(n_239),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1334),
.B(n_240),
.C(n_243),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1359),
.B(n_245),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1359),
.B(n_246),
.Y(n_1403)
);

OAI211xp5_ASAP7_75t_SL g1404 ( 
.A1(n_1353),
.A2(n_250),
.B(n_251),
.C(n_252),
.Y(n_1404)
);

NAND4xp75_ASAP7_75t_L g1405 ( 
.A(n_1344),
.B(n_255),
.C(n_256),
.D(n_261),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1395),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1395),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1377),
.Y(n_1408)
);

NOR3xp33_ASAP7_75t_L g1409 ( 
.A(n_1378),
.B(n_1356),
.C(n_1358),
.Y(n_1409)
);

NAND4xp75_ASAP7_75t_L g1410 ( 
.A(n_1393),
.B(n_1362),
.C(n_1374),
.D(n_1352),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1387),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1380),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1382),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1382),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1398),
.B(n_1369),
.Y(n_1415)
);

XOR2x2_ASAP7_75t_L g1416 ( 
.A(n_1405),
.B(n_1374),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1402),
.Y(n_1417)
);

XOR2x2_ASAP7_75t_L g1418 ( 
.A(n_1392),
.B(n_1368),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1402),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1399),
.B(n_1366),
.Y(n_1420)
);

NAND4xp75_ASAP7_75t_SL g1421 ( 
.A(n_1381),
.B(n_1375),
.C(n_1370),
.D(n_1371),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1385),
.Y(n_1422)
);

XNOR2xp5_ASAP7_75t_L g1423 ( 
.A(n_1386),
.B(n_1361),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1401),
.A2(n_1368),
.B1(n_1372),
.B2(n_1364),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1408),
.Y(n_1425)
);

XOR2xp5_ASAP7_75t_L g1426 ( 
.A(n_1423),
.B(n_1396),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1409),
.A2(n_1384),
.B1(n_1381),
.B2(n_1389),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1406),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1412),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1411),
.B(n_1402),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1406),
.Y(n_1431)
);

XOR2xp5_ASAP7_75t_L g1432 ( 
.A(n_1423),
.B(n_1390),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1417),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1407),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1413),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1418),
.A2(n_1384),
.B1(n_1404),
.B2(n_1383),
.Y(n_1436)
);

XNOR2x1_ASAP7_75t_L g1437 ( 
.A(n_1432),
.B(n_1416),
.Y(n_1437)
);

OA22x2_ASAP7_75t_L g1438 ( 
.A1(n_1436),
.A2(n_1427),
.B1(n_1426),
.B2(n_1424),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1433),
.Y(n_1439)
);

OA22x2_ASAP7_75t_L g1440 ( 
.A1(n_1429),
.A2(n_1419),
.B1(n_1417),
.B2(n_1422),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1433),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1425),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1430),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1434),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1435),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1428),
.Y(n_1446)
);

OA22x2_ASAP7_75t_L g1447 ( 
.A1(n_1431),
.A2(n_1419),
.B1(n_1417),
.B2(n_1414),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1425),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1425),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1425),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1447),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1442),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1448),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1437),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1439),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1450),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1449),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1440),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1449),
.Y(n_1459)
);

AND4x1_ASAP7_75t_L g1460 ( 
.A(n_1454),
.B(n_1367),
.C(n_1438),
.D(n_1394),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1458),
.A2(n_1410),
.B1(n_1443),
.B2(n_1444),
.Y(n_1461)
);

OA22x2_ASAP7_75t_L g1462 ( 
.A1(n_1451),
.A2(n_1455),
.B1(n_1441),
.B2(n_1452),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1456),
.Y(n_1463)
);

OAI322xp33_ASAP7_75t_L g1464 ( 
.A1(n_1451),
.A2(n_1450),
.A3(n_1445),
.B1(n_1446),
.B2(n_1420),
.C1(n_1388),
.C2(n_1400),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1461),
.A2(n_1459),
.B1(n_1457),
.B2(n_1453),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1464),
.A2(n_1394),
.B1(n_1397),
.B2(n_1379),
.C(n_1413),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1462),
.Y(n_1467)
);

AOI22x1_ASAP7_75t_L g1468 ( 
.A1(n_1460),
.A2(n_1403),
.B1(n_1391),
.B2(n_1414),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1465),
.A2(n_1463),
.B1(n_1403),
.B2(n_1415),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1467),
.A2(n_1466),
.B1(n_1468),
.B2(n_1403),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1465),
.A2(n_1354),
.B1(n_1376),
.B2(n_1365),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1467),
.B(n_1360),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1465),
.A2(n_1363),
.B(n_1376),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1472),
.B(n_1373),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1470),
.Y(n_1475)
);

AO22x1_ASAP7_75t_L g1476 ( 
.A1(n_1473),
.A2(n_1421),
.B1(n_1363),
.B2(n_273),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1469),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1471),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1474),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1477),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1475),
.B(n_271),
.Y(n_1481)
);

NAND2x1_ASAP7_75t_L g1482 ( 
.A(n_1478),
.B(n_1476),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1480),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1479),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1481),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1485),
.A2(n_1482),
.B1(n_285),
.B2(n_286),
.Y(n_1486)
);

NOR4xp25_ASAP7_75t_L g1487 ( 
.A(n_1484),
.B(n_284),
.C(n_288),
.D(n_291),
.Y(n_1487)
);

AOI211xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1483),
.A2(n_299),
.B(n_301),
.C(n_305),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1486),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1489),
.A2(n_1487),
.B1(n_1488),
.B2(n_314),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1490),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1491),
.A2(n_315),
.B1(n_319),
.B2(n_320),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1492),
.Y(n_1493)
);

AOI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1493),
.A2(n_1491),
.B1(n_326),
.B2(n_327),
.C(n_329),
.Y(n_1494)
);

AOI211xp5_ASAP7_75t_L g1495 ( 
.A1(n_1494),
.A2(n_334),
.B(n_335),
.C(n_336),
.Y(n_1495)
);


endmodule