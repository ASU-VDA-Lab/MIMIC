module fake_aes_3728_n_526 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_526);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_526;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_25), .Y(n_76) );
CKINVDCx16_ASAP7_75t_R g77 ( .A(n_50), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_74), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_51), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_32), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_21), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_48), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_72), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_36), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_49), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_58), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_40), .Y(n_87) );
BUFx2_ASAP7_75t_L g88 ( .A(n_13), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_39), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_4), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_56), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_10), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_24), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_13), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_63), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_43), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_4), .Y(n_98) );
OR2x2_ASAP7_75t_L g99 ( .A(n_64), .B(n_12), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_29), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_35), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_52), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_65), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_57), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_68), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_17), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_7), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_42), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_12), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_103), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_103), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_88), .B(n_0), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_78), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_88), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_78), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_104), .B(n_0), .Y(n_118) );
AND2x6_ASAP7_75t_L g119 ( .A(n_79), .B(n_33), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_104), .B(n_1), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_95), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_79), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
CKINVDCx6p67_ASAP7_75t_R g124 ( .A(n_77), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_95), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_80), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_96), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_93), .B(n_1), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_112), .Y(n_135) );
INVx4_ASAP7_75t_SL g136 ( .A(n_119), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_125), .B(n_98), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g138 ( .A(n_129), .B(n_99), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_119), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_124), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_115), .B(n_97), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
INVx2_ASAP7_75t_SL g143 ( .A(n_115), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_133), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_123), .B(n_101), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_124), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_133), .Y(n_147) );
OR2x2_ASAP7_75t_L g148 ( .A(n_114), .B(n_111), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_123), .B(n_98), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_126), .B(n_84), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_113), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_126), .A2(n_110), .B1(n_91), .B2(n_107), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_130), .B(n_82), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_130), .B(n_90), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_113), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_133), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_143), .B(n_131), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_142), .B(n_129), .Y(n_160) );
NOR2x2_ASAP7_75t_L g161 ( .A(n_140), .B(n_116), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_148), .B(n_127), .Y(n_162) );
NAND2xp33_ASAP7_75t_L g163 ( .A(n_143), .B(n_119), .Y(n_163) );
AND3x1_ASAP7_75t_L g164 ( .A(n_152), .B(n_120), .C(n_118), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_149), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_145), .A2(n_119), .B1(n_132), .B2(n_131), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_146), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_139), .B(n_127), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_145), .B(n_132), .Y(n_172) );
NOR2xp33_ASAP7_75t_R g173 ( .A(n_148), .B(n_76), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g174 ( .A1(n_138), .A2(n_91), .B1(n_110), .B2(n_107), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_138), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_135), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_139), .A2(n_117), .B(n_122), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_149), .A2(n_119), .B1(n_121), .B2(n_122), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_149), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_139), .B(n_87), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
NOR2x2_ASAP7_75t_L g185 ( .A(n_138), .B(n_108), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_137), .B(n_117), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_137), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_137), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_186), .B(n_138), .Y(n_190) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
NOR2xp33_ASAP7_75t_SL g192 ( .A(n_168), .B(n_139), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_165), .Y(n_193) );
BUFx4f_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_172), .A2(n_141), .B(n_153), .C(n_154), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_186), .B(n_137), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_175), .B(n_150), .Y(n_197) );
NOR2xp67_ASAP7_75t_L g198 ( .A(n_162), .B(n_153), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_160), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_166), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_181), .B(n_155), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_164), .A2(n_155), .B1(n_152), .B2(n_154), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_164), .A2(n_155), .B1(n_149), .B2(n_141), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_173), .B(n_151), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_166), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_181), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_187), .B(n_155), .Y(n_208) );
O2A1O1Ixp5_ASAP7_75t_SL g209 ( .A1(n_171), .A2(n_128), .B(n_109), .C(n_85), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_186), .B(n_156), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_160), .Y(n_211) );
NAND2x1p5_ASAP7_75t_L g212 ( .A(n_166), .B(n_156), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_188), .B(n_99), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_166), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_186), .B(n_169), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_185), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_163), .A2(n_136), .B(n_85), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_174), .A2(n_136), .B1(n_83), .B2(n_90), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_174), .A2(n_136), .B1(n_83), .B2(n_106), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_169), .B(n_136), .Y(n_220) );
OAI22xp5_ASAP7_75t_SL g221 ( .A1(n_216), .A2(n_161), .B1(n_180), .B2(n_167), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_193), .B(n_169), .Y(n_222) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_209), .A2(n_180), .B(n_179), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_193), .B(n_169), .Y(n_224) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_217), .A2(n_159), .B(n_158), .Y(n_225) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_203), .A2(n_109), .B(n_89), .Y(n_226) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_202), .A2(n_158), .B(n_184), .Y(n_227) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_195), .A2(n_158), .B(n_184), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_206), .Y(n_229) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_218), .A2(n_89), .B(n_105), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_206), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_190), .A2(n_182), .B1(n_160), .B2(n_171), .Y(n_232) );
AO31x2_ASAP7_75t_L g233 ( .A1(n_213), .A2(n_177), .A3(n_178), .B(n_165), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_191), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_201), .A2(n_177), .B(n_178), .Y(n_236) );
NOR2xp67_ASAP7_75t_L g237 ( .A(n_199), .B(n_219), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_205), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_214), .Y(n_239) );
NAND3xp33_ASAP7_75t_L g240 ( .A(n_213), .B(n_133), .C(n_106), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_201), .A2(n_183), .B(n_105), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_198), .A2(n_170), .B(n_181), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_191), .B(n_182), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_204), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_212), .A2(n_182), .B(n_147), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_199), .B(n_182), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_231), .Y(n_247) );
AOI222xp33_ASAP7_75t_L g248 ( .A1(n_221), .A2(n_196), .B1(n_215), .B2(n_197), .C1(n_108), .C2(n_210), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_233), .B(n_197), .Y(n_249) );
AND2x4_ASAP7_75t_SL g250 ( .A(n_234), .B(n_199), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_221), .A2(n_211), .B1(n_194), .B2(n_160), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_231), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_244), .A2(n_211), .B1(n_194), .B2(n_160), .Y(n_253) );
OAI22xp33_ASAP7_75t_SL g254 ( .A1(n_229), .A2(n_194), .B1(n_192), .B2(n_212), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_229), .A2(n_220), .B(n_189), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_243), .A2(n_208), .B1(n_160), .B2(n_220), .Y(n_256) );
INVx6_ASAP7_75t_L g257 ( .A(n_246), .Y(n_257) );
OAI221xp5_ASAP7_75t_L g258 ( .A1(n_240), .A2(n_208), .B1(n_207), .B2(n_189), .C(n_86), .Y(n_258) );
AOI22xp33_ASAP7_75t_SL g259 ( .A1(n_243), .A2(n_226), .B1(n_230), .B2(n_240), .Y(n_259) );
OAI221xp5_ASAP7_75t_L g260 ( .A1(n_232), .A2(n_207), .B1(n_189), .B2(n_86), .C(n_176), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_237), .A2(n_160), .B1(n_207), .B2(n_176), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_237), .A2(n_207), .B1(n_176), .B2(n_86), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_243), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_226), .A2(n_176), .B1(n_86), .B2(n_100), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_229), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_232), .A2(n_92), .B1(n_94), .B2(n_102), .Y(n_267) );
NOR2xp67_ASAP7_75t_L g268 ( .A(n_252), .B(n_235), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_247), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_265), .B(n_233), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_265), .B(n_233), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_249), .B(n_233), .Y(n_272) );
BUFx2_ASAP7_75t_SL g273 ( .A(n_247), .Y(n_273) );
AOI222xp33_ASAP7_75t_L g274 ( .A1(n_251), .A2(n_238), .B1(n_222), .B2(n_224), .C1(n_246), .C2(n_239), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_266), .B(n_233), .Y(n_275) );
INVx4_ASAP7_75t_R g276 ( .A(n_250), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_259), .B(n_233), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_257), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_257), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_257), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_257), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_263), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_261), .B(n_236), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_248), .B(n_233), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_263), .B(n_226), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_250), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_264), .B(n_226), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_256), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_270), .B(n_227), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_268), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_270), .B(n_227), .Y(n_291) );
OAI33xp33_ASAP7_75t_L g292 ( .A1(n_269), .A2(n_267), .A3(n_238), .B1(n_254), .B2(n_224), .B3(n_222), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_270), .Y(n_293) );
OAI321xp33_ASAP7_75t_L g294 ( .A1(n_277), .A2(n_262), .A3(n_260), .B1(n_258), .B2(n_253), .C(n_133), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_271), .B(n_227), .Y(n_295) );
OR2x6_ASAP7_75t_L g296 ( .A(n_273), .B(n_228), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_269), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
AOI21xp5_ASAP7_75t_SL g299 ( .A1(n_272), .A2(n_230), .B(n_255), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_276), .Y(n_300) );
AOI22xp33_ASAP7_75t_SL g301 ( .A1(n_273), .A2(n_230), .B1(n_228), .B2(n_239), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_275), .B(n_230), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_283), .B(n_236), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_275), .B(n_236), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_272), .B(n_228), .Y(n_306) );
OAI31xp33_ASAP7_75t_L g307 ( .A1(n_284), .A2(n_246), .A3(n_239), .B(n_242), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_275), .B(n_246), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_277), .B(n_245), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_284), .A2(n_246), .B1(n_242), .B2(n_223), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_272), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_277), .B(n_285), .Y(n_312) );
NOR3xp33_ASAP7_75t_L g313 ( .A(n_278), .B(n_223), .C(n_241), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_268), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_283), .Y(n_316) );
NAND4xp25_ASAP7_75t_L g317 ( .A(n_274), .B(n_2), .C(n_3), .D(n_5), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_298), .B(n_283), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_297), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_298), .B(n_283), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_298), .B(n_288), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_311), .B(n_288), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_302), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_312), .B(n_285), .Y(n_328) );
INVx5_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_289), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_311), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_312), .B(n_285), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_311), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_309), .B(n_287), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_296), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_306), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_306), .B(n_284), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_314), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_316), .B(n_279), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_303), .B(n_282), .Y(n_343) );
NAND2xp33_ASAP7_75t_SL g344 ( .A(n_300), .B(n_282), .Y(n_344) );
NAND3xp33_ASAP7_75t_SL g345 ( .A(n_301), .B(n_274), .C(n_287), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_305), .B(n_287), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_305), .B(n_279), .Y(n_347) );
NOR2x1_ASAP7_75t_L g348 ( .A(n_317), .B(n_278), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_289), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_309), .B(n_279), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_291), .B(n_281), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_289), .B(n_281), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_291), .B(n_280), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_300), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_295), .B(n_280), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_296), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_289), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_295), .B(n_280), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_316), .B(n_223), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_307), .A2(n_286), .B1(n_241), .B2(n_245), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
NOR2xp33_ASAP7_75t_SL g362 ( .A(n_354), .B(n_286), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_344), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_320), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_343), .B(n_308), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_349), .B(n_315), .Y(n_366) );
OR2x6_ASAP7_75t_L g367 ( .A(n_319), .B(n_296), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_343), .B(n_315), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_340), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_348), .B(n_292), .Y(n_370) );
AOI211x1_ASAP7_75t_L g371 ( .A1(n_345), .A2(n_307), .B(n_3), .C(n_5), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_329), .B(n_304), .Y(n_372) );
OR2x6_ASAP7_75t_L g373 ( .A(n_319), .B(n_299), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_328), .B(n_310), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_340), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_341), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_333), .B(n_304), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_351), .B(n_304), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_349), .B(n_304), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_338), .B(n_310), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_358), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_338), .B(n_299), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_357), .B(n_313), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_357), .B(n_2), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_318), .B(n_6), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_335), .B(n_286), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_341), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_358), .B(n_6), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_322), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_351), .B(n_7), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_322), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_318), .B(n_8), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_324), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_335), .B(n_9), .Y(n_394) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_337), .B(n_276), .Y(n_395) );
NOR2x1_ASAP7_75t_L g396 ( .A(n_336), .B(n_294), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_326), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_347), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_360), .B(n_144), .C(n_147), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_324), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_330), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_330), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_339), .B(n_9), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_321), .B(n_10), .Y(n_404) );
XOR2xp5_ASAP7_75t_L g405 ( .A(n_352), .B(n_11), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_347), .Y(n_406) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_336), .B(n_241), .C(n_245), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_346), .B(n_11), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_339), .B(n_14), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_323), .B(n_14), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_326), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_369), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_370), .A2(n_346), .B(n_356), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_376), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_379), .B(n_331), .Y(n_416) );
OAI22xp33_ASAP7_75t_SL g417 ( .A1(n_363), .A2(n_329), .B1(n_337), .B2(n_336), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_395), .A2(n_329), .B1(n_356), .B2(n_352), .Y(n_418) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_370), .A2(n_331), .B(n_355), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_374), .B(n_323), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_361), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_398), .B(n_325), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_364), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_405), .A2(n_355), .B1(n_353), .B2(n_329), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_406), .B(n_353), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_381), .B(n_327), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_389), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g431 ( .A1(n_403), .A2(n_332), .B(n_334), .C(n_327), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_402), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_395), .A2(n_329), .B1(n_325), .B2(n_334), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_368), .B(n_350), .Y(n_435) );
OAI32xp33_ASAP7_75t_L g436 ( .A1(n_408), .A2(n_332), .A3(n_321), .B1(n_350), .B2(n_359), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_385), .B(n_359), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_371), .A2(n_329), .B1(n_342), .B2(n_17), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_387), .Y(n_439) );
OAI321xp33_ASAP7_75t_L g440 ( .A1(n_373), .A2(n_342), .A3(n_16), .B1(n_18), .B2(n_19), .C(n_15), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_396), .A2(n_342), .B(n_225), .Y(n_441) );
AOI332xp33_ASAP7_75t_L g442 ( .A1(n_409), .A2(n_15), .A3(n_16), .B1(n_18), .B2(n_19), .B3(n_157), .C1(n_147), .C2(n_144), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_385), .B(n_225), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_411), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_365), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_379), .B(n_20), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_389), .Y(n_447) );
NAND2xp33_ASAP7_75t_SL g448 ( .A(n_392), .B(n_22), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_392), .B(n_225), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_391), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_397), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_391), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_394), .B(n_23), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_378), .B(n_26), .Y(n_454) );
OAI21xp5_ASAP7_75t_SL g455 ( .A1(n_404), .A2(n_27), .B(n_28), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_431), .B(n_383), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_412), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_416), .B(n_383), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_413), .Y(n_459) );
INVxp67_ASAP7_75t_SL g460 ( .A(n_451), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_415), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_436), .A2(n_382), .B1(n_390), .B2(n_404), .C(n_410), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_421), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_420), .B(n_380), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_451), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_425), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_417), .B(n_362), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_422), .Y(n_469) );
XOR2x2_ASAP7_75t_L g470 ( .A(n_424), .B(n_388), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_416), .B(n_366), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_414), .B(n_372), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_430), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_445), .B(n_366), .Y(n_474) );
OAI222xp33_ASAP7_75t_L g475 ( .A1(n_424), .A2(n_373), .B1(n_367), .B2(n_377), .C1(n_386), .C2(n_384), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_427), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_435), .B(n_373), .Y(n_477) );
AOI222xp33_ASAP7_75t_L g478 ( .A1(n_438), .A2(n_384), .B1(n_372), .B2(n_397), .C1(n_399), .C2(n_367), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g479 ( .A1(n_419), .A2(n_372), .B1(n_367), .B2(n_407), .C1(n_157), .C2(n_144), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_432), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_437), .B(n_407), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_444), .B(n_31), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_430), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_468), .B(n_418), .Y(n_485) );
AOI21xp33_ASAP7_75t_SL g486 ( .A1(n_468), .A2(n_455), .B(n_433), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_477), .B(n_434), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_472), .A2(n_448), .B(n_440), .Y(n_488) );
AOI32xp33_ASAP7_75t_L g489 ( .A1(n_462), .A2(n_448), .A3(n_439), .B1(n_446), .B2(n_454), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_472), .A2(n_426), .B(n_441), .C(n_429), .Y(n_490) );
OAI21xp5_ASAP7_75t_SL g491 ( .A1(n_478), .A2(n_446), .B(n_453), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_456), .B(n_452), .Y(n_492) );
INVxp67_ASAP7_75t_SL g493 ( .A(n_460), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_470), .A2(n_453), .B1(n_449), .B2(n_443), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_469), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_469), .A2(n_450), .B1(n_447), .B2(n_442), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_470), .A2(n_157), .B1(n_37), .B2(n_38), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_479), .B(n_34), .C(n_41), .D(n_44), .Y(n_498) );
AOI322xp5_ASAP7_75t_L g499 ( .A1(n_458), .A2(n_45), .A3(n_46), .B1(n_47), .B2(n_53), .C1(n_54), .C2(n_55), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_475), .A2(n_59), .B(n_60), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g501 ( .A1(n_482), .A2(n_61), .B1(n_62), .B2(n_66), .C1(n_69), .C2(n_70), .Y(n_501) );
AOI311xp33_ASAP7_75t_L g502 ( .A1(n_496), .A2(n_464), .A3(n_481), .B(n_480), .C(n_476), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_490), .A2(n_466), .B1(n_463), .B2(n_467), .C(n_457), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_485), .A2(n_461), .B1(n_459), .B2(n_477), .C(n_458), .Y(n_504) );
AOI21xp33_ASAP7_75t_L g505 ( .A1(n_497), .A2(n_483), .B(n_465), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_492), .B(n_474), .Y(n_506) );
AOI211xp5_ASAP7_75t_L g507 ( .A1(n_486), .A2(n_474), .B(n_465), .C(n_484), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_489), .A2(n_473), .B1(n_484), .B2(n_471), .C(n_75), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_487), .Y(n_509) );
NAND4xp75_ASAP7_75t_L g510 ( .A(n_488), .B(n_471), .C(n_473), .D(n_73), .Y(n_510) );
NOR3x2_ASAP7_75t_L g511 ( .A(n_510), .B(n_501), .C(n_498), .Y(n_511) );
BUFx2_ASAP7_75t_L g512 ( .A(n_509), .Y(n_512) );
BUFx12f_ASAP7_75t_L g513 ( .A(n_509), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_507), .A2(n_491), .B(n_500), .C(n_494), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_502), .B(n_495), .Y(n_515) );
AND5x1_ASAP7_75t_L g516 ( .A(n_514), .B(n_508), .C(n_504), .D(n_503), .E(n_499), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_515), .B(n_505), .C(n_493), .Y(n_517) );
NOR2x1_ASAP7_75t_L g518 ( .A(n_512), .B(n_506), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_518), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_517), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g521 ( .A1(n_520), .A2(n_513), .B1(n_516), .B2(n_511), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_519), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_522), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_523), .Y(n_524) );
XNOR2x1_ASAP7_75t_L g525 ( .A(n_524), .B(n_521), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_525), .A2(n_493), .B(n_71), .Y(n_526) );
endmodule