module real_jpeg_19194_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_281, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_281;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_278;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_0),
.A2(n_3),
.B1(n_18),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_61),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_0),
.A2(n_5),
.B1(n_61),
.B2(n_72),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_1),
.A2(n_3),
.B1(n_17),
.B2(n_18),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_1),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_1),
.A2(n_17),
.B1(n_46),
.B2(n_47),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_1),
.A2(n_5),
.B1(n_17),
.B2(n_72),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_3),
.B1(n_18),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_5),
.B1(n_57),
.B2(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_57),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_22),
.B(n_26),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_2),
.B(n_33),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_2),
.B(n_44),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_SL g170 ( 
.A1(n_2),
.A2(n_47),
.B(n_48),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_3),
.A2(n_7),
.B1(n_18),
.B2(n_31),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_23),
.B(n_57),
.C(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_4),
.Y(n_92)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_4),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_10),
.B1(n_70),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_7),
.B1(n_31),
.B2(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_5),
.B(n_99),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_7),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_225)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_18),
.B(n_21),
.C(n_24),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_10),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_36),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_34),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_27),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_19),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_19),
.B(n_62),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_24),
.Y(n_19)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_30),
.B(n_54),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_25),
.A2(n_45),
.B(n_48),
.C(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_48),
.Y(n_52)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_26),
.A2(n_49),
.B(n_57),
.C(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_28),
.B(n_38),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_33),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_33),
.A2(n_55),
.B(n_60),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_74),
.B(n_279),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_39),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_39),
.B(n_277),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_53),
.CI(n_58),
.CON(n_39),
.SN(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_44),
.B1(n_50),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_43),
.B(n_104),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_45),
.A2(n_51),
.B1(n_104),
.B2(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_45),
.A2(n_256),
.B(n_257),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_47),
.A2(n_57),
.B(n_70),
.C(n_146),
.Y(n_145)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_57),
.B(n_92),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_57),
.B(n_71),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_65),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_59),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_59),
.B(n_113),
.C(n_114),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_59),
.A2(n_101),
.B1(n_112),
.B2(n_125),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_59),
.B(n_101),
.C(n_220),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_59),
.A2(n_112),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_63),
.A2(n_65),
.B1(n_254),
.B2(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_63),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_64),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_65),
.A2(n_254),
.B1(n_255),
.B2(n_258),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_65),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_73),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_68),
.A2(n_71),
.B1(n_86),
.B2(n_89),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_71),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_72),
.B(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_276),
.B(n_278),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_249),
.A3(n_269),
.B1(n_274),
.B2(n_275),
.C(n_281),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_233),
.B(n_248),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_214),
.B(n_232),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_135),
.B(n_195),
.C(n_213),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_120),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_80),
.B(n_120),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_108),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_100),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_82),
.B(n_100),
.C(n_108),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_90),
.B2(n_91),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_84),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_83),
.A2(n_84),
.B1(n_101),
.B2(n_125),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_83),
.B(n_91),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_84),
.B(n_145),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_84),
.B(n_101),
.C(n_168),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_88),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_88),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_92),
.B(n_98),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_119),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_95),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_107),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_101),
.A2(n_105),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_103),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_122),
.B1(n_123),
.B2(n_126),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_107),
.A2(n_122),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_107),
.B(n_207),
.C(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_107),
.A2(n_122),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_107),
.A2(n_122),
.B1(n_263),
.B2(n_267),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_110),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_130),
.C(n_132),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_110),
.A2(n_113),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_110),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_110),
.B(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_152),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_128),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_160),
.C(n_163),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.C(n_129),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_121),
.B(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_122),
.B(n_254),
.C(n_258),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_122),
.B(n_267),
.C(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_129),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_142),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_194),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_189),
.B(n_193),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_177),
.B(n_188),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_165),
.B(n_176),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_155),
.B(n_164),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_147),
.B(n_154),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_151),
.B(n_153),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_157),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_163),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_163),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_180),
.C(n_187),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_163),
.B(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_167),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_169),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_174),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_197),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_211),
.B2(n_212),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_206),
.C(n_212),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_211),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_216),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_231),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_223),
.C(n_231),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_228),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_228),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_243),
.B(n_245),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_235),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_246),
.B2(n_247),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_241),
.C(n_247),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_251),
.C(n_259),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_251),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_243),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_261),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_255),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_260),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_268),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);


endmodule