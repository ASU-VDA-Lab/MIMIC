module real_jpeg_13703_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_249;
wire n_83;
wire n_166;
wire n_286;
wire n_221;
wire n_176;
wire n_215;
wire n_292;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_200;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_202;
wire n_213;
wire n_128;
wire n_179;
wire n_167;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_68),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_3),
.A2(n_29),
.B1(n_35),
.B2(n_68),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_4),
.A2(n_29),
.B1(n_35),
.B2(n_70),
.Y(n_202)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_6),
.A2(n_64),
.B1(n_65),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_6),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_6),
.A2(n_59),
.B1(n_62),
.B2(n_148),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_148),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_148),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_59),
.B1(n_62),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_7),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_29),
.B1(n_35),
.B2(n_78),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_8),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_8),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_12),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_12),
.A2(n_59),
.B1(n_62),
.B2(n_101),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_101),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_101),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_13),
.A2(n_52),
.B1(n_59),
.B2(n_62),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_14),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_14),
.A2(n_64),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_14),
.B(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_14),
.B(n_62),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_140),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_14),
.A2(n_43),
.B(n_48),
.C(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_14),
.B(n_109),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_14),
.B(n_32),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_53),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_14),
.A2(n_62),
.B(n_199),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_15),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_15),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_15),
.A2(n_36),
.B1(n_59),
.B2(n_62),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_16),
.A2(n_45),
.B1(n_59),
.B2(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_16),
.A2(n_29),
.B1(n_35),
.B2(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_16),
.A2(n_45),
.B1(n_64),
.B2(n_65),
.Y(n_280)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_271),
.B1(n_293),
.B2(n_294),
.Y(n_19)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_124),
.B(n_270),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_22),
.B(n_102),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.C(n_86),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_23),
.B(n_80),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_56),
.C(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_28),
.A2(n_32),
.B(n_37),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_28),
.A2(n_32),
.B1(n_92),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_28),
.A2(n_32),
.B1(n_136),
.B2(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_28),
.A2(n_32),
.B1(n_178),
.B2(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_28),
.A2(n_32),
.B1(n_202),
.B2(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_28),
.A2(n_32),
.B1(n_140),
.B2(n_235),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_28),
.A2(n_32),
.B1(n_228),
.B2(n_235),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_29),
.B(n_237),
.Y(n_236)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_31),
.A2(n_34),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_31),
.A2(n_90),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_35),
.A2(n_49),
.B(n_140),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_42),
.A2(n_50),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_44),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_43),
.B(n_74),
.Y(n_200)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_44),
.A2(n_62),
.A3(n_75),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_46),
.A2(n_53),
.B1(n_84),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_46),
.A2(n_53),
.B1(n_95),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_46),
.A2(n_53),
.B1(n_166),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_46),
.A2(n_53),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_46),
.A2(n_53),
.B1(n_214),
.B2(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_46),
.A2(n_53),
.B(n_111),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_50),
.A2(n_96),
.B1(n_193),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_57),
.A2(n_58),
.B1(n_147),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_57),
.A2(n_58),
.B1(n_120),
.B2(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_58),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_59),
.A2(n_61),
.A3(n_64),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_62),
.Y(n_138)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_65),
.B(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_72),
.A2(n_73),
.B1(n_143),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_72),
.A2(n_73),
.B1(n_174),
.B2(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_73),
.Y(n_109)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_85),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_82),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_82),
.A2(n_119),
.B(n_121),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_88),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_89),
.B(n_93),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_99),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_123),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_110),
.B(n_112),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_109),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_107),
.A2(n_109),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_112),
.A2(n_277),
.B1(n_289),
.B2(n_290),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_112),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_113),
.B(n_122),
.C(n_123),
.Y(n_291)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_154),
.B(n_269),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_152),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_126),
.B(n_152),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_132),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_127),
.A2(n_128),
.B1(n_131),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_131),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_132),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.C(n_145),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_145),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_185),
.B(n_263),
.C(n_268),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_179),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_156),
.B(n_179),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_169),
.C(n_171),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_157),
.A2(n_158),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_163),
.C(n_168),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_169),
.B(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_177),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_172),
.B(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_181),
.B(n_182),
.C(n_183),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_262),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_206),
.B(n_261),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_203),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_188),
.B(n_203),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_194),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_189),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_191),
.A2(n_194),
.B1(n_195),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_255),
.B(n_260),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_244),
.B(n_254),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_224),
.B(n_243),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_210),
.B(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_220),
.C(n_222),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_242),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_230),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_241),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_246),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_250),
.C(n_252),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_292),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_291),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_291),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_288),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_283),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);


endmodule