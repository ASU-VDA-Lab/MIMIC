module real_jpeg_11724_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_296, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_296;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_184;
wire n_200;
wire n_275;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_270;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_4),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_148),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_148),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_148),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_6),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_57),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_67),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_67),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_10),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_82),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_82),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_11),
.B(n_43),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_12),
.B(n_29),
.C(n_62),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_12),
.B(n_80),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_12),
.A2(n_92),
.B(n_152),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_12),
.A2(n_42),
.B(n_79),
.C(n_179),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_136),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_12),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_12),
.B(n_38),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_13),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_40),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_13),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_51),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_51),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_15),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_101),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_101),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_101),
.Y(n_227)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_123),
.B1(n_293),
.B2(n_294),
.Y(n_18)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_19),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_104),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_21),
.B(n_104),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_70),
.C(n_86),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_22),
.A2(n_23),
.B1(n_70),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_53),
.B2(n_69),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B1(n_36),
.B2(n_52),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_26),
.A2(n_36),
.B(n_69),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_26),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_31),
.B(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_27),
.A2(n_31),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_27),
.B(n_153),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_27),
.A2(n_31),
.B1(n_91),
.B2(n_241),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_28),
.A2(n_29),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_28),
.B(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_31),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_31),
.B(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_33),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_39),
.A2(n_47),
.B(n_136),
.C(n_223),
.Y(n_222)
);

AOI32xp33_ASAP7_75t_L g236 ( 
.A1(n_39),
.A2(n_42),
.A3(n_44),
.B1(n_224),
.B2(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_41),
.B(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_41),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_41),
.A2(n_45),
.B(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_41),
.A2(n_47),
.B1(n_100),
.B2(n_251),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_42),
.A2(n_43),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_47),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B1(n_65),
.B2(n_68),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_60),
.B1(n_68),
.B2(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_59),
.B1(n_78),
.B2(n_79),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_58),
.B(n_140),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_59),
.A2(n_78),
.B(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_68),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_60),
.B(n_138),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_60),
.A2(n_68),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_60),
.A2(n_68),
.B1(n_96),
.B2(n_230),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_64),
.A2(n_147),
.B(n_149),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_64),
.B(n_136),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_64),
.A2(n_149),
.B(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_70),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B(n_85),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_74),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_72),
.A2(n_135),
.B(n_137),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_72),
.A2(n_137),
.B(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_81),
.B1(n_83),
.B2(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_75),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_75),
.A2(n_83),
.B1(n_199),
.B2(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_75),
.A2(n_185),
.B(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_80),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_76),
.B(n_186),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_80),
.B(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_83),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_83),
.A2(n_98),
.B(n_200),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_86),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.C(n_99),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_87),
.A2(n_88),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_89),
.A2(n_94),
.B1(n_95),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_89),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_92),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_92),
.A2(n_93),
.B1(n_181),
.B2(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_92),
.A2(n_93),
.B1(n_207),
.B2(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_93),
.A2(n_158),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_93),
.B(n_136),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_93),
.A2(n_166),
.B(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_97),
.B(n_99),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_103),
.B(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B1(n_114),
.B2(n_116),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_123),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_287),
.B(n_292),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_275),
.B(n_286),
.Y(n_125)
);

OAI321xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_243),
.A3(n_268),
.B1(n_273),
.B2(n_274),
.C(n_296),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_216),
.B(n_242),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_193),
.B(n_215),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_174),
.B(n_192),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_154),
.B(n_173),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_132),
.B(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_139),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_134),
.B1(n_139),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_150),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_146),
.C(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_162),
.B(n_172),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_160),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_167),
.B(n_171),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_164),
.B(n_165),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_176),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_187),
.C(n_191),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_180),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_195),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_208),
.B2(n_209),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_211),
.C(n_213),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_202),
.C(n_206),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_218),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_232),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_219),
.B(n_233),
.C(n_234),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_231),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_226),
.C(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_258),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_258),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.C(n_257),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_245),
.A2(n_246),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_253),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_252),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_252),
.C(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_254),
.B(n_257),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_256),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_267),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_262),
.C(n_267),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_285),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_285),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);


endmodule