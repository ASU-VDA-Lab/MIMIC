module fake_jpeg_15037_n_258 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_258);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_27),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_44),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_17),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_16),
.B1(n_20),
.B2(n_18),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx9p33_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_23),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_69),
.B1(n_42),
.B2(n_48),
.Y(n_75)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_16),
.B1(n_15),
.B2(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_21),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_40),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_51),
.B1(n_49),
.B2(n_43),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_81),
.B1(n_89),
.B2(n_70),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_75),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_53),
.B1(n_72),
.B2(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_77),
.B1(n_90),
.B2(n_63),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_40),
.B1(n_48),
.B2(n_39),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_39),
.B1(n_33),
.B2(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_17),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_28),
.B1(n_37),
.B2(n_43),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_36),
.C(n_24),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_62),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_102),
.B1(n_56),
.B2(n_74),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_56),
.B1(n_69),
.B2(n_66),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_56),
.B1(n_66),
.B2(n_86),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_104),
.Y(n_128)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_100),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_0),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_67),
.B1(n_65),
.B2(n_68),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_108),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_55),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_109),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_55),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_78),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_93),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_85),
.B(n_84),
.C(n_83),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_123),
.B(n_124),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_78),
.B1(n_81),
.B2(n_89),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_74),
.B1(n_97),
.B2(n_49),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_122),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_92),
.C(n_55),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_125),
.C(n_127),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_94),
.C(n_101),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_79),
.B(n_15),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_79),
.B(n_22),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_55),
.C(n_74),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_132),
.B(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_99),
.B(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_97),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_104),
.B(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_149),
.B1(n_117),
.B2(n_116),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_110),
.B(n_106),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_141),
.B1(n_125),
.B2(n_118),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_110),
.B1(n_96),
.B2(n_74),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_124),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_108),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_153),
.C(n_155),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_150),
.B1(n_117),
.B2(n_133),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_112),
.B(n_103),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_68),
.B1(n_80),
.B2(n_46),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_154),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_58),
.C(n_13),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_46),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_115),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_158),
.A2(n_117),
.B1(n_46),
.B2(n_26),
.Y(n_193)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_166),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_177),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_173),
.C(n_174),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_136),
.B1(n_154),
.B2(n_140),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_176),
.B1(n_140),
.B2(n_150),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_122),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_144),
.C(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_147),
.B(n_122),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_120),
.C(n_133),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_179),
.A2(n_166),
.B1(n_163),
.B2(n_159),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_136),
.B1(n_120),
.B2(n_153),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_190),
.B1(n_182),
.B2(n_181),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_186),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_155),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_156),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_191),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_189),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_120),
.B(n_140),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_185),
.B(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_24),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_174),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_58),
.C(n_24),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_186),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_201),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_191),
.B(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_190),
.A2(n_173),
.B1(n_169),
.B2(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_205),
.B1(n_207),
.B2(n_2),
.Y(n_218)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_169),
.B1(n_158),
.B2(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_210),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_178),
.B1(n_162),
.B2(n_80),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_208),
.B(n_12),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_13),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

AOI321xp33_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_183),
.A3(n_194),
.B1(n_12),
.B2(n_13),
.C(n_25),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_220),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_58),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_218),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_26),
.C(n_25),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_221),
.C(n_222),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_12),
.C(n_3),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_26),
.C(n_25),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_200),
.B(n_205),
.C(n_203),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_224),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_217),
.A2(n_198),
.B1(n_209),
.B2(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_225),
.B(n_228),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_210),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_227),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_26),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_4),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_2),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_3),
.C(n_4),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_220),
.B1(n_212),
.B2(n_5),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_4),
.B(n_5),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_3),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_4),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_246),
.B1(n_237),
.B2(n_238),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_223),
.B(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_243),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_234),
.A2(n_224),
.B(n_5),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_5),
.C(n_6),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_249),
.B(n_250),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_244),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_248),
.A2(n_235),
.B(n_237),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_224),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_251),
.C(n_7),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_6),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_6),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_256),
.A2(n_11),
.B(n_9),
.Y(n_257)
);

OAI222xp33_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_241),
.C2(n_220),
.Y(n_258)
);


endmodule