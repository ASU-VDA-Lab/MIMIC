module real_aes_9083_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1170;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1175;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_905;
wire n_792;
wire n_503;
wire n_635;
wire n_518;
wire n_673;
wire n_1067;
wire n_878;
wire n_1192;
wire n_665;
wire n_991;
wire n_667;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_559;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_1137;
wire n_448;
wire n_556;
wire n_545;
wire n_752;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_666;
wire n_884;
wire n_537;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_1140;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_994;
wire n_495;
wire n_1072;
wire n_892;
wire n_1078;
wire n_938;
wire n_744;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_1049;
wire n_1182;
wire n_872;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_1189;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_746;
wire n_1168;
wire n_656;
wire n_1025;
wire n_1148;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_996;
wire n_523;
wire n_860;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_725;
wire n_504;
wire n_455;
wire n_973;
wire n_671;
wire n_1084;
wire n_960;
wire n_1081;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_940;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_1100;
wire n_1167;
wire n_1174;
wire n_1193;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_1006;
wire n_417;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_1142;
wire n_508;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_1145;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_1073;
wire n_735;
wire n_728;
wire n_713;
wire n_1179;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1157;
wire n_1158;
wire n_1132;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_1187;
wire n_1003;
wire n_533;
wire n_1014;
wire n_1028;
wire n_1000;
wire n_1083;
wire n_727;
wire n_1056;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_1127;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_1162;
wire n_861;
wire n_705;
wire n_1191;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_823;
wire n_1172;
wire n_863;
wire n_756;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1166;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1190;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_1045;
wire n_871;
wire n_1156;
wire n_1159;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_650;
wire n_646;
wire n_710;
wire n_743;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1185;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_1102;
wire n_447;
wire n_1101;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_802;
wire n_877;
wire n_868;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g679 ( .A(n_0), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_1), .A2(n_255), .B1(n_535), .B2(n_1006), .Y(n_1005) );
AOI222xp33_ASAP7_75t_L g941 ( .A1(n_2), .A2(n_193), .B1(n_350), .B2(n_483), .C1(n_490), .C2(n_554), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_3), .A2(n_103), .B1(n_521), .B2(n_522), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_4), .A2(n_343), .B1(n_467), .B2(n_521), .C(n_914), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_5), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_6), .A2(n_172), .B1(n_620), .B2(n_895), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_7), .A2(n_94), .B1(n_804), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_8), .A2(n_248), .B1(n_621), .B2(n_701), .Y(n_963) );
NAND2xp5_ASAP7_75t_SL g889 ( .A(n_9), .B(n_890), .Y(n_889) );
AO22x2_ASAP7_75t_L g420 ( .A1(n_10), .A2(n_234), .B1(n_421), .B2(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g1138 ( .A(n_10), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_11), .A2(n_183), .B1(n_464), .B2(n_867), .Y(n_934) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_12), .A2(n_374), .B1(n_660), .B2(n_725), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_13), .Y(n_974) );
AOI222xp33_ASAP7_75t_L g1186 ( .A1(n_14), .A2(n_64), .B1(n_344), .B2(n_553), .C1(n_564), .C2(n_878), .Y(n_1186) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_15), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_16), .Y(n_628) );
INVx1_ASAP7_75t_L g771 ( .A(n_17), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_18), .A2(n_207), .B1(n_540), .B2(n_576), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_19), .A2(n_266), .B1(n_459), .B2(n_468), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_20), .A2(n_106), .B1(n_521), .B2(n_531), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_21), .A2(n_335), .B1(n_530), .B2(n_531), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_22), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_23), .A2(n_336), .B1(n_441), .B2(n_448), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_24), .A2(n_328), .B1(n_467), .B2(n_579), .Y(n_578) );
AOI222xp33_ASAP7_75t_L g877 ( .A1(n_25), .A2(n_72), .B1(n_300), .B2(n_614), .C1(n_660), .C2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_26), .A2(n_246), .B1(n_448), .B2(n_849), .Y(n_1054) );
AOI22xp5_ASAP7_75t_SL g713 ( .A1(n_27), .A2(n_264), .B1(n_714), .B2(n_715), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_28), .A2(n_39), .B1(n_539), .B2(n_576), .C(n_919), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g1181 ( .A1(n_29), .A2(n_260), .B1(n_576), .B2(n_1182), .C(n_1183), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_30), .A2(n_269), .B1(n_464), .B2(n_630), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_31), .A2(n_1168), .B1(n_1187), .B2(n_1188), .Y(n_1167) );
INVx1_ASAP7_75t_L g1187 ( .A(n_31), .Y(n_1187) );
CKINVDCx20_ASAP7_75t_R g975 ( .A(n_32), .Y(n_975) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_33), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_34), .A2(n_261), .B1(n_804), .B2(n_867), .Y(n_1021) );
AO22x2_ASAP7_75t_L g424 ( .A1(n_35), .A2(n_124), .B1(n_421), .B2(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g1036 ( .A(n_36), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_37), .A2(n_187), .B1(n_449), .B2(n_460), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_38), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_40), .Y(n_842) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_41), .A2(n_65), .B1(n_464), .B2(n_850), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g1185 ( .A(n_42), .Y(n_1185) );
INVx1_ASAP7_75t_L g653 ( .A(n_43), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_44), .A2(n_311), .B1(n_554), .B2(n_1015), .Y(n_1014) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_45), .A2(n_66), .B1(n_466), .B2(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g747 ( .A(n_46), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_47), .A2(n_177), .B1(n_867), .B2(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g916 ( .A(n_48), .Y(n_916) );
INVx1_ASAP7_75t_L g1112 ( .A(n_49), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_50), .A2(n_224), .B1(n_497), .B2(n_549), .Y(n_651) );
AOI222xp33_ASAP7_75t_L g922 ( .A1(n_51), .A2(n_144), .B1(n_155), .B2(n_490), .C1(n_495), .C2(n_923), .Y(n_922) );
AOI222xp33_ASAP7_75t_L g550 ( .A1(n_52), .A2(n_316), .B1(n_334), .B2(n_551), .C1(n_552), .C2(n_553), .Y(n_550) );
AOI22xp5_ASAP7_75t_SL g711 ( .A1(n_53), .A2(n_332), .B1(n_625), .B2(n_712), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g942 ( .A(n_54), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_55), .A2(n_125), .B1(n_846), .B2(n_954), .Y(n_953) );
AOI22xp5_ASAP7_75t_SL g799 ( .A1(n_56), .A2(n_233), .B1(n_468), .B2(n_712), .Y(n_799) );
INVx1_ASAP7_75t_L g779 ( .A(n_57), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_58), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_59), .A2(n_190), .B1(n_448), .B2(n_1156), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_60), .A2(n_345), .B1(n_572), .B2(n_872), .Y(n_871) );
CKINVDCx16_ASAP7_75t_R g595 ( .A(n_61), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_62), .A2(n_319), .B1(n_606), .B2(n_969), .Y(n_1147) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_63), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g1179 ( .A(n_67), .Y(n_1179) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_68), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g700 ( .A1(n_69), .A2(n_263), .B1(n_621), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_70), .A2(n_380), .B1(n_433), .B2(n_583), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_71), .A2(n_290), .B1(n_568), .B2(n_608), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_73), .A2(n_93), .B1(n_554), .B2(n_572), .Y(n_1113) );
INVx1_ASAP7_75t_L g1041 ( .A(n_74), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_75), .A2(n_135), .B1(n_792), .B2(n_875), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_76), .A2(n_368), .B1(n_464), .B2(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g677 ( .A(n_77), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_78), .B(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_79), .A2(n_216), .B1(n_701), .B2(n_1003), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_80), .A2(n_230), .B1(n_540), .B2(n_544), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_81), .A2(n_244), .B1(n_846), .B2(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g993 ( .A(n_82), .Y(n_993) );
INVx1_ASAP7_75t_L g776 ( .A(n_83), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_84), .A2(n_242), .B1(n_593), .B2(n_705), .Y(n_704) );
AOI22xp5_ASAP7_75t_SL g803 ( .A1(n_85), .A2(n_97), .B1(n_593), .B2(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g757 ( .A(n_86), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_87), .A2(n_160), .B1(n_853), .B2(n_1159), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_88), .A2(n_167), .B1(n_621), .B2(n_741), .Y(n_740) );
AO22x2_ASAP7_75t_L g430 ( .A1(n_89), .A2(n_278), .B1(n_421), .B2(n_422), .Y(n_430) );
INVx1_ASAP7_75t_L g1135 ( .A(n_89), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_90), .A2(n_289), .B1(n_442), .B2(n_449), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_91), .A2(n_92), .B1(n_707), .B2(n_961), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_95), .A2(n_308), .B1(n_448), .B2(n_849), .Y(n_848) );
OA22x2_ASAP7_75t_L g516 ( .A1(n_96), .A2(n_517), .B1(n_518), .B2(n_555), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_96), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_98), .A2(n_219), .B1(n_535), .B2(n_666), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_99), .A2(n_118), .B1(n_804), .B2(n_875), .Y(n_1118) );
INVx1_ASAP7_75t_L g745 ( .A(n_100), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_101), .A2(n_109), .B1(n_552), .B2(n_725), .Y(n_1017) );
INVx1_ASAP7_75t_L g796 ( .A(n_102), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_104), .A2(n_250), .B1(n_741), .B2(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g733 ( .A(n_105), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_107), .A2(n_169), .B1(n_546), .B2(n_606), .Y(n_692) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_108), .A2(n_226), .B1(n_539), .B2(n_574), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_110), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_111), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_112), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_113), .B(n_1108), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_114), .A2(n_150), .B1(n_530), .B2(n_910), .Y(n_1053) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_115), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_116), .A2(n_258), .B1(n_442), .B2(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g1146 ( .A(n_117), .Y(n_1146) );
AOI22xp5_ASAP7_75t_L g1098 ( .A1(n_119), .A2(n_299), .B1(n_705), .B2(n_712), .Y(n_1098) );
INVx1_ASAP7_75t_L g738 ( .A(n_120), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g1073 ( .A(n_121), .Y(n_1073) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_122), .Y(n_589) );
INVx1_ASAP7_75t_L g1094 ( .A(n_123), .Y(n_1094) );
INVx1_ASAP7_75t_L g1139 ( .A(n_124), .Y(n_1139) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_126), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g1184 ( .A(n_127), .Y(n_1184) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_128), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_129), .Y(n_959) );
AOI22xp5_ASAP7_75t_L g1092 ( .A1(n_130), .A2(n_214), .B1(n_547), .B2(n_565), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_131), .A2(n_139), .B1(n_535), .B2(n_1079), .Y(n_1121) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_132), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_133), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_133), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_134), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_136), .A2(n_217), .B1(n_846), .B2(n_847), .Y(n_1154) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_137), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_138), .A2(n_279), .B1(n_606), .B2(n_969), .Y(n_968) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_140), .Y(n_472) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_141), .A2(n_551), .B(n_598), .C(n_609), .Y(n_597) );
INVx1_ASAP7_75t_L g1102 ( .A(n_142), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_143), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g1145 ( .A(n_145), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g952 ( .A(n_146), .Y(n_952) );
INVx1_ASAP7_75t_L g1122 ( .A(n_147), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_148), .A2(n_186), .B1(n_784), .B2(n_875), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_149), .A2(n_354), .B1(n_533), .B2(n_536), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_151), .A2(n_276), .B1(n_568), .B2(n_608), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_152), .A2(n_256), .B1(n_954), .B2(n_1049), .Y(n_1048) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_153), .A2(n_232), .B1(n_458), .B2(n_581), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_154), .Y(n_591) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_156), .A2(n_583), .B(n_584), .C(n_590), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_157), .A2(n_378), .B1(n_660), .B2(n_725), .Y(n_1110) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_158), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_159), .A2(n_730), .B1(n_761), .B2(n_762), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g761 ( .A(n_159), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_161), .A2(n_285), .B1(n_531), .B2(n_853), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_162), .A2(n_199), .B1(n_449), .B2(n_850), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_163), .A2(n_376), .B1(n_546), .B2(n_606), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g1169 ( .A1(n_164), .A2(n_227), .B1(n_522), .B2(n_1082), .C(n_1170), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_165), .A2(n_293), .B1(n_546), .B2(n_549), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_166), .Y(n_456) );
AND2x6_ASAP7_75t_L g401 ( .A(n_168), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_168), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_170), .A2(n_324), .B1(n_535), .B2(n_699), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_171), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_173), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_174), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_175), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_176), .A2(n_277), .B1(n_495), .B2(n_564), .Y(n_1070) );
AOI22xp33_ASAP7_75t_SL g1120 ( .A1(n_178), .A2(n_372), .B1(n_579), .B2(n_850), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_179), .A2(n_254), .B1(n_549), .B2(n_554), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_180), .A2(n_388), .B1(n_804), .B2(n_867), .Y(n_897) );
AO22x1_ASAP7_75t_L g909 ( .A1(n_181), .A2(n_196), .B1(n_910), .B2(n_912), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_182), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g908 ( .A1(n_184), .A2(n_353), .B1(n_625), .B2(n_630), .C(n_909), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_185), .A2(n_287), .B1(n_525), .B2(n_527), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g1095 ( .A1(n_188), .A2(n_394), .B1(n_496), .B2(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1065 ( .A(n_189), .Y(n_1065) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_191), .A2(n_399), .B(n_407), .C(n_1140), .Y(n_398) );
INVx1_ASAP7_75t_L g997 ( .A(n_192), .Y(n_997) );
INVx1_ASAP7_75t_L g753 ( .A(n_194), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_195), .Y(n_462) );
AOI22xp33_ASAP7_75t_SL g1099 ( .A1(n_197), .A2(n_200), .B1(n_911), .B2(n_1079), .Y(n_1099) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_198), .A2(n_265), .B1(n_421), .B2(n_425), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g1136 ( .A(n_198), .B(n_1137), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g1176 ( .A1(n_201), .A2(n_218), .B1(n_521), .B2(n_1177), .C(n_1178), .Y(n_1176) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_202), .A2(n_286), .B1(n_625), .B2(n_715), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_203), .A2(n_327), .B1(n_568), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_204), .A2(n_267), .B1(n_784), .B2(n_801), .Y(n_931) );
AOI22xp33_ASAP7_75t_SL g1100 ( .A1(n_205), .A2(n_365), .B1(n_468), .B2(n_784), .Y(n_1100) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_206), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_208), .A2(n_397), .B1(n_568), .B2(n_660), .Y(n_994) );
INVx1_ASAP7_75t_L g990 ( .A(n_209), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_210), .A2(n_352), .B1(n_707), .B2(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g996 ( .A(n_211), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_212), .Y(n_569) );
AOI22xp5_ASAP7_75t_SL g717 ( .A1(n_213), .A2(n_295), .B1(n_666), .B2(n_699), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_215), .A2(n_251), .B1(n_581), .B2(n_867), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_220), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_221), .B(n_939), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_222), .A2(n_370), .B1(n_546), .B2(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_223), .A2(n_412), .B1(n_512), .B2(n_513), .Y(n_411) );
INVx1_ASAP7_75t_L g512 ( .A(n_223), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_225), .Y(n_966) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_228), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_229), .A2(n_905), .B1(n_906), .B2(n_924), .Y(n_904) );
INVx1_ASAP7_75t_L g924 ( .A(n_229), .Y(n_924) );
INVx1_ASAP7_75t_L g1039 ( .A(n_231), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g967 ( .A(n_235), .Y(n_967) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_236), .A2(n_828), .B1(n_858), .B2(n_859), .Y(n_827) );
INVx1_ASAP7_75t_L g858 ( .A(n_236), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_237), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_238), .A2(n_253), .B1(n_464), .B2(n_467), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_239), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g1180 ( .A(n_240), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_241), .A2(n_373), .B1(n_533), .B2(n_536), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_243), .B(n_576), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_245), .A2(n_384), .B1(n_581), .B2(n_911), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_247), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_249), .A2(n_291), .B1(n_698), .B2(n_699), .Y(n_697) );
AOI22xp5_ASAP7_75t_SL g1031 ( .A1(n_252), .A2(n_1032), .B1(n_1055), .B2(n_1056), .Y(n_1031) );
INVx1_ASAP7_75t_L g1056 ( .A(n_252), .Y(n_1056) );
INVx2_ASAP7_75t_L g406 ( .A(n_257), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_259), .A2(n_342), .B1(n_497), .B2(n_660), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_262), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_268), .A2(n_284), .B1(n_625), .B2(n_705), .Y(n_868) );
INVx1_ASAP7_75t_L g1035 ( .A(n_270), .Y(n_1035) );
OA22x2_ASAP7_75t_L g765 ( .A1(n_271), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_271), .Y(n_766) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_272), .A2(n_307), .B1(n_792), .B2(n_793), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_273), .A2(n_945), .B1(n_976), .B2(n_977), .Y(n_944) );
INVx1_ASAP7_75t_L g976 ( .A(n_273), .Y(n_976) );
INVx1_ASAP7_75t_L g1045 ( .A(n_274), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_275), .A2(n_331), .B1(n_459), .B2(n_875), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_280), .A2(n_330), .B1(n_620), .B2(n_621), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_281), .A2(n_379), .B1(n_707), .B2(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g650 ( .A(n_282), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_283), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_288), .A2(n_367), .B1(n_698), .B2(n_1077), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_292), .A2(n_333), .B1(n_539), .B2(n_543), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g888 ( .A(n_294), .B(n_576), .Y(n_888) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_296), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_297), .A2(n_348), .B1(n_954), .B2(n_1162), .Y(n_1161) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_298), .A2(n_382), .B1(n_576), .B2(n_604), .Y(n_870) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_301), .A2(n_396), .B1(n_630), .B2(n_707), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_302), .Y(n_810) );
INVx1_ASAP7_75t_L g421 ( .A(n_303), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_303), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_304), .A2(n_310), .B1(n_539), .B2(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g991 ( .A(n_305), .Y(n_991) );
INVx1_ASAP7_75t_L g750 ( .A(n_306), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_309), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_312), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_313), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_314), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g1101 ( .A1(n_315), .A2(n_357), .B1(n_536), .B2(n_875), .Y(n_1101) );
INVx1_ASAP7_75t_L g739 ( .A(n_317), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_318), .Y(n_818) );
INVx1_ASAP7_75t_L g1066 ( .A(n_320), .Y(n_1066) );
CKINVDCx20_ASAP7_75t_R g1174 ( .A(n_321), .Y(n_1174) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_322), .A2(n_366), .B1(n_547), .B2(n_572), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_323), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_325), .B(n_495), .Y(n_1042) );
CKINVDCx20_ASAP7_75t_R g1149 ( .A(n_326), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_329), .A2(n_358), .B1(n_608), .B2(n_725), .Y(n_940) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_337), .Y(n_684) );
AND2x2_ASAP7_75t_L g405 ( .A(n_338), .B(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_SL g1061 ( .A1(n_339), .A2(n_1062), .B1(n_1083), .B2(n_1084), .Y(n_1061) );
INVx1_ASAP7_75t_L g1084 ( .A(n_339), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_340), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g402 ( .A(n_341), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_346), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_347), .B(n_939), .Y(n_1109) );
INVx1_ASAP7_75t_L g760 ( .A(n_349), .Y(n_760) );
INVx1_ASAP7_75t_L g681 ( .A(n_351), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_355), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_356), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g780 ( .A(n_359), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_360), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_361), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_362), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_363), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_364), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g1171 ( .A(n_369), .Y(n_1171) );
INVx1_ASAP7_75t_L g631 ( .A(n_371), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_375), .B(n_939), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_377), .A2(n_1142), .B1(n_1163), .B2(n_1164), .Y(n_1141) );
CKINVDCx20_ASAP7_75t_R g1163 ( .A(n_377), .Y(n_1163) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_381), .Y(n_626) );
INVx1_ASAP7_75t_L g773 ( .A(n_383), .Y(n_773) );
INVx1_ASAP7_75t_L g1044 ( .A(n_385), .Y(n_1044) );
INVx1_ASAP7_75t_L g915 ( .A(n_386), .Y(n_915) );
XNOR2xp5_ASAP7_75t_L g557 ( .A(n_387), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g735 ( .A(n_389), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g1151 ( .A(n_390), .Y(n_1151) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_391), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_392), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_393), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_395), .Y(n_1013) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1131 ( .A(n_402), .Y(n_1131) );
OAI21xp5_ASAP7_75t_L g1193 ( .A1(n_403), .A2(n_1130), .B(n_1194), .Y(n_1193) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_821), .B1(n_1125), .B2(n_1126), .C(n_1127), .Y(n_407) );
INVx1_ASAP7_75t_L g1126 ( .A(n_408), .Y(n_1126) );
XOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_641), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_514), .B1(n_639), .B2(n_640), .Y(n_409) );
INVx3_ASAP7_75t_L g639 ( .A(n_410), .Y(n_639) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g513 ( .A(n_412), .Y(n_513) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_413), .B(n_470), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_452), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_431), .B1(n_432), .B2(n_439), .C(n_440), .Y(n_414) );
INVx2_ASAP7_75t_SL g531 ( .A(n_415), .Y(n_531) );
INVx4_ASAP7_75t_L g593 ( .A(n_415), .Y(n_593) );
INVx3_ASAP7_75t_L g625 ( .A(n_415), .Y(n_625) );
INVx11_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx11_ASAP7_75t_L g680 ( .A(n_416), .Y(n_680) );
AND2x6_ASAP7_75t_L g416 ( .A(n_417), .B(n_426), .Y(n_416) );
AND2x4_ASAP7_75t_L g542 ( .A(n_417), .B(n_461), .Y(n_542) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g475 ( .A(n_418), .B(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_424), .Y(n_418) );
AND2x2_ASAP7_75t_L g437 ( .A(n_419), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g447 ( .A(n_419), .B(n_424), .Y(n_447) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g487 ( .A(n_420), .B(n_428), .Y(n_487) );
AND2x2_ASAP7_75t_L g492 ( .A(n_420), .B(n_424), .Y(n_492) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_423), .Y(n_425) );
INVx2_ASAP7_75t_L g438 ( .A(n_424), .Y(n_438) );
INVx1_ASAP7_75t_L g451 ( .A(n_424), .Y(n_451) );
AND2x2_ASAP7_75t_L g455 ( .A(n_426), .B(n_437), .Y(n_455) );
AND2x4_ASAP7_75t_L g466 ( .A(n_426), .B(n_447), .Y(n_466) );
AND2x6_ASAP7_75t_L g491 ( .A(n_426), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
AND2x2_ASAP7_75t_L g461 ( .A(n_427), .B(n_430), .Y(n_461) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_428), .B(n_430), .Y(n_436) );
AND2x2_ASAP7_75t_L g445 ( .A(n_428), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g446 ( .A(n_430), .Y(n_446) );
INVx1_ASAP7_75t_L g486 ( .A(n_430), .Y(n_486) );
INVx2_ASAP7_75t_L g1049 ( .A(n_432), .Y(n_1049) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g912 ( .A(n_433), .Y(n_912) );
BUFx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g536 ( .A(n_434), .Y(n_536) );
BUFx3_ASAP7_75t_L g581 ( .A(n_434), .Y(n_581) );
INVx1_ASAP7_75t_L g674 ( .A(n_434), .Y(n_674) );
BUFx3_ASAP7_75t_L g699 ( .A(n_434), .Y(n_699) );
BUFx3_ASAP7_75t_L g804 ( .A(n_434), .Y(n_804) );
BUFx2_ASAP7_75t_SL g961 ( .A(n_434), .Y(n_961) );
BUFx2_ASAP7_75t_SL g1077 ( .A(n_434), .Y(n_1077) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
AND2x2_ASAP7_75t_L g666 ( .A(n_435), .B(n_504), .Y(n_666) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x6_ASAP7_75t_L g450 ( .A(n_436), .B(n_451), .Y(n_450) );
AND2x4_ASAP7_75t_L g460 ( .A(n_437), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g469 ( .A(n_437), .B(n_445), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_437), .B(n_445), .Y(n_634) );
AND2x2_ASAP7_75t_L g485 ( .A(n_438), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g504 ( .A(n_438), .Y(n_504) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx4_ASAP7_75t_L g526 ( .A(n_443), .Y(n_526) );
INVx1_ASAP7_75t_L g620 ( .A(n_443), .Y(n_620) );
INVx3_ASAP7_75t_L g712 ( .A(n_443), .Y(n_712) );
BUFx3_ASAP7_75t_L g742 ( .A(n_443), .Y(n_742) );
INVx5_ASAP7_75t_L g850 ( .A(n_443), .Y(n_850) );
INVx8_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_445), .B(n_447), .Y(n_586) );
INVx1_ASAP7_75t_L g511 ( .A(n_446), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_447), .B(n_461), .Y(n_480) );
AND2x6_ASAP7_75t_L g544 ( .A(n_447), .B(n_461), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g917 ( .A(n_448), .Y(n_917) );
BUFx4f_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g527 ( .A(n_449), .Y(n_527) );
BUFx2_ASAP7_75t_L g895 ( .A(n_449), .Y(n_895) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_449), .Y(n_1003) );
INVx6_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g621 ( .A(n_450), .Y(n_621) );
INVx1_ASAP7_75t_L g793 ( .A(n_450), .Y(n_793) );
INVx1_ASAP7_75t_SL g1079 ( .A(n_450), .Y(n_1079) );
INVx1_ASAP7_75t_L g548 ( .A(n_451), .Y(n_548) );
OAI221xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_456), .B1(n_457), .B2(n_462), .C(n_463), .Y(n_452) );
INVx2_ASAP7_75t_L g1082 ( .A(n_453), .Y(n_1082) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx3_ASAP7_75t_L g530 ( .A(n_454), .Y(n_530) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_454), .Y(n_630) );
BUFx3_ASAP7_75t_L g846 ( .A(n_454), .Y(n_846) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_SL g583 ( .A(n_455), .Y(n_583) );
INVx2_ASAP7_75t_L g668 ( .A(n_455), .Y(n_668) );
BUFx2_ASAP7_75t_SL g714 ( .A(n_455), .Y(n_714) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_460), .Y(n_535) );
INVx2_ASAP7_75t_L g663 ( .A(n_460), .Y(n_663) );
BUFx3_ASAP7_75t_L g792 ( .A(n_460), .Y(n_792) );
BUFx3_ASAP7_75t_L g911 ( .A(n_460), .Y(n_911) );
INVx1_ASAP7_75t_L g476 ( .A(n_461), .Y(n_476) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g521 ( .A(n_465), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_465), .A2(n_623), .B1(n_624), .B2(n_626), .Y(n_622) );
OAI22xp5_ASAP7_75t_SL g667 ( .A1(n_465), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_667) );
INVx2_ASAP7_75t_L g705 ( .A(n_465), .Y(n_705) );
OAI221xp5_ASAP7_75t_SL g737 ( .A1(n_465), .A2(n_632), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_737) );
INVx2_ASAP7_75t_L g853 ( .A(n_465), .Y(n_853) );
INVx6_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g579 ( .A(n_466), .Y(n_579) );
BUFx3_ASAP7_75t_L g715 ( .A(n_466), .Y(n_715) );
BUFx3_ASAP7_75t_L g790 ( .A(n_466), .Y(n_790) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g523 ( .A(n_468), .Y(n_523) );
BUFx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g708 ( .A(n_469), .Y(n_708) );
BUFx3_ASAP7_75t_L g857 ( .A(n_469), .Y(n_857) );
BUFx3_ASAP7_75t_L g867 ( .A(n_469), .Y(n_867) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_481), .C(n_500), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_477), .B2(n_478), .Y(n_471) );
OAI221xp5_ASAP7_75t_SL g965 ( .A1(n_473), .A2(n_774), .B1(n_966), .B2(n_967), .C(n_968), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_473), .A2(n_774), .B1(n_990), .B2(n_991), .Y(n_989) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_473), .A2(n_602), .B1(n_1065), .B2(n_1066), .Y(n_1064) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g746 ( .A(n_474), .Y(n_746) );
INVx2_ASAP7_75t_L g832 ( .A(n_474), .Y(n_832) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_475), .A2(n_650), .B(n_651), .Y(n_649) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_475), .Y(n_772) );
OAI22xp5_ASAP7_75t_SL g807 ( .A1(n_478), .A2(n_808), .B1(n_809), .B2(n_810), .Y(n_807) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_SL g1037 ( .A(n_479), .Y(n_1037) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g602 ( .A(n_480), .Y(n_602) );
OAI222xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_488), .B1(n_489), .B2(n_493), .C1(n_494), .C2(n_499), .Y(n_481) );
OAI222xp33_ASAP7_75t_L g1148 ( .A1(n_482), .A2(n_494), .B1(n_884), .B2(n_1149), .C1(n_1150), .C2(n_1151), .Y(n_1148) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx4f_ASAP7_75t_SL g552 ( .A(n_484), .Y(n_552) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_484), .Y(n_565) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_484), .Y(n_660) );
BUFx2_ASAP7_75t_L g752 ( .A(n_484), .Y(n_752) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g498 ( .A(n_486), .Y(n_498) );
AND2x4_ASAP7_75t_L g497 ( .A(n_487), .B(n_498), .Y(n_497) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_487), .B(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g547 ( .A(n_487), .B(n_548), .Y(n_547) );
OAI21xp5_ASAP7_75t_SL g687 ( .A1(n_489), .A2(n_688), .B(n_689), .Y(n_687) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g749 ( .A(n_490), .Y(n_749) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx3_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
INVx2_ASAP7_75t_L g561 ( .A(n_491), .Y(n_561) );
INVx2_ASAP7_75t_SL g657 ( .A(n_491), .Y(n_657) );
INVx4_ASAP7_75t_L g815 ( .A(n_491), .Y(n_815) );
INVx2_ASAP7_75t_L g884 ( .A(n_491), .Y(n_884) );
INVx1_ASAP7_75t_L g509 ( .A(n_492), .Y(n_509) );
AND2x4_ASAP7_75t_L g549 ( .A(n_492), .B(n_511), .Y(n_549) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g837 ( .A(n_496), .Y(n_837) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx12f_ASAP7_75t_L g554 ( .A(n_497), .Y(n_554) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_497), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_505), .B2(n_506), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g1071 ( .A1(n_502), .A2(n_1072), .B1(n_1073), .B2(n_1074), .Y(n_1071) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_503), .A2(n_602), .B1(n_653), .B2(n_654), .Y(n_652) );
INVx4_ASAP7_75t_L g759 ( .A(n_503), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_503), .A2(n_611), .B1(n_779), .B2(n_780), .Y(n_778) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_503), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_503), .A2(n_506), .B1(n_920), .B2(n_921), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_503), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_506), .A2(n_757), .B1(n_758), .B2(n_760), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_506), .A2(n_840), .B1(n_841), .B2(n_842), .Y(n_839) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g1074 ( .A(n_507), .Y(n_1074) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g998 ( .A(n_508), .Y(n_998) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g640 ( .A(n_514), .Y(n_640) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_556), .B1(n_637), .B2(n_638), .Y(n_515) );
INVx1_ASAP7_75t_L g638 ( .A(n_516), .Y(n_638) );
INVx1_ASAP7_75t_SL g555 ( .A(n_518), .Y(n_555) );
NAND4xp75_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .C(n_537), .D(n_550), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g702 ( .A(n_526), .Y(n_702) );
INVx1_ASAP7_75t_L g588 ( .A(n_527), .Y(n_588) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .Y(n_528) );
INVx1_ASAP7_75t_L g734 ( .A(n_531), .Y(n_734) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g1177 ( .A(n_534), .Y(n_1177) );
INVx4_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_SL g537 ( .A(n_538), .B(n_545), .Y(n_537) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx5_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g604 ( .A(n_541), .Y(n_604) );
INVx2_ASAP7_75t_L g890 ( .A(n_541), .Y(n_890) );
INVx2_ASAP7_75t_L g939 ( .A(n_541), .Y(n_939) );
INVx4_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx4f_ASAP7_75t_L g576 ( .A(n_544), .Y(n_576) );
INVx1_ASAP7_75t_SL g695 ( .A(n_544), .Y(n_695) );
BUFx2_ASAP7_75t_L g1108 ( .A(n_544), .Y(n_1108) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g725 ( .A(n_547), .Y(n_725) );
BUFx2_ASAP7_75t_L g872 ( .A(n_547), .Y(n_872) );
INVx1_ASAP7_75t_L g970 ( .A(n_547), .Y(n_970) );
BUFx3_ASAP7_75t_L g572 ( .A(n_549), .Y(n_572) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_549), .Y(n_608) );
BUFx2_ASAP7_75t_SL g1015 ( .A(n_549), .Y(n_1015) );
BUFx2_ASAP7_75t_SL g1096 ( .A(n_549), .Y(n_1096) );
INVx3_ASAP7_75t_L g1069 ( .A(n_551), .Y(n_1069) );
INVx1_ASAP7_75t_L g972 ( .A(n_552), .Y(n_972) );
BUFx4f_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g615 ( .A(n_554), .Y(n_615) );
INVx1_ASAP7_75t_L g637 ( .A(n_556), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_594), .B1(n_635), .B2(n_636), .Y(n_556) );
INVx1_ASAP7_75t_L g636 ( .A(n_557), .Y(n_636) );
NAND3x1_ASAP7_75t_L g558 ( .A(n_559), .B(n_577), .C(n_582), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_570), .Y(n_559) );
OAI222xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B1(n_563), .B2(n_566), .C1(n_567), .C2(n_569), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g720 ( .A1(n_561), .A2(n_721), .B(n_722), .Y(n_720) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g611 ( .A(n_565), .Y(n_611) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx4f_ASAP7_75t_L g755 ( .A(n_568), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
OAI22xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_585), .A2(n_915), .B1(n_916), .B2(n_917), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_585), .A2(n_588), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
BUFx2_ASAP7_75t_R g585 ( .A(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_586), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g635 ( .A(n_594), .Y(n_635) );
XNOR2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_616), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_603), .C(n_605), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_600), .A2(n_832), .B1(n_1145), .B2(n_1146), .C(n_1147), .Y(n_1144) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_602), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_744) );
BUFx3_ASAP7_75t_L g774 ( .A(n_602), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_602), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_830) );
OA211x2_ASAP7_75t_L g936 ( .A1(n_602), .A2(n_937), .B(n_938), .C(n_940), .Y(n_936) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_612), .B2(n_613), .Y(n_609) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_622), .C(n_627), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_631), .B2(n_632), .Y(n_627) );
OAI221xp5_ASAP7_75t_SL g732 ( .A1(n_629), .A2(n_733), .B1(n_734), .B2(n_735), .C(n_736), .Y(n_732) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_634), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B1(n_728), .B2(n_820), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
XNOR2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_682), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
XOR2x2_ASAP7_75t_L g794 ( .A(n_646), .B(n_795), .Y(n_794) );
XNOR2x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_681), .Y(n_646) );
AND3x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_661), .C(n_671), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .C(n_655), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_655) );
OAI222xp33_ASAP7_75t_L g971 ( .A1(n_657), .A2(n_837), .B1(n_972), .B2(n_973), .C1(n_974), .C2(n_975), .Y(n_971) );
OAI222xp33_ASAP7_75t_L g834 ( .A1(n_659), .A2(n_749), .B1(n_835), .B2(n_836), .C1(n_837), .C2(n_838), .Y(n_834) );
INVx3_ASAP7_75t_L g923 ( .A(n_659), .Y(n_923) );
INVx4_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g690 ( .A(n_660), .Y(n_690) );
INVx2_ASAP7_75t_L g817 ( .A(n_660), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_667), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_664), .B(n_665), .Y(n_662) );
INVx2_ASAP7_75t_L g698 ( .A(n_663), .Y(n_698) );
INVx1_ASAP7_75t_L g847 ( .A(n_663), .Y(n_847) );
INVx3_ASAP7_75t_L g801 ( .A(n_668), .Y(n_801) );
INVx3_ASAP7_75t_L g875 ( .A(n_668), .Y(n_875) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_676), .C(n_678), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx5_ASAP7_75t_SL g784 ( .A(n_680), .Y(n_784) );
INVx1_ASAP7_75t_L g949 ( .A(n_680), .Y(n_949) );
INVx2_ASAP7_75t_L g1051 ( .A(n_680), .Y(n_1051) );
INVx2_ASAP7_75t_SL g1117 ( .A(n_680), .Y(n_1117) );
INVx4_ASAP7_75t_L g1173 ( .A(n_680), .Y(n_1173) );
XOR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_709), .Y(n_682) );
XNOR2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_696), .C(n_703), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_691), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .Y(n_696) );
INVx1_ASAP7_75t_L g1175 ( .A(n_699), .Y(n_1175) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
BUFx4f_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g955 ( .A(n_708), .Y(n_955) );
XOR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_727), .Y(n_709) );
NAND4xp75_ASAP7_75t_SL g710 ( .A(n_711), .B(n_713), .C(n_716), .D(n_719), .Y(n_710) );
INVx1_ASAP7_75t_L g951 ( .A(n_715), .Y(n_951) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_723), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx2_ASAP7_75t_L g820 ( .A(n_728), .Y(n_820) );
XNOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_763), .Y(n_728) );
INVx1_ASAP7_75t_L g762 ( .A(n_730), .Y(n_762) );
AND2x2_ASAP7_75t_SL g730 ( .A(n_731), .B(n_743), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_737), .Y(n_731) );
INVx3_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .C(n_756), .Y(n_743) );
OAI221xp5_ASAP7_75t_SL g748 ( .A1(n_749), .A2(n_750), .B1(n_751), .B2(n_753), .C(n_754), .Y(n_748) );
OAI21xp33_ASAP7_75t_L g775 ( .A1(n_749), .A2(n_776), .B(n_777), .Y(n_775) );
OAI21xp33_ASAP7_75t_SL g992 ( .A1(n_749), .A2(n_993), .B(n_994), .Y(n_992) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_749), .A2(n_1039), .B1(n_1040), .B2(n_1041), .C(n_1042), .Y(n_1038) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_758), .A2(n_998), .B1(n_1184), .B2(n_1185), .Y(n_1183) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx3_ASAP7_75t_SL g809 ( .A(n_759), .Y(n_809) );
AO22x2_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_794), .B2(n_819), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_781), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_775), .C(n_778), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_770) );
OAI21xp5_ASAP7_75t_SL g811 ( .A1(n_772), .A2(n_812), .B(n_813), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_772), .A2(n_1035), .B1(n_1036), .B2(n_1037), .Y(n_1034) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_786), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_785), .Y(n_782) );
INVx1_ASAP7_75t_L g1007 ( .A(n_784), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_791), .Y(n_786) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx3_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
BUFx2_ASAP7_75t_L g958 ( .A(n_792), .Y(n_958) );
INVx2_ASAP7_75t_L g819 ( .A(n_794), .Y(n_819) );
XNOR2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
NAND3x1_ASAP7_75t_SL g797 ( .A(n_798), .B(n_802), .C(n_806), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
BUFx2_ASAP7_75t_L g1162 ( .A(n_804), .Y(n_1162) );
NOR3xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_811), .C(n_814), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_809), .A2(n_998), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
OAI22xp5_ASAP7_75t_SL g814 ( .A1(n_815), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_814) );
INVx4_ASAP7_75t_L g878 ( .A(n_815), .Y(n_878) );
INVx1_ASAP7_75t_L g1125 ( .A(n_821), .Y(n_1125) );
XNOR2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_979), .Y(n_821) );
XOR2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_901), .Y(n_822) );
INVx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
BUFx3_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_827), .B1(n_860), .B2(n_861), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g859 ( .A(n_828), .Y(n_859) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_843), .Y(n_828) );
NOR3xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_834), .C(n_839), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_844), .B(n_851), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .Y(n_844) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
BUFx2_ASAP7_75t_L g1156 ( .A(n_850), .Y(n_1156) );
NAND2xp5_ASAP7_75t_SL g851 ( .A(n_852), .B(n_854), .Y(n_851) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AO22x2_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_880), .B2(n_900), .Y(n_861) );
AO22x1_ASAP7_75t_SL g927 ( .A1(n_862), .A2(n_863), .B1(n_928), .B2(n_943), .Y(n_927) );
INVx2_ASAP7_75t_SL g862 ( .A(n_863), .Y(n_862) );
XOR2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_879), .Y(n_863) );
NAND4xp75_ASAP7_75t_L g864 ( .A(n_865), .B(n_869), .C(n_873), .D(n_877), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_868), .Y(n_865) );
AND2x2_ASAP7_75t_SL g869 ( .A(n_870), .B(n_871), .Y(n_869) );
AND2x2_ASAP7_75t_L g873 ( .A(n_874), .B(n_876), .Y(n_873) );
INVx4_ASAP7_75t_SL g900 ( .A(n_880), .Y(n_900) );
OA22x2_ASAP7_75t_L g1030 ( .A1(n_880), .A2(n_900), .B1(n_1031), .B2(n_1057), .Y(n_1030) );
XOR2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_899), .Y(n_880) );
NAND3x1_ASAP7_75t_L g881 ( .A(n_882), .B(n_892), .C(n_896), .Y(n_881) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_887), .Y(n_882) );
OAI21xp5_ASAP7_75t_SL g883 ( .A1(n_884), .A2(n_885), .B(n_886), .Y(n_883) );
OAI21xp5_ASAP7_75t_L g1012 ( .A1(n_884), .A2(n_1013), .B(n_1014), .Y(n_1012) );
OAI21xp5_ASAP7_75t_L g1093 ( .A1(n_884), .A2(n_1094), .B(n_1095), .Y(n_1093) );
OAI21xp5_ASAP7_75t_SL g1111 ( .A1(n_884), .A2(n_1112), .B(n_1113), .Y(n_1111) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .C(n_891), .Y(n_887) );
BUFx2_ASAP7_75t_L g1182 ( .A(n_890), .Y(n_1182) );
AND2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
XNOR2xp5_ASAP7_75t_SL g901 ( .A(n_902), .B(n_925), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx2_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AND4x1_ASAP7_75t_L g907 ( .A(n_908), .B(n_913), .C(n_918), .D(n_922), .Y(n_907) );
BUFx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g1040 ( .A(n_923), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_927), .B1(n_944), .B2(n_978), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx2_ASAP7_75t_SL g943 ( .A(n_928), .Y(n_943) );
XOR2x2_ASAP7_75t_L g928 ( .A(n_929), .B(n_942), .Y(n_928) );
NAND4xp75_ASAP7_75t_L g929 ( .A(n_930), .B(n_933), .C(n_936), .D(n_941), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .Y(n_930) );
AND2x2_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
INVx1_ASAP7_75t_L g978 ( .A(n_944), .Y(n_978) );
INVx1_ASAP7_75t_L g977 ( .A(n_945), .Y(n_977) );
AND2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_964), .Y(n_945) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_947), .B(n_956), .Y(n_946) );
OAI221xp5_ASAP7_75t_SL g947 ( .A1(n_948), .A2(n_950), .B1(n_951), .B2(n_952), .C(n_953), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
OAI221xp5_ASAP7_75t_SL g956 ( .A1(n_957), .A2(n_959), .B1(n_960), .B2(n_962), .C(n_963), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
NOR2xp33_ASAP7_75t_SL g964 ( .A(n_965), .B(n_971), .Y(n_964) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
XOR2xp5_ASAP7_75t_L g979 ( .A(n_980), .B(n_1028), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
BUFx2_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
AO22x1_ASAP7_75t_L g982 ( .A1(n_983), .A2(n_984), .B1(n_1009), .B2(n_1027), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx1_ASAP7_75t_SL g986 ( .A(n_987), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_988), .B(n_999), .Y(n_987) );
NOR3xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_992), .C(n_995), .Y(n_988) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1004), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1002), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1008), .Y(n_1004) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx3_ASAP7_75t_SL g1027 ( .A(n_1009), .Y(n_1027) );
XOR2x2_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1026), .Y(n_1009) );
NAND2xp5_ASAP7_75t_SL g1010 ( .A(n_1011), .B(n_1019), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1016), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1018), .Y(n_1016) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1023), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1022), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g1028 ( .A1(n_1029), .A2(n_1030), .B1(n_1058), .B2(n_1059), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1031), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1055 ( .A(n_1032), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1046), .Y(n_1032) );
NOR3xp33_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1038), .C(n_1043), .Y(n_1033) );
NOR2xp33_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1052), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1050), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1054), .Y(n_1052) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
OA22x2_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1085), .B1(n_1123), .B2(n_1124), .Y(n_1060) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1061), .Y(n_1123) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_1062), .Y(n_1083) );
AND2x2_ASAP7_75t_SL g1062 ( .A(n_1063), .B(n_1075), .Y(n_1062) );
NOR3xp33_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1067), .C(n_1071), .Y(n_1063) );
OAI21xp33_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1069), .B(n_1070), .Y(n_1067) );
AND4x1_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1078), .C(n_1080), .D(n_1081), .Y(n_1075) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1085), .Y(n_1124) );
XOR2x2_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1103), .Y(n_1085) );
XOR2x2_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1102), .Y(n_1086) );
NAND4xp75_ASAP7_75t_SL g1087 ( .A(n_1088), .B(n_1097), .C(n_1100), .D(n_1101), .Y(n_1087) );
NOR2xp67_ASAP7_75t_SL g1088 ( .A(n_1089), .B(n_1093), .Y(n_1088) );
NAND3xp33_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1091), .C(n_1092), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1099), .Y(n_1097) );
XOR2x2_ASAP7_75t_SL g1103 ( .A(n_1104), .B(n_1122), .Y(n_1103) );
NAND2x1p5_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1114), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1111), .Y(n_1105) );
NAND3xp33_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1109), .C(n_1110), .Y(n_1106) );
NOR2x1_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1119), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1118), .Y(n_1115) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1117), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
INVx1_ASAP7_75t_SL g1127 ( .A(n_1128), .Y(n_1127) );
NOR2x1_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1133), .Y(n_1128) );
OR2x2_ASAP7_75t_SL g1191 ( .A(n_1129), .B(n_1134), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1132), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1130), .B(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1131), .B(n_1166), .Y(n_1194) );
CKINVDCx16_ASAP7_75t_R g1166 ( .A(n_1132), .Y(n_1166) );
CKINVDCx20_ASAP7_75t_R g1133 ( .A(n_1134), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1139), .Y(n_1137) );
OAI222xp33_ASAP7_75t_L g1140 ( .A1(n_1141), .A2(n_1165), .B1(n_1167), .B2(n_1187), .C1(n_1189), .C2(n_1192), .Y(n_1140) );
INVx1_ASAP7_75t_SL g1164 ( .A(n_1142), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1152), .Y(n_1142) );
NOR2xp33_ASAP7_75t_SL g1143 ( .A(n_1144), .B(n_1148), .Y(n_1143) );
NOR2xp33_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1157), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1155), .Y(n_1153) );
NAND2xp5_ASAP7_75t_SL g1157 ( .A(n_1158), .B(n_1161), .Y(n_1157) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1168), .Y(n_1188) );
AND4x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1176), .C(n_1181), .D(n_1186), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_1171), .A2(n_1172), .B1(n_1174), .B2(n_1175), .Y(n_1170) );
INVx1_ASAP7_75t_SL g1172 ( .A(n_1173), .Y(n_1172) );
CKINVDCx20_ASAP7_75t_R g1189 ( .A(n_1190), .Y(n_1189) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_1191), .Y(n_1190) );
CKINVDCx16_ASAP7_75t_R g1192 ( .A(n_1193), .Y(n_1192) );
endmodule