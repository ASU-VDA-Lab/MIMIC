module fake_jpeg_20888_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_22),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_10),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_20),
.B1(n_10),
.B2(n_16),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_18),
.B(n_25),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_20),
.B1(n_13),
.B2(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_38),
.C(n_40),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_41),
.B1(n_33),
.B2(n_26),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_28),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_29),
.C(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_33),
.B1(n_30),
.B2(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp67_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_15),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_46),
.B(n_35),
.Y(n_50)
);

OA21x2_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_30),
.B(n_15),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_14),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_37),
.C(n_17),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_46),
.B(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_14),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_19),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_56),
.C(n_17),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_42),
.C(n_19),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_58),
.B(n_60),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_4),
.C(n_5),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_1),
.B(n_3),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_6),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_55),
.A3(n_56),
.B1(n_17),
.B2(n_11),
.C1(n_14),
.C2(n_7),
.Y(n_64)
);

OAI21x1_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_60),
.B(n_58),
.Y(n_68)
);

XNOR2x2_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_6),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_7),
.B(n_9),
.Y(n_70)
);


endmodule