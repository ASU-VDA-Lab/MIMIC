module fake_jpeg_25188_n_181 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx11_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_29),
.B1(n_19),
.B2(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_31),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_24),
.B1(n_29),
.B2(n_28),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_52),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_25),
.B(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_45),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_29),
.B1(n_28),
.B2(n_20),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_48),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_51),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_10),
.B1(n_25),
.B2(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_56),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_36),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_11),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_41),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_74),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_44),
.C(n_51),
.Y(n_74)
);

XOR2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_44),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_23),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_35),
.B1(n_38),
.B2(n_36),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_79),
.B1(n_63),
.B2(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_53),
.B1(n_63),
.B2(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_23),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_64),
.B1(n_60),
.B2(n_66),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_88),
.B1(n_93),
.B2(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_91),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_35),
.B1(n_38),
.B2(n_46),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_54),
.B(n_1),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_12),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_12),
.Y(n_94)
);

OA21x2_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_12),
.B(n_17),
.Y(n_110)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_73),
.B1(n_78),
.B2(n_70),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_101),
.B1(n_42),
.B2(n_11),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_72),
.B1(n_42),
.B2(n_14),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_30),
.C(n_54),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_112),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_15),
.B(n_16),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_93),
.B(n_84),
.C(n_17),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_122),
.B(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_20),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_103),
.B(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_123),
.B(n_5),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_54),
.B1(n_11),
.B2(n_16),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_103),
.B1(n_102),
.B2(n_101),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_37),
.B1(n_21),
.B2(n_18),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_26),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_106),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_108),
.C(n_129),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_132),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_131),
.A2(n_137),
.B1(n_140),
.B2(n_117),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_106),
.B(n_98),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_127),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_123),
.B1(n_125),
.B2(n_128),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_105),
.B1(n_20),
.B2(n_37),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_20),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_30),
.C(n_21),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_141),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_114),
.B(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_145),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_148),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_27),
.B1(n_30),
.B2(n_7),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_150),
.A2(n_138),
.B1(n_141),
.B2(n_136),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_158),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_130),
.B(n_7),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_157),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_5),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_8),
.B(n_1),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_5),
.B(n_9),
.Y(n_157)
);

OAI21x1_ASAP7_75t_SL g158 ( 
.A1(n_150),
.A2(n_9),
.B(n_8),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_18),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_146),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_0),
.B(n_2),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_164),
.C(n_0),
.Y(n_171)
);

AOI21x1_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_151),
.B(n_8),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_151),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_13),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_160),
.B(n_3),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_170),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_13),
.B1(n_18),
.B2(n_3),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_171),
.A2(n_172),
.B(n_4),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_0),
.B(n_2),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_0),
.B(n_4),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_4),
.B(n_173),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_4),
.B(n_177),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_179),
.Y(n_181)
);


endmodule