module fake_jpeg_30565_n_289 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_11),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_8),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_19),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_60),
.B(n_61),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_41),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_26),
.B1(n_39),
.B2(n_17),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_65),
.A2(n_75),
.B1(n_34),
.B2(n_2),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_26),
.B1(n_20),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_72),
.B1(n_81),
.B2(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_70),
.B(n_77),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_26),
.B1(n_38),
.B2(n_36),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_17),
.B1(n_37),
.B2(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_73),
.A2(n_83),
.B1(n_92),
.B2(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_17),
.B1(n_37),
.B2(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_20),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_38),
.B(n_33),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.Y(n_121)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_29),
.B1(n_24),
.B2(n_37),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_30),
.B1(n_35),
.B2(n_23),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_53),
.A2(n_37),
.B1(n_33),
.B2(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_32),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_35),
.B1(n_30),
.B2(n_25),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_45),
.A2(n_35),
.B1(n_30),
.B2(n_25),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_25),
.B1(n_23),
.B2(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_45),
.A2(n_23),
.B1(n_32),
.B2(n_34),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_32),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_34),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_43),
.A2(n_21),
.B1(n_34),
.B2(n_3),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_56),
.B(n_9),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_10),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_43),
.A2(n_34),
.B1(n_7),
.B2(n_3),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_43),
.A2(n_34),
.B1(n_7),
.B2(n_3),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_107),
.A2(n_121),
.B(n_128),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_102),
.B1(n_80),
.B2(n_99),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_80),
.B1(n_94),
.B2(n_97),
.Y(n_138)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_119),
.Y(n_148)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_127),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_125),
.Y(n_169)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_135),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_75),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_5),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_12),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_151),
.B1(n_154),
.B2(n_156),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_63),
.B1(n_64),
.B2(n_94),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_169),
.B1(n_168),
.B2(n_148),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_87),
.B(n_61),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_143),
.B(n_141),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_66),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_163),
.C(n_111),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_63),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_152),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_106),
.A2(n_97),
.B1(n_64),
.B2(n_74),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_132),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_89),
.B1(n_71),
.B2(n_86),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_108),
.A2(n_89),
.B1(n_71),
.B2(n_86),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_74),
.B1(n_62),
.B2(n_68),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_161),
.B1(n_137),
.B2(n_150),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_62),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_140),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_109),
.A2(n_68),
.B1(n_13),
.B2(n_14),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_16),
.C(n_124),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_16),
.B(n_135),
.Y(n_164)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_166),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_111),
.B(n_134),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_130),
.B(n_114),
.C(n_133),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_114),
.B1(n_115),
.B2(n_123),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_115),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_114),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_177),
.Y(n_207)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

XNOR2x2_ASAP7_75t_SL g204 ( 
.A(n_176),
.B(n_189),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_167),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_178),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_162),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_125),
.B1(n_117),
.B2(n_118),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_190),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_122),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_187),
.B(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_126),
.B(n_125),
.C(n_122),
.D(n_113),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_157),
.A2(n_137),
.B1(n_150),
.B2(n_148),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_197),
.B(n_199),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_198),
.B1(n_144),
.B2(n_140),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_138),
.B1(n_139),
.B2(n_147),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_160),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_156),
.B1(n_154),
.B2(n_150),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_165),
.A2(n_143),
.B(n_166),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_208),
.B1(n_213),
.B2(n_193),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_144),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_216),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_198),
.A2(n_169),
.B1(n_139),
.B2(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_175),
.C(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_226),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_219),
.A2(n_192),
.B1(n_191),
.B2(n_183),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_225),
.Y(n_239)
);

XNOR2x2_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_176),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_236),
.B(n_238),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_218),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_175),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_235),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_171),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_231),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_181),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_234),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_183),
.B1(n_174),
.B2(n_176),
.Y(n_234)
);

AOI221xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_185),
.B1(n_197),
.B2(n_189),
.C(n_194),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_194),
.B1(n_197),
.B2(n_180),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_212),
.B(n_213),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_204),
.B(n_234),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_216),
.C(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_221),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_203),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_251),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_203),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_250),
.B(n_206),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_254),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_262),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_248),
.B1(n_222),
.B2(n_250),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_209),
.C(n_237),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_217),
.C(n_206),
.Y(n_265)
);

OAI31xp33_ASAP7_75t_L g263 ( 
.A1(n_256),
.A2(n_245),
.A3(n_242),
.B(n_239),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_249),
.A2(n_225),
.B1(n_238),
.B2(n_237),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_211),
.Y(n_268)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_243),
.C(n_249),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_200),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_242),
.B1(n_228),
.B2(n_204),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_205),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_204),
.B1(n_240),
.B2(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_230),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_258),
.C(n_217),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_255),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_273),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_253),
.B(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_263),
.A2(n_232),
.B1(n_226),
.B2(n_258),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_275),
.B(n_268),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_264),
.Y(n_280)
);

NAND2x1_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_270),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_277),
.B(n_281),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_284),
.B(n_280),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_282),
.C(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_285),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_278),
.Y(n_289)
);


endmodule