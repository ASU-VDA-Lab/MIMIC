module fake_jpeg_6263_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_37),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_45),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_27),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_12),
.C(n_20),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_21),
.B1(n_15),
.B2(n_28),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_15),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_14),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_73),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_28),
.B1(n_21),
.B2(n_15),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_71),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_44),
.B1(n_54),
.B2(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_12),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_22),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_21),
.B1(n_38),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_54),
.B1(n_14),
.B2(n_49),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_38),
.A3(n_24),
.B1(n_14),
.B2(n_26),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_43),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g79 ( 
.A(n_50),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_45),
.B1(n_44),
.B2(n_49),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_85),
.A2(n_99),
.B1(n_24),
.B2(n_26),
.Y(n_120)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_86),
.B(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_17),
.B1(n_68),
.B2(n_61),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_94),
.B1(n_97),
.B2(n_74),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_24),
.B(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_99),
.A2(n_62),
.B1(n_67),
.B2(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_106),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_76),
.C(n_59),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_94),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_108),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_75),
.B1(n_72),
.B2(n_46),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_117),
.Y(n_138)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_96),
.B(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_125),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_90),
.B(n_83),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_132),
.B(n_135),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_109),
.B1(n_111),
.B2(n_103),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_97),
.B(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_26),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

XOR2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_104),
.Y(n_139)
);

AOI321xp33_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_146),
.A3(n_150),
.B1(n_23),
.B2(n_19),
.C(n_3),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_116),
.C(n_105),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_115),
.B1(n_118),
.B2(n_107),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_148),
.A2(n_136),
.B(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_151),
.B(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_129),
.B(n_138),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_153),
.B(n_155),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_150),
.C(n_145),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_142),
.A3(n_144),
.B1(n_140),
.B2(n_147),
.C1(n_143),
.C2(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_157),
.B(n_19),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_24),
.C(n_26),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_23),
.C(n_4),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_23),
.C(n_10),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_1),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_165),
.B(n_1),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_1),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_158),
.B1(n_9),
.B2(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_167),
.B(n_169),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_23),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_168),
.C(n_8),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_171),
.Y(n_175)
);


endmodule