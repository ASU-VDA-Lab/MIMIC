module fake_netlist_5_651_n_1209 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1209);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1209;

wire n_924;
wire n_676;
wire n_431;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_615;
wire n_469;
wire n_851;
wire n_1060;
wire n_1141;
wire n_785;
wire n_855;
wire n_389;
wire n_843;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_605;
wire n_776;
wire n_928;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_620;
wire n_367;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_525;
wire n_397;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_372;
wire n_677;
wire n_443;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_1203;
wire n_821;
wire n_714;
wire n_447;
wire n_368;
wire n_433;
wire n_604;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1048;
wire n_932;
wire n_417;
wire n_946;
wire n_1008;
wire n_612;
wire n_1001;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_640;
wire n_559;
wire n_968;
wire n_624;
wire n_825;
wire n_1010;
wire n_877;
wire n_739;
wire n_508;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_1090;
wire n_1200;
wire n_633;
wire n_1192;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_1143;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_1182;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_579;
wire n_394;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_883;
wire n_1135;
wire n_752;
wire n_906;
wire n_905;
wire n_1163;
wire n_519;
wire n_406;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_918;
wire n_942;
wire n_381;
wire n_1147;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_618;
wire n_940;
wire n_896;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1172;
wire n_976;
wire n_1096;
wire n_1095;
wire n_379;
wire n_428;
wire n_570;
wire n_457;
wire n_514;
wire n_833;
wire n_1045;
wire n_1079;
wire n_1208;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_1201;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_795;
wire n_1009;
wire n_1148;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_1149;
wire n_882;
wire n_398;
wire n_1146;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_763;
wire n_522;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_1204;
wire n_580;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_670;
wire n_486;
wire n_816;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_1177;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_813;
wire n_1159;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_801;
wire n_369;
wire n_675;
wire n_888;
wire n_613;
wire n_871;
wire n_1119;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_517;
wire n_482;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_903;
wire n_1006;
wire n_740;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_1061;
wire n_477;
wire n_571;
wire n_461;
wire n_693;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_1193;
wire n_567;
wire n_1113;
wire n_652;
wire n_778;
wire n_1122;
wire n_1197;
wire n_1111;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_466;
wire n_1164;
wire n_420;
wire n_630;
wire n_1202;
wire n_632;
wire n_699;
wire n_489;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_1053;
wire n_1101;
wire n_585;
wire n_1106;
wire n_1190;
wire n_616;
wire n_953;
wire n_601;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_679;
wire n_513;
wire n_607;
wire n_407;
wire n_527;
wire n_425;
wire n_710;
wire n_707;
wire n_857;
wire n_695;
wire n_832;
wire n_1072;
wire n_560;
wire n_656;
wire n_1094;
wire n_561;
wire n_1044;
wire n_1205;
wire n_937;
wire n_393;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_1156;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_754;
wire n_712;
wire n_847;
wire n_1136;
wire n_815;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_529;
wire n_735;
wire n_702;
wire n_822;
wire n_412;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1160;
wire n_1080;
wire n_1162;
wire n_491;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1207;
wire n_1181;
wire n_1196;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_868;
wire n_803;
wire n_1092;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_1186;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_1189;
wire n_1029;
wire n_626;
wire n_925;
wire n_1180;
wire n_1206;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_784;

BUFx10_ASAP7_75t_L g354 ( 
.A(n_11),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_102),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_266),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_349),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_279),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_197),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_114),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_37),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_178),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_214),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_155),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_182),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_331),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_322),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_59),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_220),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_162),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_292),
.B(n_353),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_287),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_86),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_151),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_199),
.B(n_272),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_23),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_36),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_325),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_191),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_290),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_207),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_253),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_241),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_317),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_15),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_237),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_264),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_86),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_141),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_250),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_350),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_79),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_294),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_39),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_306),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_213),
.B(n_175),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_92),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_238),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_218),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_234),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_145),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_227),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_138),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_20),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_324),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_198),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_157),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_309),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_39),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_45),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_29),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_94),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_113),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_67),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_256),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_318),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_159),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_115),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_150),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_267),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_308),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_239),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_29),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_278),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_206),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_156),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_196),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_224),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_222),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_174),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_270),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_255),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_247),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_305),
.B(n_148),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_70),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_165),
.B(n_83),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_327),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_208),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_140),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_284),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_43),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_158),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_179),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_63),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_212),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_166),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_101),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_78),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_263),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_105),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_37),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_85),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_184),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_203),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_315),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_117),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_258),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_343),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_341),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_169),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_13),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_288),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_236),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_85),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_259),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_24),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_242),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_89),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_200),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_67),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_55),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_323),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_38),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_100),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_89),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_43),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_194),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_344),
.B(n_12),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_254),
.B(n_164),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_176),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_185),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_119),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_314),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_245),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_50),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_321),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_82),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_120),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_244),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_160),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_57),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_123),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_271),
.Y(n_499)
);

CKINVDCx14_ASAP7_75t_R g500 ( 
.A(n_276),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_171),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_269),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_289),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_152),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_248),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_71),
.Y(n_506)
);

INVxp33_ASAP7_75t_SL g507 ( 
.A(n_186),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_217),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_144),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_17),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_312),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_352),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_225),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_296),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_480),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_372),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_365),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_457),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_356),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_480),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_355),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_377),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_382),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_356),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_356),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_358),
.A2(n_361),
.B(n_359),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_400),
.B(n_0),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_491),
.B(n_1),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_393),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_356),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_365),
.B(n_2),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_474),
.B(n_2),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_391),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_426),
.B(n_3),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_357),
.B(n_3),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_391),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_391),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_357),
.B(n_421),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_403),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_421),
.B(n_4),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_470),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_426),
.B(n_5),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_500),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_470),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_410),
.Y(n_545)
);

OAI22x1_ASAP7_75t_L g546 ( 
.A1(n_474),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_473),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_388),
.A2(n_110),
.B(n_109),
.Y(n_548)
);

BUFx8_ASAP7_75t_SL g549 ( 
.A(n_479),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_429),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_423),
.A2(n_112),
.B(n_111),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_473),
.Y(n_553)
);

CKINVDCx6p67_ASAP7_75t_R g554 ( 
.A(n_354),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_473),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_460),
.B(n_13),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

AOI22x1_ASAP7_75t_SL g558 ( 
.A1(n_479),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_450),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_473),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_458),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_476),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_439),
.B(n_18),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_506),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_466),
.B(n_19),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_501),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_466),
.B(n_19),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_362),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_366),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_477),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_501),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_381),
.B(n_20),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_381),
.B(n_21),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_501),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_501),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_354),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_396),
.B(n_21),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_373),
.B(n_22),
.Y(n_580)
);

OA21x2_ASAP7_75t_L g581 ( 
.A1(n_367),
.A2(n_369),
.B(n_368),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_504),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_504),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_504),
.Y(n_584)
);

AOI22x1_ASAP7_75t_SL g585 ( 
.A1(n_415),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_363),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_511),
.Y(n_587)
);

OA21x2_ASAP7_75t_L g588 ( 
.A1(n_370),
.A2(n_25),
.B(n_26),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_442),
.B(n_25),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_544),
.B(n_420),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_519),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_582),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_582),
.Y(n_593)
);

CKINVDCx6p67_ASAP7_75t_R g594 ( 
.A(n_545),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_520),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_573),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_519),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_538),
.B(n_412),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_589),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_589),
.B(n_504),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_574),
.B(n_507),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_527),
.B(n_484),
.C(n_390),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_576),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_570),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_577),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_565),
.B(n_411),
.Y(n_606)
);

AND3x2_ASAP7_75t_L g607 ( 
.A(n_575),
.B(n_433),
.C(n_427),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_571),
.Y(n_608)
);

INVx8_ASAP7_75t_L g609 ( 
.A(n_537),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_517),
.B(n_483),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_557),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_564),
.B(n_580),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_521),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_531),
.B(n_475),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_532),
.Y(n_615)
);

BUFx6f_ASAP7_75t_SL g616 ( 
.A(n_531),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_586),
.Y(n_617)
);

AND3x2_ASAP7_75t_L g618 ( 
.A(n_528),
.B(n_451),
.C(n_449),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_519),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_524),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_524),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_525),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_587),
.B(n_511),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_522),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_580),
.B(n_467),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_525),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_525),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_525),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_530),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_526),
.B(n_452),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_530),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_552),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_581),
.B(n_495),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_631),
.B(n_581),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_613),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_601),
.B(n_578),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_612),
.A2(n_564),
.B(n_572),
.C(n_540),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_634),
.B(n_600),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_624),
.B(n_578),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_598),
.B(n_579),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_610),
.B(n_534),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_611),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_597),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_615),
.B(n_554),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_606),
.B(n_615),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_614),
.B(n_535),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_614),
.B(n_535),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_617),
.B(n_542),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_599),
.B(n_515),
.Y(n_651)
);

NOR3xp33_ASAP7_75t_L g652 ( 
.A(n_602),
.B(n_541),
.C(n_626),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_625),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_599),
.B(n_556),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_604),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_608),
.Y(n_656)
);

NOR3xp33_ASAP7_75t_L g657 ( 
.A(n_626),
.B(n_541),
.C(n_543),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_623),
.B(n_547),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_592),
.B(n_530),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_599),
.B(n_567),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_619),
.B(n_560),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_592),
.B(n_533),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_620),
.Y(n_663)
);

BUFx6f_ASAP7_75t_SL g664 ( 
.A(n_633),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_621),
.Y(n_665)
);

NAND2x1p5_ASAP7_75t_L g666 ( 
.A(n_595),
.B(n_588),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_593),
.B(n_533),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_590),
.B(n_569),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_596),
.B(n_398),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_596),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_593),
.B(n_533),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_603),
.B(n_398),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_605),
.B(n_533),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_622),
.B(n_513),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_622),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_627),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_627),
.B(n_536),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_616),
.B(n_409),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_628),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_628),
.B(n_536),
.Y(n_680)
);

INVx6_ASAP7_75t_L g681 ( 
.A(n_594),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_616),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_629),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_630),
.B(n_536),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_616),
.B(n_462),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_632),
.B(n_560),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_648),
.A2(n_649),
.B1(n_642),
.B2(n_640),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_670),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_651),
.B(n_594),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_647),
.B(n_650),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_637),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_636),
.B(n_632),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_640),
.A2(n_609),
.B(n_584),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_639),
.A2(n_562),
.B(n_550),
.C(n_559),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_665),
.Y(n_695)
);

CKINVDCx10_ASAP7_75t_R g696 ( 
.A(n_664),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_653),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_666),
.A2(n_551),
.B(n_548),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_652),
.A2(n_375),
.B(n_402),
.C(n_379),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_678),
.B(n_378),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_643),
.B(n_374),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_638),
.A2(n_588),
.B(n_440),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_644),
.B(n_654),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_660),
.A2(n_383),
.B1(n_485),
.B2(n_487),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_655),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_685),
.B(n_549),
.Y(n_706)
);

O2A1O1Ixp5_ASAP7_75t_L g707 ( 
.A1(n_641),
.A2(n_387),
.B(n_394),
.C(n_384),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_643),
.B(n_395),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_657),
.A2(n_499),
.B1(n_360),
.B2(n_364),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_646),
.B(n_550),
.Y(n_710)
);

INVx11_ASAP7_75t_L g711 ( 
.A(n_681),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_676),
.B(n_399),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_668),
.A2(n_546),
.B1(n_406),
.B2(n_407),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_669),
.B(n_549),
.Y(n_714)
);

CKINVDCx6p67_ASAP7_75t_R g715 ( 
.A(n_664),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_672),
.A2(n_562),
.B(n_529),
.C(n_561),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_682),
.A2(n_413),
.B1(n_414),
.B2(n_408),
.Y(n_717)
);

BUFx12f_ASAP7_75t_L g718 ( 
.A(n_681),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_656),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_663),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_679),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_674),
.B(n_397),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_675),
.B(n_607),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_683),
.Y(n_724)
);

AO21x2_ASAP7_75t_L g725 ( 
.A1(n_677),
.A2(n_431),
.B(n_430),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_680),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_680),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_635),
.A2(n_434),
.B(n_443),
.C(n_432),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_645),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_684),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_659),
.A2(n_667),
.B(n_662),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_673),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_673),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_659),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_662),
.B(n_472),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_667),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_671),
.Y(n_737)
);

NOR2x1_ASAP7_75t_L g738 ( 
.A(n_671),
.B(n_446),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_661),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_686),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_658),
.B(n_459),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_642),
.B(n_380),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_655),
.Y(n_743)
);

AO21x1_ASAP7_75t_L g744 ( 
.A1(n_648),
.A2(n_465),
.B(n_464),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_636),
.A2(n_496),
.B(n_494),
.Y(n_745)
);

AND2x6_ASAP7_75t_L g746 ( 
.A(n_636),
.B(n_503),
.Y(n_746)
);

BUFx4f_ASAP7_75t_SL g747 ( 
.A(n_638),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_669),
.B(n_523),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_655),
.Y(n_749)
);

AOI21x1_ASAP7_75t_L g750 ( 
.A1(n_636),
.A2(n_509),
.B(n_505),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_681),
.B(n_482),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_642),
.B(n_514),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_642),
.B(n_371),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_642),
.B(n_618),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_642),
.B(n_376),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_670),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_669),
.B(n_563),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_670),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_642),
.B(n_566),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_642),
.B(n_481),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_642),
.A2(n_539),
.B(n_386),
.C(n_389),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_636),
.A2(n_555),
.B(n_553),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_655),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_642),
.A2(n_513),
.B1(n_417),
.B2(n_418),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_642),
.B(n_385),
.Y(n_765)
);

AND2x6_ASAP7_75t_L g766 ( 
.A(n_727),
.B(n_730),
.Y(n_766)
);

O2A1O1Ixp5_ASAP7_75t_L g767 ( 
.A1(n_702),
.A2(n_518),
.B(n_516),
.C(n_392),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_691),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_697),
.Y(n_769)
);

OAI22x1_ASAP7_75t_L g770 ( 
.A1(n_714),
.A2(n_558),
.B1(n_585),
.B2(n_441),
.Y(n_770)
);

NOR2x1_ASAP7_75t_L g771 ( 
.A(n_690),
.B(n_493),
.Y(n_771)
);

OAI22x1_ASAP7_75t_L g772 ( 
.A1(n_742),
.A2(n_453),
.B1(n_456),
.B2(n_416),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_719),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_755),
.B(n_401),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_718),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_733),
.B(n_734),
.Y(n_776)
);

O2A1O1Ixp5_ASAP7_75t_L g777 ( 
.A1(n_699),
.A2(n_405),
.B(n_419),
.C(n_404),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_752),
.A2(n_424),
.B(n_425),
.C(n_422),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_692),
.A2(n_568),
.B(n_555),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_765),
.A2(n_435),
.B(n_436),
.C(n_428),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_731),
.A2(n_568),
.B(n_555),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_759),
.B(n_437),
.Y(n_782)
);

BUFx4f_ASAP7_75t_L g783 ( 
.A(n_715),
.Y(n_783)
);

AOI21xp33_ASAP7_75t_L g784 ( 
.A1(n_704),
.A2(n_510),
.B(n_497),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_710),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_756),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_736),
.A2(n_583),
.B(n_444),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_760),
.B(n_481),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_762),
.A2(n_750),
.B(n_739),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_689),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_705),
.Y(n_791)
);

AOI221xp5_ASAP7_75t_L g792 ( 
.A1(n_764),
.A2(n_448),
.B1(n_455),
.B2(n_445),
.C(n_438),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_746),
.A2(n_463),
.B(n_461),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_758),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_694),
.A2(n_469),
.B(n_471),
.C(n_468),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_722),
.Y(n_796)
);

NAND2x1p5_ASAP7_75t_L g797 ( 
.A(n_705),
.B(n_583),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_737),
.B(n_478),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_693),
.A2(n_118),
.B(n_116),
.Y(n_799)
);

OAI21x1_ASAP7_75t_L g800 ( 
.A1(n_695),
.A2(n_122),
.B(n_121),
.Y(n_800)
);

INVx5_ASAP7_75t_L g801 ( 
.A(n_746),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_726),
.A2(n_488),
.B(n_486),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_732),
.B(n_489),
.Y(n_803)
);

AND2x6_ASAP7_75t_SL g804 ( 
.A(n_706),
.B(n_26),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_753),
.B(n_490),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_703),
.A2(n_498),
.B(n_502),
.C(n_492),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_746),
.A2(n_512),
.B(n_508),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_705),
.B(n_124),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_724),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_720),
.Y(n_810)
);

OAI21xp33_ASAP7_75t_L g811 ( 
.A1(n_713),
.A2(n_27),
.B(n_28),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_746),
.A2(n_126),
.B(n_125),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_761),
.A2(n_128),
.B(n_127),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_735),
.B(n_30),
.Y(n_814)
);

AOI21x1_ASAP7_75t_L g815 ( 
.A1(n_741),
.A2(n_130),
.B(n_129),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_729),
.B(n_30),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_749),
.B(n_131),
.Y(n_817)
);

INVx5_ASAP7_75t_L g818 ( 
.A(n_763),
.Y(n_818)
);

AOI221x1_ASAP7_75t_SL g819 ( 
.A1(n_717),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.C(n_34),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_721),
.B(n_31),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_700),
.B(n_32),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_754),
.B(n_33),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_747),
.B(n_34),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_712),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_701),
.A2(n_133),
.B(n_132),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_708),
.A2(n_135),
.B(n_134),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_709),
.A2(n_137),
.B(n_136),
.Y(n_827)
);

AO31x2_ASAP7_75t_L g828 ( 
.A1(n_744),
.A2(n_38),
.A3(n_35),
.B(n_36),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_763),
.B(n_139),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_711),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_743),
.B(n_40),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_748),
.B(n_41),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_757),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_707),
.A2(n_143),
.B(n_146),
.C(n_142),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_763),
.B(n_147),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_751),
.B(n_41),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_740),
.B(n_42),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_716),
.B(n_44),
.Y(n_838)
);

AO21x2_ASAP7_75t_L g839 ( 
.A1(n_725),
.A2(n_153),
.B(n_149),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_738),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_723),
.B(n_154),
.Y(n_841)
);

INVx5_ASAP7_75t_L g842 ( 
.A(n_696),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_728),
.B(n_46),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_687),
.B(n_47),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_705),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_698),
.A2(n_163),
.B(n_161),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_687),
.B(n_47),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_687),
.B(n_48),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_742),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_849)
);

AO31x2_ASAP7_75t_L g850 ( 
.A1(n_744),
.A2(n_53),
.A3(n_51),
.B(n_52),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_745),
.A2(n_168),
.B(n_167),
.Y(n_851)
);

AOI21xp33_ASAP7_75t_L g852 ( 
.A1(n_742),
.A2(n_53),
.B(n_54),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_687),
.B(n_54),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_687),
.A2(n_172),
.B1(n_173),
.B2(n_170),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_698),
.A2(n_351),
.B(n_177),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_745),
.A2(n_181),
.B(n_180),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_760),
.B(n_55),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_687),
.B(n_56),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_698),
.A2(n_187),
.B(n_183),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_718),
.B(n_188),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_745),
.A2(n_190),
.B(n_189),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_688),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_687),
.B(n_56),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_745),
.A2(n_193),
.B(n_192),
.Y(n_864)
);

OAI22x1_ASAP7_75t_L g865 ( 
.A1(n_714),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_865)
);

NAND2x1p5_ASAP7_75t_L g866 ( 
.A(n_705),
.B(n_195),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_718),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_745),
.A2(n_202),
.B(n_201),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_745),
.A2(n_205),
.B(n_204),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_745),
.A2(n_210),
.B(n_209),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_760),
.B(n_60),
.Y(n_871)
);

NAND2x1p5_ASAP7_75t_L g872 ( 
.A(n_705),
.B(n_211),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_687),
.B(n_61),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_687),
.B(n_62),
.Y(n_874)
);

AOI211xp5_ASAP7_75t_L g875 ( 
.A1(n_742),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_875)
);

OA22x2_ASAP7_75t_L g876 ( 
.A1(n_760),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_691),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_742),
.A2(n_65),
.B(n_68),
.C(n_69),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_742),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_879)
);

AOI21xp33_ASAP7_75t_L g880 ( 
.A1(n_742),
.A2(n_71),
.B(n_72),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_851),
.A2(n_216),
.B(n_215),
.Y(n_881)
);

BUFx2_ASAP7_75t_SL g882 ( 
.A(n_818),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_785),
.B(n_72),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_775),
.B(n_73),
.Y(n_884)
);

AO21x2_ASAP7_75t_L g885 ( 
.A1(n_856),
.A2(n_221),
.B(n_219),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_796),
.B(n_73),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_773),
.B(n_74),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_789),
.A2(n_226),
.B(n_223),
.Y(n_888)
);

INVx6_ASAP7_75t_L g889 ( 
.A(n_818),
.Y(n_889)
);

BUFx12f_ASAP7_75t_L g890 ( 
.A(n_830),
.Y(n_890)
);

OAI21x1_ASAP7_75t_SL g891 ( 
.A1(n_861),
.A2(n_229),
.B(n_228),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_768),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_767),
.A2(n_231),
.B(n_230),
.Y(n_893)
);

AO21x2_ASAP7_75t_L g894 ( 
.A1(n_864),
.A2(n_233),
.B(n_232),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_867),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_781),
.A2(n_869),
.B(n_868),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_769),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_SL g898 ( 
.A1(n_822),
.A2(n_273),
.B(n_345),
.C(n_342),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_791),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_818),
.B(n_235),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_791),
.Y(n_901)
);

AOI21xp33_ASAP7_75t_L g902 ( 
.A1(n_844),
.A2(n_75),
.B(n_76),
.Y(n_902)
);

BUFx2_ASAP7_75t_SL g903 ( 
.A(n_791),
.Y(n_903)
);

INVx8_ASAP7_75t_L g904 ( 
.A(n_845),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_824),
.A2(n_275),
.B(n_340),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_846),
.A2(n_274),
.B(n_339),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_777),
.A2(n_277),
.B(n_338),
.Y(n_907)
);

OAI21x1_ASAP7_75t_SL g908 ( 
.A1(n_827),
.A2(n_268),
.B(n_337),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_855),
.A2(n_265),
.B(n_336),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_847),
.A2(n_280),
.B(n_335),
.Y(n_910)
);

OA21x2_ASAP7_75t_L g911 ( 
.A1(n_813),
.A2(n_262),
.B(n_334),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_782),
.B(n_77),
.Y(n_912)
);

AOI21xp33_ASAP7_75t_L g913 ( 
.A1(n_848),
.A2(n_77),
.B(n_78),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_814),
.B(n_79),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_853),
.A2(n_281),
.B(n_333),
.Y(n_915)
);

AO21x2_ASAP7_75t_L g916 ( 
.A1(n_826),
.A2(n_282),
.B(n_332),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_L g917 ( 
.A(n_821),
.B(n_80),
.C(n_81),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_836),
.B(n_80),
.C(n_81),
.Y(n_918)
);

OA21x2_ASAP7_75t_L g919 ( 
.A1(n_779),
.A2(n_283),
.B(n_330),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_859),
.A2(n_261),
.B(n_329),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_858),
.A2(n_260),
.B(n_328),
.Y(n_921)
);

AO21x2_ASAP7_75t_L g922 ( 
.A1(n_812),
.A2(n_257),
.B(n_326),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_783),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_863),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_788),
.B(n_84),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_877),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_810),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_790),
.B(n_87),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_771),
.B(n_88),
.Y(n_929)
);

AO21x1_ASAP7_75t_L g930 ( 
.A1(n_873),
.A2(n_88),
.B(n_90),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_786),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_841),
.B(n_240),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_783),
.Y(n_933)
);

AOI22x1_ASAP7_75t_L g934 ( 
.A1(n_772),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_833),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_799),
.A2(n_286),
.B(n_319),
.Y(n_936)
);

CKINVDCx11_ASAP7_75t_R g937 ( 
.A(n_804),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_809),
.Y(n_938)
);

AO21x2_ASAP7_75t_L g939 ( 
.A1(n_874),
.A2(n_252),
.B(n_316),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_774),
.A2(n_251),
.B(n_313),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_808),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_766),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_803),
.A2(n_249),
.B1(n_311),
.B2(n_310),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_829),
.Y(n_944)
);

BUFx6f_ASAP7_75t_SL g945 ( 
.A(n_841),
.Y(n_945)
);

NOR2x1_ASAP7_75t_SL g946 ( 
.A(n_801),
.B(n_246),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_857),
.B(n_93),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_800),
.A2(n_291),
.B(n_307),
.Y(n_948)
);

AO21x2_ASAP7_75t_L g949 ( 
.A1(n_870),
.A2(n_243),
.B(n_303),
.Y(n_949)
);

AO21x2_ASAP7_75t_L g950 ( 
.A1(n_780),
.A2(n_347),
.B(n_302),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_794),
.Y(n_951)
);

BUFx12f_ASAP7_75t_L g952 ( 
.A(n_842),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_862),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_842),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_811),
.A2(n_94),
.B(n_95),
.C(n_96),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_805),
.B(n_301),
.Y(n_956)
);

CKINVDCx11_ASAP7_75t_R g957 ( 
.A(n_842),
.Y(n_957)
);

INVx6_ASAP7_75t_L g958 ( 
.A(n_831),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_815),
.A2(n_300),
.B(n_299),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_871),
.B(n_95),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_766),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_866),
.Y(n_962)
);

CKINVDCx14_ASAP7_75t_R g963 ( 
.A(n_823),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_837),
.A2(n_298),
.B(n_297),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_860),
.B(n_295),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_832),
.B(n_96),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_834),
.A2(n_97),
.B(n_98),
.Y(n_967)
);

AND2x6_ASAP7_75t_L g968 ( 
.A(n_840),
.B(n_98),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_825),
.A2(n_99),
.B(n_102),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_798),
.A2(n_108),
.B(n_104),
.Y(n_970)
);

AOI22x1_ASAP7_75t_L g971 ( 
.A1(n_865),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_776),
.B(n_103),
.Y(n_972)
);

BUFx2_ASAP7_75t_R g973 ( 
.A(n_820),
.Y(n_973)
);

BUFx10_ASAP7_75t_L g974 ( 
.A(n_776),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_816),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_784),
.B(n_106),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_797),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_872),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_876),
.Y(n_979)
);

INVx5_ASAP7_75t_L g980 ( 
.A(n_801),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_787),
.A2(n_107),
.B(n_108),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_770),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_838),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_L g984 ( 
.A(n_792),
.B(n_875),
.C(n_852),
.Y(n_984)
);

AO21x2_ASAP7_75t_L g985 ( 
.A1(n_795),
.A2(n_778),
.B(n_793),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_854),
.A2(n_835),
.B(n_817),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_802),
.A2(n_807),
.B(n_843),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_828),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_806),
.B(n_880),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_828),
.Y(n_990)
);

INVx6_ASAP7_75t_L g991 ( 
.A(n_819),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_849),
.B(n_878),
.Y(n_992)
);

BUFx2_ASAP7_75t_R g993 ( 
.A(n_839),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_892),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_897),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_897),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_883),
.B(n_879),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_957),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_901),
.Y(n_999)
);

CKINVDCx11_ASAP7_75t_R g1000 ( 
.A(n_952),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_901),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_895),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_926),
.Y(n_1003)
);

OR2x6_ASAP7_75t_L g1004 ( 
.A(n_944),
.B(n_882),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_931),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_938),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_881),
.A2(n_984),
.B(n_989),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_889),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_974),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_941),
.B(n_850),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_927),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_979),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_951),
.Y(n_1013)
);

CKINVDCx11_ASAP7_75t_R g1014 ( 
.A(n_890),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_951),
.Y(n_1015)
);

AO21x1_ASAP7_75t_SL g1016 ( 
.A1(n_910),
.A2(n_921),
.B(n_915),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_954),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_928),
.B(n_925),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_976),
.A2(n_991),
.B1(n_971),
.B2(n_992),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_953),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_990),
.A2(n_988),
.B(n_983),
.Y(n_1021)
);

BUFx8_ASAP7_75t_L g1022 ( 
.A(n_945),
.Y(n_1022)
);

BUFx10_ASAP7_75t_L g1023 ( 
.A(n_945),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_889),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_906),
.A2(n_920),
.B(n_909),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_904),
.Y(n_1026)
);

AO21x2_ASAP7_75t_L g1027 ( 
.A1(n_893),
.A2(n_990),
.B(n_908),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_904),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_923),
.Y(n_1029)
);

CKINVDCx11_ASAP7_75t_R g1030 ( 
.A(n_937),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_901),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_963),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_935),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_942),
.B(n_980),
.Y(n_1034)
);

AOI221xp5_ASAP7_75t_L g1035 ( 
.A1(n_902),
.A2(n_913),
.B1(n_929),
.B2(n_886),
.C(n_917),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_960),
.B(n_975),
.Y(n_1036)
);

AO21x2_ASAP7_75t_L g1037 ( 
.A1(n_891),
.A2(n_907),
.B(n_987),
.Y(n_1037)
);

OAI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_991),
.A2(n_971),
.B1(n_918),
.B2(n_887),
.Y(n_1038)
);

CKINVDCx11_ASAP7_75t_R g1039 ( 
.A(n_884),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_966),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_899),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_955),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_934),
.A2(n_924),
.B1(n_930),
.B2(n_968),
.Y(n_1043)
);

NOR2x1_ASAP7_75t_SL g1044 ( 
.A(n_980),
.B(n_961),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_932),
.A2(n_912),
.B1(n_914),
.B2(n_947),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_903),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_958),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_972),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_958),
.Y(n_1049)
);

BUFx2_ASAP7_75t_SL g1050 ( 
.A(n_933),
.Y(n_1050)
);

OR2x6_ASAP7_75t_L g1051 ( 
.A(n_978),
.B(n_962),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_982),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_962),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_977),
.Y(n_1054)
);

NAND2x1p5_ASAP7_75t_L g1055 ( 
.A(n_965),
.B(n_986),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_934),
.A2(n_968),
.B1(n_970),
.B2(n_922),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_969),
.Y(n_1057)
);

OA21x2_ASAP7_75t_L g1058 ( 
.A1(n_967),
.A2(n_888),
.B(n_981),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_900),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_936),
.A2(n_948),
.B(n_959),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_884),
.Y(n_1061)
);

AO21x2_ASAP7_75t_L g1062 ( 
.A1(n_985),
.A2(n_885),
.B(n_894),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_968),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_922),
.A2(n_885),
.B1(n_894),
.B2(n_911),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_946),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_973),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_939),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1021),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1018),
.B(n_956),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_994),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_995),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_1024),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_997),
.B(n_964),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1036),
.B(n_950),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1012),
.B(n_950),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_1045),
.B(n_993),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_996),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_SL g1078 ( 
.A1(n_1067),
.A2(n_896),
.B1(n_916),
.B2(n_949),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1040),
.B(n_940),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1019),
.B(n_949),
.Y(n_1080)
);

AOI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_1035),
.A2(n_898),
.B(n_943),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1029),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1007),
.B(n_919),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1003),
.Y(n_1084)
);

NOR2x1_ASAP7_75t_L g1085 ( 
.A(n_1002),
.B(n_905),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1007),
.B(n_1048),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_1054),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1005),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1006),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1011),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1047),
.B(n_1049),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1047),
.B(n_1049),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_1033),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1038),
.A2(n_1016),
.B1(n_1043),
.B2(n_1042),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1013),
.B(n_1015),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1038),
.A2(n_1043),
.B1(n_1056),
.B2(n_1039),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1020),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_1051),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_1051),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1056),
.A2(n_1055),
.B(n_1065),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1067),
.A2(n_1051),
.B1(n_1064),
.B2(n_1052),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_SL g1102 ( 
.A1(n_1063),
.A2(n_1066),
.B1(n_1022),
.B2(n_1061),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1041),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1063),
.B(n_1055),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_1046),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1066),
.B(n_1053),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_1008),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1064),
.A2(n_1004),
.B1(n_1010),
.B2(n_1059),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1004),
.B(n_1050),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_1008),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_999),
.B(n_1031),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_1023),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_1023),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1044),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1001),
.B(n_1017),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1026),
.B(n_1028),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1098),
.B(n_1009),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1103),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1086),
.B(n_1027),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_1082),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1103),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1086),
.B(n_1027),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1070),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1071),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1068),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1077),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_1068),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1091),
.B(n_1057),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1092),
.B(n_1034),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1084),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_1082),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1088),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1076),
.A2(n_1032),
.B1(n_998),
.B2(n_1039),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1073),
.B(n_1062),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1072),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1076),
.A2(n_1032),
.B1(n_1037),
.B2(n_998),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1089),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1099),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1090),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1096),
.A2(n_1000),
.B1(n_1030),
.B2(n_1014),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1072),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1096),
.A2(n_1000),
.B1(n_1030),
.B2(n_1014),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1106),
.B(n_1058),
.Y(n_1143)
);

BUFx2_ASAP7_75t_SL g1144 ( 
.A(n_1110),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1094),
.B(n_1058),
.Y(n_1145)
);

AND2x4_ASAP7_75t_SL g1146 ( 
.A(n_1115),
.B(n_1025),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1069),
.B(n_1060),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1095),
.B(n_1074),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1097),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1087),
.Y(n_1150)
);

NOR2x1_ASAP7_75t_L g1151 ( 
.A(n_1085),
.B(n_1079),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1125),
.Y(n_1152)
);

NOR2xp67_ASAP7_75t_L g1153 ( 
.A(n_1131),
.B(n_1112),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1118),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1148),
.B(n_1080),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1134),
.B(n_1075),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1128),
.B(n_1093),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1121),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1149),
.B(n_1105),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1136),
.B(n_1081),
.C(n_1078),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1134),
.B(n_1083),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1123),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1143),
.B(n_1083),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1119),
.B(n_1122),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1129),
.B(n_1124),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1146),
.B(n_1100),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1126),
.B(n_1104),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1150),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1130),
.B(n_1101),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1132),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1137),
.B(n_1104),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1139),
.B(n_1095),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1164),
.B(n_1147),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1161),
.B(n_1156),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1162),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1167),
.B(n_1127),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1163),
.B(n_1145),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1152),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1165),
.B(n_1157),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1170),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1160),
.B(n_1136),
.C(n_1151),
.Y(n_1181)
);

NOR2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1169),
.B(n_1113),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1153),
.A2(n_1140),
.B(n_1142),
.Y(n_1183)
);

AOI33xp33_ASAP7_75t_L g1184 ( 
.A1(n_1154),
.A2(n_1142),
.A3(n_1140),
.B1(n_1102),
.B2(n_1078),
.B3(n_1133),
.Y(n_1184)
);

OAI21xp33_ASAP7_75t_L g1185 ( 
.A1(n_1184),
.A2(n_1102),
.B(n_1172),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1181),
.B(n_1184),
.C(n_1183),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1182),
.A2(n_1159),
.B(n_1138),
.C(n_1120),
.Y(n_1187)
);

AOI32xp33_ASAP7_75t_L g1188 ( 
.A1(n_1173),
.A2(n_1155),
.A3(n_1166),
.B1(n_1171),
.B2(n_1167),
.Y(n_1188)
);

OAI21xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1174),
.A2(n_1173),
.B(n_1177),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1186),
.A2(n_1166),
.B1(n_1179),
.B2(n_1176),
.Y(n_1190)
);

OAI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1185),
.A2(n_1180),
.B1(n_1175),
.B2(n_1141),
.C(n_1135),
.Y(n_1191)
);

AOI221xp5_ASAP7_75t_L g1192 ( 
.A1(n_1191),
.A2(n_1185),
.B1(n_1187),
.B2(n_1189),
.C(n_1188),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_L g1193 ( 
.A(n_1190),
.B(n_1178),
.C(n_1158),
.Y(n_1193)
);

NOR3xp33_ASAP7_75t_L g1194 ( 
.A(n_1192),
.B(n_1131),
.C(n_1109),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1193),
.B(n_1150),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1192),
.B(n_1150),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1195),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_SL g1198 ( 
.A(n_1196),
.B(n_1108),
.C(n_1114),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_1197),
.B(n_1198),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1199),
.B(n_1194),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1200),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1201),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1202),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1203),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1204),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1205),
.A2(n_1116),
.B(n_1107),
.Y(n_1206)
);

AOI21xp33_ASAP7_75t_SL g1207 ( 
.A1(n_1206),
.A2(n_1117),
.B(n_1111),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1207),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1208),
.A2(n_1144),
.B1(n_1168),
.B2(n_1117),
.Y(n_1209)
);


endmodule