module fake_jpeg_361_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_45),
.Y(n_58)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_67),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_45),
.B1(n_47),
.B2(n_41),
.Y(n_61)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_69),
.B1(n_62),
.B2(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_36),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_36),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_22),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_4),
.Y(n_98)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_40),
.B(n_37),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_6),
.B(n_7),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_64),
.B1(n_1),
.B2(n_2),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_96),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_82),
.B1(n_70),
.B2(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_98),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_3),
.CI(n_4),
.CON(n_96),
.SN(n_96)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_100),
.B(n_21),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_107),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_7),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_111),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_25),
.C(n_33),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_108),
.C(n_27),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_24),
.C(n_32),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_8),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_8),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_117),
.B1(n_101),
.B2(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_125),
.C(n_34),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_110),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_130),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_115),
.B(n_102),
.Y(n_132)
);

AO21x2_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_9),
.B(n_10),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_133),
.A2(n_119),
.B1(n_120),
.B2(n_125),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_120),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_139),
.B1(n_135),
.B2(n_137),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_126),
.B(n_122),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_124),
.B(n_14),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_13),
.C(n_18),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_19),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_20),
.Y(n_146)
);


endmodule