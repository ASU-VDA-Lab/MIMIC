module fake_netlist_1_5460_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_3), .B(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
NOR2x1p5_ASAP7_75t_L g16 ( .A(n_12), .B(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_13), .B(n_1), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_12), .B(n_14), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_15), .B(n_11), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_16), .Y(n_23) );
INVxp67_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVxp67_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OAI21xp33_ASAP7_75t_SL g27 ( .A1(n_25), .A2(n_21), .B(n_19), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_18), .B1(n_2), .B2(n_3), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_18), .B1(n_2), .B2(n_4), .Y(n_29) );
NAND5xp2_ASAP7_75t_L g30 ( .A(n_28), .B(n_1), .C(n_4), .D(n_5), .E(n_6), .Y(n_30) );
OR2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_6), .Y(n_31) );
INVx1_ASAP7_75t_SL g32 ( .A(n_27), .Y(n_32) );
INVx1_ASAP7_75t_SL g33 ( .A(n_31), .Y(n_33) );
HB1xp67_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
INVx2_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
AOI322xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_7), .A3(n_9), .B1(n_30), .B2(n_32), .C1(n_33), .C2(n_34), .Y(n_36) );
endmodule