module fake_netlist_1_11603_n_662 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_662);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_662;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_490;
wire n_247;
wire n_613;
wire n_393;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx5_ASAP7_75t_L g76 ( .A(n_62), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_41), .Y(n_77) );
INVxp33_ASAP7_75t_SL g78 ( .A(n_35), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_34), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_63), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_10), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_74), .Y(n_82) );
NOR2xp67_ASAP7_75t_L g83 ( .A(n_71), .B(n_0), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_72), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_20), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_16), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_1), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_3), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_65), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_7), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_50), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_54), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_49), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_22), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_11), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_18), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_55), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_67), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_47), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_27), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_29), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_37), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_42), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_58), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_53), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_9), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_19), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_5), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_60), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_7), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_8), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_28), .B(n_40), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_59), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_32), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_68), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_24), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_15), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_46), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_109), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_105), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_109), .B(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_79), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_105), .B(n_2), .Y(n_126) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_92), .B(n_75), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_76), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_89), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_90), .B(n_2), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_93), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_81), .B(n_3), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_76), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_86), .B(n_4), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_106), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_110), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_106), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_110), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_91), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_118), .B(n_10), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_80), .B(n_11), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_118), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_94), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_101), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_115), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_87), .B(n_12), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
AOI22x1_ASAP7_75t_SL g152 ( .A1(n_95), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_112), .B(n_13), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_116), .B(n_14), .Y(n_154) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_83), .A2(n_44), .B(n_17), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_76), .Y(n_156) );
INVx6_ASAP7_75t_L g157 ( .A(n_76), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_88), .B(n_16), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_107), .Y(n_159) );
INVxp67_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_112), .B(n_21), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_124), .B(n_76), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_124), .B(n_76), .Y(n_163) );
OAI22xp33_ASAP7_75t_SL g164 ( .A1(n_142), .A2(n_113), .B1(n_78), .B2(n_119), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_122), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_127), .B(n_117), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_128), .B(n_78), .Y(n_167) );
OAI22x1_ASAP7_75t_L g168 ( .A1(n_140), .A2(n_152), .B1(n_113), .B2(n_132), .Y(n_168) );
BUFx10_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_123), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_126), .B(n_114), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_128), .B(n_117), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_130), .B(n_98), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_130), .B(n_98), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_127), .B(n_77), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_123), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_126), .B(n_95), .Y(n_179) );
NOR2x1p5_ASAP7_75t_L g180 ( .A(n_132), .B(n_97), .Y(n_180) );
INVx4_ASAP7_75t_SL g181 ( .A(n_157), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_133), .B(n_84), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_123), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_160), .B(n_102), .Y(n_184) );
INVx5_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_133), .B(n_100), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_127), .B(n_99), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_146), .B(n_85), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_122), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_146), .B(n_96), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_143), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_122), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_147), .B(n_103), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_147), .B(n_103), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_148), .B(n_91), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_143), .Y(n_199) );
INVxp33_ASAP7_75t_SL g200 ( .A(n_144), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_148), .B(n_23), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_161), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_149), .B(n_25), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_126), .Y(n_205) );
NAND3xp33_ASAP7_75t_L g206 ( .A(n_150), .B(n_26), .C(n_30), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_150), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_126), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_149), .B(n_151), .Y(n_209) );
NAND2xp33_ASAP7_75t_R g210 ( .A(n_144), .B(n_31), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_151), .B(n_33), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_172), .B(n_154), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_172), .B(n_154), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_191), .A2(n_150), .B1(n_139), .B2(n_159), .Y(n_215) );
O2A1O1Ixp5_ASAP7_75t_L g216 ( .A1(n_205), .A2(n_156), .B(n_153), .C(n_137), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_205), .Y(n_217) );
OR2x2_ASAP7_75t_L g218 ( .A(n_195), .B(n_158), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_207), .B(n_156), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_212), .B(n_156), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_174), .B(n_156), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_169), .B(n_158), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_167), .B(n_137), .Y(n_224) );
BUFx3_ASAP7_75t_L g225 ( .A(n_189), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_174), .B(n_135), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_208), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_194), .B(n_135), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_170), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_204), .B(n_136), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_194), .B(n_157), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_190), .B(n_121), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_190), .B(n_121), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_166), .A2(n_142), .B1(n_140), .B2(n_152), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_173), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_176), .B(n_121), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g237 ( .A1(n_197), .A2(n_139), .B1(n_159), .B2(n_121), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_169), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_191), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_188), .B(n_139), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_188), .B(n_139), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_192), .A2(n_159), .B1(n_136), .B2(n_129), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_202), .B(n_136), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_177), .A2(n_125), .B1(n_129), .B2(n_159), .Y(n_244) );
O2A1O1Ixp5_ASAP7_75t_L g245 ( .A1(n_209), .A2(n_125), .B(n_129), .C(n_155), .Y(n_245) );
AND2x6_ASAP7_75t_SL g246 ( .A(n_179), .B(n_159), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_193), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_184), .B(n_125), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_182), .B(n_159), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_196), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_199), .B(n_145), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_186), .B(n_155), .Y(n_252) );
INVx4_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
NAND2x1_ASAP7_75t_L g254 ( .A(n_178), .B(n_155), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_183), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
INVx5_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
OR2x6_ASAP7_75t_L g258 ( .A(n_179), .B(n_155), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_187), .A2(n_145), .B1(n_141), .B2(n_134), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_171), .B(n_145), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g261 ( .A1(n_200), .A2(n_145), .B1(n_141), .B2(n_134), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_197), .B(n_145), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_171), .B(n_145), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_171), .B(n_141), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_171), .B(n_141), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_180), .A2(n_141), .B1(n_134), .B2(n_131), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_162), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_162), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_171), .B(n_141), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_206), .B(n_134), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_163), .B(n_175), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_217), .B(n_181), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_217), .Y(n_274) );
BUFx12f_ASAP7_75t_L g275 ( .A(n_238), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_218), .B(n_198), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_254), .A2(n_163), .B(n_185), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_217), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_224), .A2(n_211), .B(n_201), .C(n_131), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_234), .A2(n_210), .B1(n_134), .B2(n_131), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_223), .B(n_164), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g282 ( .A1(n_228), .A2(n_168), .B(n_134), .C(n_131), .Y(n_282) );
AOI21x1_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_270), .B(n_251), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_267), .B(n_175), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_213), .B(n_175), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_258), .A2(n_185), .B(n_131), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_258), .A2(n_185), .B(n_131), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_224), .A2(n_185), .B(n_38), .C(n_39), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_243), .Y(n_289) );
CKINVDCx11_ASAP7_75t_R g290 ( .A(n_246), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_227), .Y(n_291) );
CKINVDCx14_ASAP7_75t_R g292 ( .A(n_266), .Y(n_292) );
CKINVDCx8_ASAP7_75t_R g293 ( .A(n_262), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_226), .A2(n_36), .B(n_43), .C(n_45), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_268), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_245), .A2(n_48), .B(n_51), .Y(n_296) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_253), .B(n_52), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_239), .Y(n_299) );
AO32x1_ASAP7_75t_L g300 ( .A1(n_247), .A2(n_56), .A3(n_57), .B1(n_61), .B2(n_64), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_225), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_214), .B(n_66), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_232), .B(n_69), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_239), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_233), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_229), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_255), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_235), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_255), .B(n_70), .Y(n_309) );
OR2x6_ASAP7_75t_L g310 ( .A(n_253), .B(n_256), .Y(n_310) );
O2A1O1Ixp5_ASAP7_75t_SL g311 ( .A1(n_270), .A2(n_73), .B(n_251), .C(n_249), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_221), .B(n_240), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_253), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_219), .A2(n_220), .B(n_230), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_237), .B(n_225), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_241), .B(n_236), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_247), .Y(n_317) );
AO32x2_ASAP7_75t_L g318 ( .A1(n_216), .A2(n_262), .A3(n_264), .B1(n_263), .B2(n_265), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_231), .B(n_248), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_257), .B(n_219), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_230), .B(n_215), .Y(n_321) );
AO31x2_ASAP7_75t_L g322 ( .A1(n_280), .A2(n_260), .A3(n_269), .B(n_222), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_295), .B(n_220), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_272), .A2(n_222), .B(n_215), .Y(n_324) );
NAND3x1_ASAP7_75t_L g325 ( .A(n_281), .B(n_261), .C(n_259), .Y(n_325) );
OR2x6_ASAP7_75t_L g326 ( .A(n_275), .B(n_271), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_296), .A2(n_250), .B(n_242), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_276), .B(n_244), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g330 ( .A1(n_282), .A2(n_250), .B(n_242), .C(n_271), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_277), .A2(n_257), .B(n_302), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_312), .A2(n_257), .B(n_319), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_312), .A2(n_257), .B1(n_280), .B2(n_305), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_314), .A2(n_303), .B(n_279), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_316), .A2(n_289), .B(n_305), .C(n_315), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_283), .A2(n_311), .B(n_287), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_321), .A2(n_306), .B(n_308), .C(n_285), .Y(n_337) );
AOI221xp5_ASAP7_75t_SL g338 ( .A1(n_321), .A2(n_288), .B1(n_286), .B2(n_294), .C(n_304), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_290), .B(n_292), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_310), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g341 ( .A1(n_307), .A2(n_299), .B(n_291), .C(n_298), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_309), .A2(n_273), .B(n_284), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_320), .A2(n_297), .B(n_278), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_310), .B(n_317), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_274), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_274), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_300), .A2(n_318), .B(n_297), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_SL g349 ( .A1(n_278), .A2(n_318), .B(n_293), .C(n_300), .Y(n_349) );
AO31x2_ASAP7_75t_L g350 ( .A1(n_318), .A2(n_300), .A3(n_320), .B(n_313), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_313), .A2(n_252), .B(n_254), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_313), .B(n_295), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_272), .A2(n_252), .B(n_254), .Y(n_353) );
AO31x2_ASAP7_75t_L g354 ( .A1(n_333), .A2(n_334), .A3(n_353), .B(n_351), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_340), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_343), .A2(n_349), .B(n_333), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_344), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_343), .A2(n_331), .B(n_337), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_328), .B(n_335), .Y(n_359) );
BUFx2_ASAP7_75t_SL g360 ( .A(n_346), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_348), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_323), .A2(n_329), .B1(n_339), .B2(n_352), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_341), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_323), .B(n_325), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_338), .B(n_332), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_345), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_324), .B(n_342), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_347), .B(n_326), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g370 ( .A1(n_338), .A2(n_330), .B(n_348), .C(n_322), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_326), .A2(n_179), .B1(n_127), .B2(n_281), .Y(n_371) );
OA21x2_ASAP7_75t_L g372 ( .A1(n_322), .A2(n_350), .B(n_326), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_350), .A2(n_336), .B(n_343), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_350), .Y(n_374) );
AND2x6_ASAP7_75t_L g375 ( .A(n_322), .B(n_343), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_353), .A2(n_252), .B(n_334), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_337), .A2(n_335), .B(n_328), .C(n_282), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_327), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_352), .B(n_295), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_328), .A2(n_179), .B1(n_127), .B2(n_281), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_354), .B(n_374), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_370), .A2(n_376), .B(n_365), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_359), .B(n_364), .Y(n_383) );
HB1xp67_ASAP7_75t_SL g384 ( .A(n_360), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_368), .A2(n_356), .B(n_373), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_354), .B(n_374), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_359), .B(n_363), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_361), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_372), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_358), .A2(n_365), .B(n_378), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_363), .B(n_372), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_372), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_366), .A2(n_378), .B(n_377), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_372), .Y(n_394) );
AO21x2_ASAP7_75t_L g395 ( .A1(n_373), .A2(n_366), .B(n_369), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_360), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_361), .B(n_357), .Y(n_397) );
AO21x2_ASAP7_75t_L g398 ( .A1(n_354), .A2(n_375), .B(n_361), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_354), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_361), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_354), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_375), .Y(n_402) );
AO21x2_ASAP7_75t_L g403 ( .A1(n_375), .A2(n_379), .B(n_367), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_375), .A2(n_379), .B(n_367), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_375), .Y(n_405) );
OAI21x1_ASAP7_75t_L g406 ( .A1(n_375), .A2(n_355), .B(n_362), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_357), .B(n_371), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_375), .B(n_380), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_355), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_411), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_411), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_391), .B(n_381), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_387), .B(n_383), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_391), .B(n_381), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_397), .B(n_391), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_387), .B(n_383), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_411), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_397), .B(n_383), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_389), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_381), .B(n_386), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_384), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_381), .B(n_386), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_381), .B(n_386), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_405), .B(n_402), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_388), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_388), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_408), .A2(n_407), .B1(n_387), .B2(n_403), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_386), .B(n_399), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_400), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_386), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_386), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_396), .B(n_407), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_389), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_399), .B(n_401), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_408), .B(n_399), .Y(n_441) );
AND2x4_ASAP7_75t_SL g442 ( .A(n_384), .B(n_410), .Y(n_442) );
INVx5_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_405), .B(n_402), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_403), .B(n_404), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_408), .B(n_399), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_401), .B(n_398), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_392), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_389), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_407), .A2(n_403), .B1(n_404), .B2(n_410), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_405), .B(n_402), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_401), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_401), .B(n_398), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_382), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_439), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_439), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_419), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_421), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_426), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_414), .B(n_416), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
OAI21xp5_ASAP7_75t_SL g463 ( .A1(n_442), .A2(n_394), .B(n_410), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_415), .B(n_409), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_425), .B(n_394), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_425), .B(n_394), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_412), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_412), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_418), .B(n_404), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_442), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_413), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_422), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_413), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_413), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_452), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_414), .B(n_404), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_414), .B(n_404), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_442), .B(n_394), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_418), .B(n_404), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_424), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_425), .B(n_394), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_422), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_416), .B(n_403), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_424), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_416), .B(n_417), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_449), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_420), .B(n_403), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_452), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_417), .B(n_403), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_427), .B(n_392), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_438), .B(n_409), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_454), .B(n_409), .C(n_406), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_422), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_449), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_427), .B(n_398), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_420), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_447), .B(n_406), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_427), .B(n_398), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_443), .B(n_392), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
NOR2xp33_ASAP7_75t_SL g503 ( .A(n_443), .B(n_392), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_423), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_423), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_447), .B(n_406), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_428), .B(n_402), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_428), .B(n_398), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_428), .B(n_395), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_434), .B(n_395), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_456), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_456), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_487), .B(n_441), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_466), .B(n_453), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_502), .B(n_437), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_471), .B(n_437), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_457), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_490), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_487), .B(n_441), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_457), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_467), .B(n_446), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_459), .B(n_446), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_455), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_458), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_461), .B(n_434), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_461), .B(n_434), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_497), .B(n_453), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_496), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_464), .B(n_453), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_492), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_498), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_482), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_497), .B(n_454), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_460), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_465), .B(n_433), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_500), .B(n_454), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_496), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_477), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_477), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_500), .B(n_430), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_469), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_471), .B(n_436), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_472), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_490), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_470), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_470), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_508), .B(n_430), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_508), .B(n_436), .Y(n_551) );
NAND2x1_ASAP7_75t_L g552 ( .A(n_492), .B(n_448), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_493), .B(n_440), .Y(n_553) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_480), .B(n_443), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_504), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_481), .B(n_440), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_481), .B(n_448), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_463), .A2(n_406), .B(n_450), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_473), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_473), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_478), .B(n_445), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_491), .B(n_451), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_504), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_555), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_528), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_556), .B(n_489), .Y(n_566) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_554), .B(n_494), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_539), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_525), .B(n_492), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_511), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_511), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_532), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_533), .B(n_491), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_555), .Y(n_574) );
INVxp33_ASAP7_75t_L g575 ( .A(n_552), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_525), .B(n_466), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_552), .A2(n_503), .B1(n_489), .B2(n_445), .Y(n_577) );
AND2x2_ASAP7_75t_SL g578 ( .A(n_530), .B(n_478), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_535), .A2(n_495), .B(n_484), .C(n_474), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_533), .B(n_479), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_554), .B(n_443), .Y(n_581) );
OAI22xp33_ASAP7_75t_SL g582 ( .A1(n_554), .A2(n_501), .B1(n_443), .B2(n_483), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_545), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_538), .B(n_479), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_538), .B(n_485), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_534), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_536), .Y(n_587) );
AO21x1_ASAP7_75t_L g588 ( .A1(n_558), .A2(n_475), .B(n_476), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_526), .B(n_483), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_563), .Y(n_591) );
OAI222xp33_ASAP7_75t_L g592 ( .A1(n_530), .A2(n_485), .B1(n_499), .B2(n_506), .C1(n_443), .C2(n_466), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_537), .A2(n_509), .B1(n_510), .B2(n_507), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_557), .Y(n_594) );
OAI21xp33_ASAP7_75t_SL g595 ( .A1(n_526), .A2(n_509), .B(n_510), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_556), .B(n_483), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_557), .Y(n_597) );
NAND2xp33_ASAP7_75t_L g598 ( .A(n_530), .B(n_443), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_561), .A2(n_468), .B(n_507), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_523), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_524), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_564), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_583), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_564), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_595), .A2(n_553), .B1(n_521), .B2(n_529), .C(n_522), .Y(n_605) );
OAI21xp33_ASAP7_75t_SL g606 ( .A1(n_578), .A2(n_513), .B(n_519), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_594), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_594), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_565), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_601), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g611 ( .A1(n_575), .A2(n_514), .B(n_513), .C(n_519), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_600), .Y(n_612) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_579), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_566), .B(n_527), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_568), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_573), .B(n_527), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_570), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_571), .Y(n_618) );
AOI222xp33_ASAP7_75t_SL g619 ( .A1(n_597), .A2(n_512), .B1(n_517), .B2(n_520), .C1(n_540), .C2(n_541), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_572), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_593), .B(n_561), .Y(n_621) );
AOI322xp5_ASAP7_75t_L g622 ( .A1(n_578), .A2(n_542), .A3(n_550), .B1(n_551), .B2(n_562), .C1(n_514), .C2(n_468), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_SL g623 ( .A1(n_575), .A2(n_544), .B(n_516), .C(n_515), .Y(n_623) );
AOI21xp33_ASAP7_75t_SL g624 ( .A1(n_577), .A2(n_544), .B(n_516), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_608), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_606), .A2(n_567), .B(n_588), .C(n_582), .Y(n_626) );
OAI322xp33_ASAP7_75t_SL g627 ( .A1(n_621), .A2(n_580), .A3(n_584), .B1(n_585), .B2(n_590), .C1(n_587), .C2(n_586), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_623), .A2(n_598), .B(n_567), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_623), .A2(n_598), .B(n_581), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_617), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_613), .A2(n_577), .B(n_592), .C(n_581), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_605), .A2(n_593), .B1(n_599), .B2(n_514), .C(n_550), .Y(n_632) );
AOI322xp5_ASAP7_75t_L g633 ( .A1(n_613), .A2(n_569), .A3(n_576), .B1(n_589), .B2(n_551), .C1(n_542), .C2(n_468), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_603), .A2(n_507), .B1(n_596), .B2(n_429), .Y(n_634) );
AOI222xp33_ASAP7_75t_L g635 ( .A1(n_607), .A2(n_591), .B1(n_574), .B2(n_548), .C1(n_560), .C2(n_559), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_609), .B(n_591), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_611), .A2(n_515), .B1(n_574), .B2(n_549), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_611), .A2(n_543), .B(n_546), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g639 ( .A1(n_631), .A2(n_624), .B(n_612), .C(n_620), .Y(n_639) );
AOI322xp5_ASAP7_75t_L g640 ( .A1(n_632), .A2(n_610), .A3(n_615), .B1(n_622), .B2(n_619), .C1(n_618), .C2(n_604), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_627), .A2(n_604), .B1(n_602), .B2(n_614), .C(n_616), .Y(n_641) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_628), .A2(n_602), .B1(n_547), .B2(n_518), .Y(n_642) );
OAI211xp5_ASAP7_75t_L g643 ( .A1(n_626), .A2(n_518), .B(n_547), .C(n_563), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_625), .A2(n_476), .B1(n_475), .B2(n_451), .C1(n_444), .C2(n_429), .Y(n_644) );
AOI211xp5_ASAP7_75t_SL g645 ( .A1(n_629), .A2(n_390), .B(n_393), .C(n_451), .Y(n_645) );
AOI322xp5_ASAP7_75t_L g646 ( .A1(n_634), .A2(n_451), .A3(n_444), .B1(n_429), .B2(n_462), .C1(n_505), .C2(n_431), .Y(n_646) );
XNOR2x1_ASAP7_75t_L g647 ( .A(n_642), .B(n_637), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_640), .B(n_633), .C(n_638), .D(n_635), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_639), .B(n_630), .C(n_636), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_643), .B(n_390), .C(n_393), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_641), .A2(n_444), .B1(n_429), .B2(n_462), .C(n_505), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_648), .A2(n_645), .B1(n_644), .B2(n_646), .C(n_444), .Y(n_652) );
NOR2xp67_ASAP7_75t_SL g653 ( .A(n_649), .B(n_385), .Y(n_653) );
OAI21xp33_ASAP7_75t_L g654 ( .A1(n_647), .A2(n_423), .B(n_435), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_653), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_652), .Y(n_656) );
XOR2xp5_ASAP7_75t_L g657 ( .A(n_656), .B(n_650), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_657), .Y(n_658) );
OAI222xp33_ASAP7_75t_L g659 ( .A1(n_658), .A2(n_655), .B1(n_654), .B2(n_651), .C1(n_432), .C2(n_435), .Y(n_659) );
INVxp67_ASAP7_75t_L g660 ( .A(n_659), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g661 ( .A1(n_660), .A2(n_431), .B(n_435), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_661), .A2(n_382), .B1(n_385), .B2(n_395), .Y(n_662) );
endmodule