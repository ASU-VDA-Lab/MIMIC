module fake_ibex_810_n_3749 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_768, n_338, n_173, n_696, n_796, n_797, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_3749);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_768;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_3749;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3023;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3529;
wire n_1711;
wire n_3222;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_2252;
wire n_1982;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_3544;
wire n_2557;
wire n_2523;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3498;
wire n_2986;
wire n_3238;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_3385;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_3137;
wire n_2459;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_3337;
wire n_1263;
wire n_2465;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_961;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_991;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_3289;
wire n_2619;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_3512;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3493;
wire n_2447;
wire n_3044;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_3121;
wire n_2232;
wire n_2898;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2803;
wire n_2433;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_3102;
wire n_2872;
wire n_2790;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3543;
wire n_1734;
wire n_3143;
wire n_3655;
wire n_3742;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_3225;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_999;
wire n_2634;
wire n_2982;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3622;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2653;
wire n_2855;
wire n_2357;
wire n_2618;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2749;
wire n_888;
wire n_2378;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

BUFx10_ASAP7_75t_L g798 ( 
.A(n_88),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_96),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_156),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_77),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_613),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_402),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_726),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_409),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_137),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_573),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_47),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_609),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_735),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_101),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_449),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_209),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_709),
.Y(n_814)
);

BUFx10_ASAP7_75t_L g815 ( 
.A(n_469),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_229),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_379),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_719),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_544),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_579),
.B(n_330),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_164),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_520),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_510),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_60),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_763),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_194),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_643),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_787),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_174),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_230),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_442),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_603),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_203),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_503),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_785),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_510),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_260),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_545),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_360),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_223),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_788),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_375),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_212),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_686),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_272),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_406),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_782),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_603),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_574),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_580),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_570),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_598),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_256),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_175),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_688),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_16),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_382),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_309),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_512),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_225),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_624),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_795),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_391),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_126),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_281),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_379),
.Y(n_866)
);

BUFx5_ASAP7_75t_L g867 ( 
.A(n_503),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_228),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_29),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_740),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_13),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_354),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_55),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_131),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_343),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_255),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_575),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_756),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_714),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_206),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_728),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_449),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_368),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_264),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_252),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_171),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_698),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_308),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_242),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_277),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_780),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_484),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_519),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_265),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_548),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_369),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_566),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_581),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_319),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_267),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_288),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_293),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_57),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_40),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_562),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_513),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_581),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_464),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_188),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_548),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_27),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_1),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_240),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_555),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_710),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_403),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_312),
.Y(n_917)
);

CKINVDCx16_ASAP7_75t_R g918 ( 
.A(n_30),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_8),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_789),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_653),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_649),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_457),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_226),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_125),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_723),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_288),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_447),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_782),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_439),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_22),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_422),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_706),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_712),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_623),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_25),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_150),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_656),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_637),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_620),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_391),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_778),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_285),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_250),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_466),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_120),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_556),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_99),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_590),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_587),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_279),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_750),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_33),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_522),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_5),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_129),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_38),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_470),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_155),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_186),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_99),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_95),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_200),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_470),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_339),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_174),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_509),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_142),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_645),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_404),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_27),
.Y(n_971)
);

BUFx10_ASAP7_75t_L g972 ( 
.A(n_44),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_715),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_387),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_294),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_730),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_322),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_197),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_0),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_259),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_1),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_545),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_166),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_732),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_202),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_342),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_585),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_232),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_387),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_541),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_493),
.Y(n_991)
);

BUFx5_ASAP7_75t_L g992 ( 
.A(n_210),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_543),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_682),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_794),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_306),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_360),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_596),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_93),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_401),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_605),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_570),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_681),
.B(n_647),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_428),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_478),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_71),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_413),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_516),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_37),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_553),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_500),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_335),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_193),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_272),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_495),
.B(n_117),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_292),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_520),
.Y(n_1017)
);

BUFx10_ASAP7_75t_L g1018 ( 
.A(n_115),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_714),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_715),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_212),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_156),
.Y(n_1022)
);

INVxp67_ASAP7_75t_SL g1023 ( 
.A(n_489),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_611),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_458),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_340),
.Y(n_1026)
);

BUFx2_ASAP7_75t_SL g1027 ( 
.A(n_491),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_412),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_431),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_471),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_184),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_427),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_732),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_328),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_530),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_521),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_691),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_123),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_468),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_633),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_162),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_74),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_473),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_402),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_425),
.Y(n_1045)
);

NOR2xp67_ASAP7_75t_L g1046 ( 
.A(n_197),
.B(n_133),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_111),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_636),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_157),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_647),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_194),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_331),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_119),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_140),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_694),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_369),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_345),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_252),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_569),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_55),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_375),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_685),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_47),
.B(n_8),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_182),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_208),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_240),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_111),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_313),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_95),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_181),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_588),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_678),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_670),
.Y(n_1073)
);

BUFx2_ASAP7_75t_SL g1074 ( 
.A(n_772),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_602),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_264),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_410),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_724),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_152),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_514),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_64),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_14),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_112),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_141),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_552),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_692),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_249),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_640),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_679),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_628),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_678),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_357),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_323),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_275),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_703),
.Y(n_1095)
);

XNOR2x2_ASAP7_75t_R g1096 ( 
.A(n_365),
.B(n_584),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_412),
.Y(n_1097)
);

CKINVDCx14_ASAP7_75t_R g1098 ( 
.A(n_120),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_452),
.Y(n_1099)
);

BUFx10_ASAP7_75t_L g1100 ( 
.A(n_741),
.Y(n_1100)
);

BUFx5_ASAP7_75t_L g1101 ( 
.A(n_672),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_580),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_537),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_646),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_251),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_774),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_160),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_512),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_164),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_504),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_18),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_406),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_430),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_749),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_83),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_632),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_150),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_38),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_242),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_192),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_0),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_437),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_376),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_525),
.Y(n_1124)
);

BUFx10_ASAP7_75t_L g1125 ( 
.A(n_421),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_546),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_529),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_514),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_767),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_208),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_330),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_118),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_389),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_619),
.Y(n_1134)
);

BUFx5_ASAP7_75t_L g1135 ( 
.A(n_454),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_467),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_481),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_661),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_129),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_228),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_98),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_724),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_502),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_441),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_543),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_654),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_344),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_424),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_568),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_625),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_184),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_100),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_26),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_274),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_632),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_516),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_485),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_590),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_45),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_144),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_58),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_558),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_70),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_673),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_312),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_201),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_128),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_215),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_597),
.Y(n_1169)
);

CKINVDCx16_ASAP7_75t_R g1170 ( 
.A(n_236),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_163),
.Y(n_1171)
);

CKINVDCx16_ASAP7_75t_R g1172 ( 
.A(n_68),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_496),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_705),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_628),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_657),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_115),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_690),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_36),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_338),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_539),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_586),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_147),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_610),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_343),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_190),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_867),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1098),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1098),
.A2(n_909),
.B1(n_1043),
.B2(n_850),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_863),
.B(n_2),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_850),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_883),
.B(n_2),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_798),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_798),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_909),
.Y(n_1195)
);

BUFx8_ASAP7_75t_SL g1196 ( 
.A(n_800),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_812),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1043),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_905),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_893),
.B(n_3),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1107),
.Y(n_1201)
);

CKINVDCx6p67_ASAP7_75t_R g1202 ( 
.A(n_798),
.Y(n_1202)
);

CKINVDCx16_ASAP7_75t_R g1203 ( 
.A(n_869),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1166),
.B(n_1171),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_906),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1107),
.B(n_6),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_815),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1136),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_841),
.A2(n_791),
.B(n_790),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_918),
.B(n_6),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_815),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_839),
.A2(n_793),
.B(n_792),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_867),
.Y(n_1213)
);

BUFx12f_ASAP7_75t_L g1214 ( 
.A(n_815),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_867),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_933),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1136),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_839),
.A2(n_797),
.B(n_796),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_972),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_972),
.Y(n_1220)
);

BUFx8_ASAP7_75t_SL g1221 ( 
.A(n_800),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1036),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_867),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_972),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_814),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_867),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_812),
.Y(n_1227)
);

BUFx8_ASAP7_75t_SL g1228 ( 
.A(n_827),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_856),
.B(n_7),
.Y(n_1229)
);

CKINVDCx6p67_ASAP7_75t_R g1230 ( 
.A(n_1018),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_998),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_SL g1232 ( 
.A(n_920),
.B(n_9),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_856),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1054),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1185),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_812),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_857),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_857),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_914),
.B(n_10),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_914),
.B(n_11),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_867),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_992),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_932),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_992),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_803),
.B(n_12),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1160),
.B(n_1170),
.Y(n_1246)
);

BUFx8_ASAP7_75t_SL g1247 ( 
.A(n_827),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_932),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_962),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_992),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_992),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1172),
.A2(n_823),
.B1(n_824),
.B2(n_822),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_831),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_992),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_962),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_822),
.B(n_823),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_992),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1018),
.Y(n_1258)
);

AOI22x1_ASAP7_75t_SL g1259 ( 
.A1(n_831),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_824),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_992),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_826),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1018),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1069),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1101),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1090),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1101),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1090),
.Y(n_1268)
);

INVx6_ASAP7_75t_L g1269 ( 
.A(n_1069),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_812),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1157),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_826),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1101),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_828),
.B(n_18),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1157),
.B(n_17),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_SL g1276 ( 
.A1(n_834),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_828),
.B(n_20),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1182),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_829),
.B(n_21),
.Y(n_1279)
);

BUFx8_ASAP7_75t_L g1280 ( 
.A(n_1063),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_829),
.B(n_23),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1069),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1182),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1101),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_825),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1101),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_830),
.A2(n_786),
.B1(n_787),
.B2(n_785),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_843),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1100),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1100),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1260),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1283),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1193),
.B(n_920),
.Y(n_1293)
);

INVxp67_ASAP7_75t_SL g1294 ( 
.A(n_1199),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1238),
.B(n_1101),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1212),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1269),
.Y(n_1297)
);

CKINVDCx6p67_ASAP7_75t_R g1298 ( 
.A(n_1211),
.Y(n_1298)
);

INVx5_ASAP7_75t_L g1299 ( 
.A(n_1229),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1229),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1275),
.B(n_1101),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1238),
.B(n_1135),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1204),
.B(n_1180),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1227),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1285),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1269),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1285),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1205),
.B(n_1100),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1285),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1275),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1269),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1243),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1187),
.B(n_1135),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1187),
.B(n_1135),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1266),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1213),
.B(n_1135),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1213),
.B(n_1135),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1211),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1215),
.B(n_1135),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1223),
.B(n_862),
.Y(n_1320)
);

NAND2xp33_ASAP7_75t_SL g1321 ( 
.A(n_1188),
.B(n_1210),
.Y(n_1321)
);

AND3x2_ASAP7_75t_L g1322 ( 
.A(n_1232),
.B(n_1096),
.C(n_1023),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1223),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1239),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1214),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1226),
.B(n_995),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1240),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1226),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1241),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1241),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1242),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1242),
.B(n_825),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1260),
.Y(n_1333)
);

AO21x2_ASAP7_75t_L g1334 ( 
.A1(n_1218),
.A2(n_802),
.B(n_801),
.Y(n_1334)
);

AOI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1244),
.A2(n_853),
.B(n_843),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1250),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1191),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1250),
.B(n_825),
.Y(n_1338)
);

NAND2xp33_ASAP7_75t_L g1339 ( 
.A(n_1188),
.B(n_825),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1195),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1251),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1253),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1254),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1193),
.B(n_799),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1216),
.B(n_1125),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1254),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1257),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1194),
.B(n_1207),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1257),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1272),
.A2(n_832),
.B1(n_833),
.B2(n_830),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1222),
.B(n_1125),
.Y(n_1351)
);

CKINVDCx16_ASAP7_75t_R g1352 ( 
.A(n_1203),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1214),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1272),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1261),
.Y(n_1355)
);

AND3x2_ASAP7_75t_L g1356 ( 
.A(n_1234),
.B(n_1235),
.C(n_1199),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1261),
.B(n_854),
.Y(n_1357)
);

BUFx10_ASAP7_75t_L g1358 ( 
.A(n_1258),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1201),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1196),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1265),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1208),
.Y(n_1362)
);

AND2x6_ASAP7_75t_L g1363 ( 
.A(n_1189),
.B(n_854),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1246),
.B(n_1176),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1265),
.Y(n_1365)
);

INVx6_ASAP7_75t_L g1366 ( 
.A(n_1263),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1217),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1197),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1225),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1263),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1267),
.B(n_854),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1267),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1273),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1194),
.B(n_805),
.Y(n_1374)
);

BUFx4f_ASAP7_75t_L g1375 ( 
.A(n_1202),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1273),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1233),
.Y(n_1377)
);

AND2x2_ASAP7_75t_SL g1378 ( 
.A(n_1190),
.B(n_1015),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1237),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1284),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1248),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1207),
.B(n_806),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1249),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1284),
.Y(n_1384)
);

INVxp33_ASAP7_75t_SL g1385 ( 
.A(n_1252),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1286),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1255),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1264),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1230),
.B(n_1125),
.Y(n_1389)
);

NOR2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1264),
.B(n_1180),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1268),
.Y(n_1391)
);

AND3x2_ASAP7_75t_L g1392 ( 
.A(n_1192),
.B(n_1200),
.C(n_1278),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1271),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1288),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1256),
.B(n_833),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1219),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1219),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1220),
.Y(n_1398)
);

BUFx10_ASAP7_75t_L g1399 ( 
.A(n_1245),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_SL g1400 ( 
.A(n_1196),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1224),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1224),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1282),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1289),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1289),
.B(n_853),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1197),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1236),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_L g1408 ( 
.A(n_1290),
.B(n_916),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1236),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1290),
.B(n_1280),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1280),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1209),
.B(n_916),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1236),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1270),
.Y(n_1414)
);

NOR2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1221),
.B(n_832),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1270),
.B(n_895),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1270),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1270),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1274),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1277),
.B(n_895),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1279),
.B(n_1281),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1198),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1231),
.B(n_1173),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1262),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1287),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1276),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1259),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1221),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1253),
.A2(n_836),
.B1(n_838),
.B2(n_835),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1228),
.B(n_1014),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1228),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1247),
.B(n_807),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1247),
.Y(n_1433)
);

AND2x6_ASAP7_75t_L g1434 ( 
.A(n_1229),
.B(n_968),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1206),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1283),
.Y(n_1436)
);

NAND2xp33_ASAP7_75t_SL g1437 ( 
.A(n_1188),
.B(n_968),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1205),
.B(n_835),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1206),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1229),
.B(n_968),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1199),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1283),
.Y(n_1442)
);

NAND2xp33_ASAP7_75t_L g1443 ( 
.A(n_1188),
.B(n_978),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1206),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1206),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1206),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1283),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1206),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1231),
.A2(n_844),
.B1(n_861),
.B2(n_834),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1441),
.B(n_836),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1297),
.B(n_808),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1306),
.B(n_813),
.Y(n_1452)
);

NOR2xp67_ASAP7_75t_L g1453 ( 
.A(n_1299),
.B(n_912),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1419),
.B(n_1421),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1421),
.B(n_838),
.Y(n_1455)
);

NOR3xp33_ASAP7_75t_L g1456 ( 
.A(n_1449),
.B(n_837),
.C(n_818),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1294),
.B(n_1181),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1293),
.B(n_1173),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1441),
.B(n_1175),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1420),
.B(n_1175),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1397),
.B(n_819),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1395),
.B(n_1176),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1396),
.B(n_846),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1366),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1294),
.B(n_1303),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1348),
.B(n_1177),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1399),
.B(n_1025),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1366),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1348),
.B(n_1177),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1438),
.B(n_1308),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1292),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1366),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1398),
.B(n_1401),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1402),
.B(n_1181),
.Y(n_1474)
);

BUFx5_ASAP7_75t_L g1475 ( 
.A(n_1434),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1403),
.B(n_1183),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1404),
.B(n_1183),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1337),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1291),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1344),
.B(n_848),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1433),
.B(n_1411),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1436),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1344),
.B(n_849),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1374),
.B(n_1184),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1374),
.B(n_858),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1340),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1375),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1382),
.B(n_1184),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1359),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1345),
.B(n_866),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1364),
.B(n_868),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1312),
.B(n_873),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1362),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1333),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1439),
.B(n_875),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1367),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1315),
.B(n_876),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1435),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1311),
.B(n_878),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1435),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1444),
.B(n_1446),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1351),
.B(n_880),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1445),
.Y(n_1503)
);

BUFx5_ASAP7_75t_L g1504 ( 
.A(n_1434),
.Y(n_1504)
);

NOR3xp33_ASAP7_75t_L g1505 ( 
.A(n_1449),
.B(n_882),
.C(n_842),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1298),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1442),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1324),
.B(n_884),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1378),
.B(n_885),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1327),
.B(n_888),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1300),
.B(n_1038),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1296),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1352),
.B(n_896),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1311),
.B(n_890),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1445),
.Y(n_1515)
);

INVx8_ASAP7_75t_L g1516 ( 
.A(n_1434),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1448),
.B(n_892),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1447),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1422),
.A2(n_942),
.B1(n_951),
.B2(n_931),
.C(n_904),
.Y(n_1519)
);

AND2x2_ASAP7_75t_SL g1520 ( 
.A(n_1375),
.B(n_945),
.Y(n_1520)
);

INVx8_ASAP7_75t_L g1521 ( 
.A(n_1434),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1335),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1429),
.B(n_958),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1448),
.B(n_901),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1394),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1387),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1358),
.B(n_902),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1342),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1425),
.A2(n_810),
.B1(n_811),
.B2(n_809),
.C(n_804),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1388),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1310),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1405),
.B(n_1295),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1299),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1299),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1422),
.A2(n_817),
.B1(n_821),
.B2(n_816),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1369),
.Y(n_1536)
);

INVx4_ASAP7_75t_L g1537 ( 
.A(n_1358),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1318),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1295),
.B(n_907),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1377),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1302),
.B(n_908),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1379),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1381),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1304),
.Y(n_1544)
);

INVxp67_ASAP7_75t_L g1545 ( 
.A(n_1354),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1325),
.B(n_910),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1353),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1370),
.B(n_913),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1302),
.B(n_915),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1378),
.B(n_921),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1437),
.B(n_1077),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1383),
.B(n_922),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1389),
.B(n_923),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1410),
.B(n_925),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1305),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1356),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1391),
.B(n_1393),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1301),
.B(n_926),
.Y(n_1558)
);

BUFx8_ASAP7_75t_L g1559 ( 
.A(n_1400),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1350),
.B(n_1093),
.Y(n_1560)
);

BUFx8_ASAP7_75t_L g1561 ( 
.A(n_1400),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1410),
.B(n_928),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1440),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1320),
.B(n_929),
.Y(n_1564)
);

INVxp33_ASAP7_75t_L g1565 ( 
.A(n_1430),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1416),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1307),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1385),
.B(n_930),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1309),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1356),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1320),
.B(n_934),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_SL g1572 ( 
.A(n_1433),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1363),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1416),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1385),
.B(n_935),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1326),
.B(n_937),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1363),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1334),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1326),
.B(n_938),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1412),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1334),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1322),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1363),
.B(n_939),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1424),
.A2(n_840),
.B1(n_847),
.B2(n_845),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1423),
.B(n_964),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1321),
.B(n_1093),
.Y(n_1586)
);

A2O1A1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1425),
.A2(n_851),
.B(n_855),
.C(n_852),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1321),
.B(n_1093),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1363),
.B(n_940),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1363),
.B(n_941),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1392),
.B(n_943),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1392),
.B(n_944),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1408),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1412),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1339),
.B(n_947),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1339),
.B(n_952),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1323),
.B(n_953),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_SL g1598 ( 
.A(n_1428),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1443),
.B(n_954),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1390),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1328),
.B(n_960),
.Y(n_1601)
);

INVx8_ASAP7_75t_L g1602 ( 
.A(n_1360),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1342),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1443),
.B(n_961),
.Y(n_1604)
);

NOR3xp33_ASAP7_75t_L g1605 ( 
.A(n_1426),
.B(n_977),
.C(n_971),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1332),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1432),
.B(n_963),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1313),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1432),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1329),
.B(n_976),
.Y(n_1610)
);

AND2x6_ASAP7_75t_L g1611 ( 
.A(n_1426),
.B(n_945),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1314),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1427),
.A2(n_982),
.B1(n_983),
.B2(n_980),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1332),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1329),
.B(n_985),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1330),
.B(n_986),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1330),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1314),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1331),
.B(n_987),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1336),
.B(n_994),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1338),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1338),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1431),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1316),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_L g1625 ( 
.A(n_1316),
.B(n_999),
.C(n_997),
.Y(n_1625)
);

NAND2x1_ASAP7_75t_L g1626 ( 
.A(n_1341),
.B(n_1016),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1322),
.B(n_1001),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1343),
.B(n_1002),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1346),
.B(n_1005),
.Y(n_1629)
);

NOR2xp67_ASAP7_75t_L g1630 ( 
.A(n_1317),
.B(n_1017),
.Y(n_1630)
);

INVx8_ASAP7_75t_L g1631 ( 
.A(n_1407),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1347),
.B(n_1008),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1349),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1357),
.Y(n_1634)
);

NAND2xp33_ASAP7_75t_L g1635 ( 
.A(n_1355),
.B(n_1113),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1319),
.A2(n_859),
.B(n_864),
.C(n_860),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1415),
.A2(n_871),
.B1(n_872),
.B2(n_870),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1361),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1365),
.B(n_1010),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1372),
.B(n_1133),
.Y(n_1640)
);

BUFx5_ASAP7_75t_L g1641 ( 
.A(n_1371),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1371),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1373),
.B(n_1011),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1376),
.A2(n_1019),
.B1(n_1020),
.B2(n_1013),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1380),
.B(n_1021),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1384),
.B(n_1386),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1407),
.B(n_1133),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1414),
.B(n_1022),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1407),
.B(n_1133),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1407),
.B(n_1024),
.Y(n_1650)
);

AOI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1406),
.A2(n_886),
.B1(n_887),
.B2(n_879),
.C(n_877),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1418),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1418),
.B(n_1031),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1368),
.B(n_1163),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1409),
.B(n_1032),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1368),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_SL g1657 ( 
.A(n_1368),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1413),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1417),
.A2(n_891),
.B1(n_894),
.B2(n_889),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1297),
.B(n_1033),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1454),
.A2(n_897),
.B(n_899),
.C(n_898),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1631),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1537),
.B(n_820),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1532),
.A2(n_903),
.B(n_900),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1530),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1457),
.B(n_1034),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1522),
.A2(n_1581),
.B(n_1578),
.Y(n_1667)
);

NOR2xp67_ASAP7_75t_L g1668 ( 
.A(n_1556),
.B(n_19),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1465),
.B(n_844),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1479),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1455),
.B(n_1035),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1587),
.A2(n_917),
.B(n_919),
.C(n_911),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1498),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1460),
.B(n_1039),
.Y(n_1674)
);

CKINVDCx10_ASAP7_75t_R g1675 ( 
.A(n_1572),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1494),
.B(n_861),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1450),
.A2(n_874),
.B1(n_881),
.B2(n_865),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1545),
.B(n_865),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1501),
.A2(n_936),
.B(n_927),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1633),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1566),
.A2(n_948),
.B(n_946),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1608),
.A2(n_950),
.B(n_949),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1459),
.B(n_1509),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1537),
.B(n_1042),
.Y(n_1684)
);

OAI321xp33_ASAP7_75t_L g1685 ( 
.A1(n_1519),
.A2(n_1584),
.A3(n_957),
.B1(n_955),
.B2(n_965),
.C(n_956),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1538),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1612),
.A2(n_1624),
.B(n_1618),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1631),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1478),
.A2(n_881),
.B1(n_924),
.B2(n_874),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1633),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1486),
.A2(n_1493),
.B1(n_1496),
.B2(n_1489),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1547),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1643),
.B(n_1047),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1646),
.A2(n_1557),
.B(n_1541),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1539),
.A2(n_967),
.B(n_966),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1506),
.Y(n_1696)
);

O2A1O1Ixp33_ASAP7_75t_L g1697 ( 
.A1(n_1456),
.A2(n_970),
.B(n_973),
.C(n_969),
.Y(n_1697)
);

AO21x1_ASAP7_75t_L g1698 ( 
.A1(n_1586),
.A2(n_975),
.B(n_974),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1536),
.A2(n_981),
.B(n_984),
.C(n_979),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1611),
.A2(n_1074),
.B1(n_1027),
.B2(n_959),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1500),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1549),
.A2(n_1473),
.B(n_1495),
.Y(n_1702)
);

A2O1A1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1540),
.A2(n_991),
.B(n_993),
.C(n_989),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1645),
.B(n_1491),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1638),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1563),
.A2(n_1004),
.B(n_1000),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1462),
.B(n_1048),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1574),
.A2(n_1007),
.B(n_1006),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1531),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1558),
.A2(n_1012),
.B(n_1009),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1480),
.B(n_1483),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1550),
.B(n_924),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1503),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1515),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1559),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1568),
.A2(n_1051),
.B1(n_1052),
.B2(n_1049),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1464),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_L g1718 ( 
.A(n_1575),
.B(n_1179),
.C(n_1167),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1485),
.B(n_1053),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1636),
.A2(n_1617),
.B(n_1543),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1542),
.A2(n_1029),
.B(n_1028),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1458),
.B(n_1055),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1484),
.B(n_1488),
.Y(n_1723)
);

INVx4_ASAP7_75t_L g1724 ( 
.A(n_1516),
.Y(n_1724)
);

BUFx8_ASAP7_75t_L g1725 ( 
.A(n_1572),
.Y(n_1725)
);

AO21x1_ASAP7_75t_L g1726 ( 
.A1(n_1588),
.A2(n_1041),
.B(n_1040),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1466),
.B(n_1058),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1553),
.B(n_1470),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1573),
.A2(n_959),
.B1(n_996),
.B2(n_990),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1469),
.B(n_1060),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1471),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1526),
.B(n_1061),
.Y(n_1732)
);

AOI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1512),
.A2(n_1050),
.B(n_1045),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1516),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_R g1735 ( 
.A(n_1528),
.B(n_990),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1631),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1653),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1516),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1585),
.B(n_1490),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1502),
.B(n_1065),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1474),
.A2(n_1059),
.B(n_1057),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1513),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1577),
.A2(n_996),
.B1(n_1037),
.B2(n_1026),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1472),
.Y(n_1744)
);

OAI321xp33_ASAP7_75t_L g1745 ( 
.A1(n_1584),
.A2(n_1068),
.A3(n_1062),
.B1(n_1075),
.B2(n_1070),
.C(n_1064),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1535),
.B(n_1066),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1476),
.A2(n_1083),
.B(n_1082),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1609),
.B(n_1026),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1554),
.B(n_1562),
.Y(n_1749)
);

INVx4_ASAP7_75t_L g1750 ( 
.A(n_1521),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1565),
.B(n_1623),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1521),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1546),
.B(n_1037),
.Y(n_1753)
);

AO21x1_ASAP7_75t_L g1754 ( 
.A1(n_1626),
.A2(n_1089),
.B(n_1087),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1468),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1630),
.A2(n_1477),
.B(n_1625),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1508),
.A2(n_1510),
.B(n_1517),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1524),
.A2(n_1095),
.B(n_1092),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1548),
.B(n_1056),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1552),
.A2(n_1056),
.B1(n_1086),
.B2(n_1072),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1492),
.A2(n_1110),
.B(n_1111),
.C(n_1104),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1523),
.B(n_1072),
.Y(n_1762)
);

AOI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1453),
.A2(n_1116),
.B(n_1115),
.Y(n_1763)
);

NOR3xp33_ASAP7_75t_L g1764 ( 
.A(n_1505),
.B(n_1030),
.C(n_988),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1527),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1580),
.A2(n_1120),
.B(n_1119),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1481),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1607),
.B(n_1497),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1499),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1521),
.Y(n_1770)
);

INVx4_ASAP7_75t_L g1771 ( 
.A(n_1481),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1611),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1611),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1561),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1560),
.B(n_1067),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1582),
.Y(n_1776)
);

INVx4_ASAP7_75t_L g1777 ( 
.A(n_1475),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1597),
.B(n_1071),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1601),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1594),
.A2(n_1126),
.B(n_1124),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1594),
.A2(n_1132),
.B(n_1127),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1594),
.A2(n_1138),
.B(n_1137),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1603),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1610),
.B(n_1073),
.Y(n_1784)
);

A2O1A1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1595),
.A2(n_1144),
.B(n_1145),
.C(n_1141),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1514),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1644),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1642),
.A2(n_1148),
.B(n_1146),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1570),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1564),
.A2(n_1152),
.B(n_1150),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1615),
.B(n_1079),
.Y(n_1791)
);

A2O1A1Ixp33_ASAP7_75t_L g1792 ( 
.A1(n_1596),
.A2(n_1159),
.B(n_1162),
.C(n_1153),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1520),
.A2(n_1080),
.B1(n_1084),
.B2(n_1081),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1591),
.B(n_1086),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1616),
.B(n_1085),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1599),
.A2(n_1174),
.B(n_1178),
.C(n_1165),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1571),
.A2(n_1078),
.B(n_1076),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1650),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1619),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1576),
.A2(n_1118),
.B(n_1097),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1463),
.B(n_1088),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1579),
.A2(n_1161),
.B(n_1156),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1482),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1593),
.A2(n_1046),
.B(n_1003),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1620),
.A2(n_1094),
.B(n_1091),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1628),
.A2(n_1103),
.B(n_1102),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1507),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1629),
.A2(n_1639),
.B(n_1632),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1529),
.B(n_1105),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1533),
.A2(n_1108),
.B(n_1106),
.Y(n_1810)
);

A2O1A1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1604),
.A2(n_1099),
.B(n_1117),
.C(n_1044),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1621),
.A2(n_1114),
.B(n_1112),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1656),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1534),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1467),
.A2(n_1122),
.B(n_1121),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1487),
.B(n_1109),
.Y(n_1816)
);

NAND2xp33_ASAP7_75t_L g1817 ( 
.A(n_1504),
.B(n_1123),
.Y(n_1817)
);

O2A1O1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1605),
.A2(n_1142),
.B(n_1140),
.C(n_1109),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1622),
.A2(n_1129),
.B(n_1128),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1592),
.B(n_1140),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1637),
.A2(n_1461),
.B1(n_1589),
.B2(n_1583),
.Y(n_1821)
);

AND2x2_ASAP7_75t_SL g1822 ( 
.A(n_1627),
.B(n_23),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1518),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1561),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1634),
.A2(n_1131),
.B(n_1130),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1656),
.Y(n_1826)
);

O2A1O1Ixp5_ASAP7_75t_L g1827 ( 
.A1(n_1551),
.A2(n_1139),
.B(n_1143),
.C(n_1134),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1659),
.A2(n_1149),
.B(n_1151),
.C(n_1147),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1602),
.Y(n_1829)
);

O2A1O1Ixp33_ASAP7_75t_L g1830 ( 
.A1(n_1613),
.A2(n_1155),
.B(n_1158),
.C(n_1154),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1590),
.A2(n_1168),
.B(n_1169),
.C(n_1164),
.Y(n_1831)
);

BUFx4f_ASAP7_75t_L g1832 ( 
.A(n_1602),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_SL g1833 ( 
.A(n_1504),
.B(n_1186),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1659),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1637),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1651),
.B(n_24),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1600),
.Y(n_1837)
);

O2A1O1Ixp5_ASAP7_75t_L g1838 ( 
.A1(n_1511),
.A2(n_28),
.B(n_25),
.C(n_26),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1648),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1451),
.B(n_28),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1452),
.B(n_30),
.Y(n_1841)
);

NOR2xp67_ASAP7_75t_L g1842 ( 
.A(n_1660),
.B(n_31),
.Y(n_1842)
);

INVx11_ASAP7_75t_L g1843 ( 
.A(n_1598),
.Y(n_1843)
);

OAI21xp33_ASAP7_75t_L g1844 ( 
.A1(n_1655),
.A2(n_31),
.B(n_32),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1544),
.B(n_34),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_L g1846 ( 
.A(n_1635),
.B(n_35),
.C(n_36),
.Y(n_1846)
);

INVx3_ASAP7_75t_L g1847 ( 
.A(n_1657),
.Y(n_1847)
);

BUFx12f_ASAP7_75t_L g1848 ( 
.A(n_1598),
.Y(n_1848)
);

OAI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1555),
.A2(n_1569),
.B(n_1567),
.Y(n_1849)
);

OAI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1652),
.A2(n_39),
.B(n_40),
.Y(n_1850)
);

NOR3xp33_ASAP7_75t_L g1851 ( 
.A(n_1647),
.B(n_1649),
.C(n_1640),
.Y(n_1851)
);

BUFx2_ASAP7_75t_SL g1852 ( 
.A(n_1657),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1606),
.B(n_41),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1658),
.A2(n_42),
.B(n_43),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1641),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1654),
.A2(n_46),
.B(n_48),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1641),
.B(n_48),
.Y(n_1857)
);

INVxp33_ASAP7_75t_SL g1858 ( 
.A(n_1641),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1614),
.B(n_49),
.Y(n_1859)
);

O2A1O1Ixp33_ASAP7_75t_L g1860 ( 
.A1(n_1454),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1525),
.Y(n_1861)
);

BUFx12f_ASAP7_75t_L g1862 ( 
.A(n_1559),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1465),
.B(n_53),
.Y(n_1863)
);

O2A1O1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1454),
.A2(n_57),
.B(n_54),
.C(n_56),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1454),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1865)
);

O2A1O1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1454),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1454),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1465),
.B(n_62),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1454),
.B(n_63),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1454),
.B(n_64),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1454),
.B(n_65),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1457),
.B(n_784),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1454),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1465),
.B(n_66),
.Y(n_1874)
);

INVx4_ASAP7_75t_SL g1875 ( 
.A(n_1573),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1454),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1454),
.B(n_67),
.Y(n_1877)
);

A2O1A1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1454),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1878)
);

AO22x1_ASAP7_75t_L g1879 ( 
.A1(n_1528),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_1879)
);

CKINVDCx10_ASAP7_75t_R g1880 ( 
.A(n_1572),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1631),
.Y(n_1881)
);

A2O1A1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1454),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_1882)
);

NOR3xp33_ASAP7_75t_L g1883 ( 
.A(n_1568),
.B(n_76),
.C(n_78),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1454),
.A2(n_78),
.B(n_79),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1454),
.B(n_79),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1631),
.Y(n_1886)
);

OAI21xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1454),
.A2(n_80),
.B(n_81),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1454),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1454),
.Y(n_1889)
);

AO21x1_ASAP7_75t_L g1890 ( 
.A1(n_1578),
.A2(n_84),
.B(n_85),
.Y(n_1890)
);

AND2x6_ASAP7_75t_L g1891 ( 
.A(n_1573),
.B(n_84),
.Y(n_1891)
);

AO21x1_ASAP7_75t_L g1892 ( 
.A1(n_1578),
.A2(n_85),
.B(n_86),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1454),
.A2(n_86),
.B(n_87),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1454),
.A2(n_87),
.B(n_89),
.Y(n_1894)
);

AND2x2_ASAP7_75t_SL g1895 ( 
.A(n_1582),
.B(n_89),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1454),
.B(n_90),
.Y(n_1896)
);

AOI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1568),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1897)
);

AND2x6_ASAP7_75t_L g1898 ( 
.A(n_1573),
.B(n_91),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1454),
.B(n_92),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1873),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1876),
.Y(n_1901)
);

BUFx12f_ASAP7_75t_L g1902 ( 
.A(n_1862),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1677),
.B(n_94),
.Y(n_1903)
);

AOI21x1_ASAP7_75t_L g1904 ( 
.A1(n_1763),
.A2(n_1667),
.B(n_1857),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1675),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1889),
.B(n_97),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1813),
.Y(n_1907)
);

AO21x1_ASAP7_75t_L g1908 ( 
.A1(n_1850),
.A2(n_97),
.B(n_98),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1834),
.B(n_100),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1694),
.A2(n_101),
.B(n_102),
.Y(n_1910)
);

NAND2x1p5_ASAP7_75t_L g1911 ( 
.A(n_1724),
.B(n_102),
.Y(n_1911)
);

O2A1O1Ixp5_ASAP7_75t_L g1912 ( 
.A1(n_1840),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1725),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1723),
.B(n_105),
.Y(n_1914)
);

NAND2x1_ASAP7_75t_L g1915 ( 
.A(n_1662),
.B(n_106),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1691),
.B(n_106),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1702),
.B(n_107),
.Y(n_1917)
);

AOI21xp33_ASAP7_75t_L g1918 ( 
.A1(n_1841),
.A2(n_108),
.B(n_109),
.Y(n_1918)
);

AO31x2_ASAP7_75t_L g1919 ( 
.A1(n_1890),
.A2(n_110),
.A3(n_108),
.B(n_109),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1861),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1687),
.A2(n_110),
.B(n_112),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1808),
.A2(n_113),
.B(n_114),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1845),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1757),
.A2(n_116),
.B(n_117),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1686),
.B(n_118),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1683),
.B(n_121),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1670),
.Y(n_1927)
);

AO31x2_ASAP7_75t_L g1928 ( 
.A1(n_1892),
.A2(n_124),
.A3(n_122),
.B(n_123),
.Y(n_1928)
);

AO21x1_ASAP7_75t_L g1929 ( 
.A1(n_1850),
.A2(n_122),
.B(n_125),
.Y(n_1929)
);

NAND2x1p5_ASAP7_75t_L g1930 ( 
.A(n_1724),
.B(n_126),
.Y(n_1930)
);

BUFx12f_ASAP7_75t_L g1931 ( 
.A(n_1725),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1665),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1728),
.A2(n_130),
.B1(n_127),
.B2(n_128),
.C(n_131),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1739),
.B(n_127),
.Y(n_1934)
);

NAND2x1_ASAP7_75t_L g1935 ( 
.A(n_1662),
.B(n_130),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1669),
.B(n_132),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1779),
.B(n_1799),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1720),
.A2(n_134),
.B(n_135),
.Y(n_1938)
);

NAND2x1p5_ASAP7_75t_L g1939 ( 
.A(n_1738),
.B(n_136),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1845),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_1940)
);

NAND3x1_ASAP7_75t_L g1941 ( 
.A(n_1764),
.B(n_143),
.C(n_145),
.Y(n_1941)
);

OAI21x1_ASAP7_75t_L g1942 ( 
.A1(n_1720),
.A2(n_145),
.B(n_146),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1835),
.B(n_148),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1711),
.B(n_148),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1689),
.B(n_149),
.Y(n_1945)
);

OAI21x1_ASAP7_75t_L g1946 ( 
.A1(n_1772),
.A2(n_151),
.B(n_152),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1704),
.A2(n_153),
.B(n_154),
.Y(n_1947)
);

OAI22x1_ASAP7_75t_L g1948 ( 
.A1(n_1816),
.A2(n_1678),
.B1(n_1742),
.B2(n_1771),
.Y(n_1948)
);

AOI21x1_ASAP7_75t_L g1949 ( 
.A1(n_1859),
.A2(n_153),
.B(n_154),
.Y(n_1949)
);

AOI21x1_ASAP7_75t_L g1950 ( 
.A1(n_1773),
.A2(n_155),
.B(n_157),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1735),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1771),
.B(n_158),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1695),
.A2(n_158),
.B(n_159),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1709),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1688),
.Y(n_1955)
);

NAND2xp33_ASAP7_75t_SL g1956 ( 
.A(n_1738),
.B(n_776),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1880),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1768),
.B(n_161),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1737),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1750),
.B(n_165),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1721),
.B(n_1681),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1713),
.Y(n_1962)
);

OAI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1869),
.A2(n_166),
.B(n_167),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1899),
.A2(n_167),
.B(n_168),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1721),
.B(n_168),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1749),
.B(n_169),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1750),
.B(n_169),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1788),
.B(n_170),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1849),
.A2(n_1756),
.B(n_1813),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1748),
.A2(n_175),
.B1(n_172),
.B2(n_173),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1870),
.A2(n_1877),
.B(n_1871),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1733),
.A2(n_176),
.B(n_177),
.Y(n_1972)
);

AND2x4_ASAP7_75t_L g1973 ( 
.A(n_1770),
.B(n_176),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1872),
.B(n_177),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1885),
.A2(n_178),
.B(n_179),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1762),
.B(n_178),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1787),
.B(n_180),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1714),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1676),
.B(n_180),
.Y(n_1979)
);

OAI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1760),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1863),
.B(n_185),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1712),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1783),
.Y(n_1983)
);

BUFx8_ASAP7_75t_SL g1984 ( 
.A(n_1715),
.Y(n_1984)
);

OAI21x1_ASAP7_75t_SL g1985 ( 
.A1(n_1754),
.A2(n_191),
.B(n_192),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_SL g1986 ( 
.A1(n_1729),
.A2(n_193),
.B(n_195),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1753),
.B(n_774),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_SL g1988 ( 
.A1(n_1788),
.A2(n_195),
.B(n_196),
.Y(n_1988)
);

OAI21xp33_ASAP7_75t_L g1989 ( 
.A1(n_1759),
.A2(n_196),
.B(n_198),
.Y(n_1989)
);

AOI21x1_ASAP7_75t_L g1990 ( 
.A1(n_1842),
.A2(n_198),
.B(n_199),
.Y(n_1990)
);

OAI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1896),
.A2(n_1664),
.B(n_1710),
.Y(n_1991)
);

OAI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1790),
.A2(n_202),
.B(n_203),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1868),
.B(n_1874),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1816),
.Y(n_1994)
);

O2A1O1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1811),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_1995)
);

AOI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1826),
.A2(n_204),
.B(n_205),
.Y(n_1996)
);

AOI221x1_ASAP7_75t_L g1997 ( 
.A1(n_1844),
.A2(n_210),
.B1(n_207),
.B2(n_209),
.C(n_211),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1692),
.B(n_207),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1833),
.B(n_211),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1785),
.B(n_213),
.Y(n_2000)
);

NAND2x1p5_ASAP7_75t_L g2001 ( 
.A(n_1770),
.B(n_213),
.Y(n_2001)
);

O2A1O1Ixp33_ASAP7_75t_L g2002 ( 
.A1(n_1761),
.A2(n_1661),
.B(n_1697),
.C(n_1792),
.Y(n_2002)
);

NOR2x1_ASAP7_75t_SL g2003 ( 
.A(n_1852),
.B(n_215),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1826),
.A2(n_214),
.B(n_216),
.Y(n_2004)
);

A2O1A1Ixp33_ASAP7_75t_L g2005 ( 
.A1(n_1741),
.A2(n_217),
.B(n_214),
.C(n_216),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1796),
.B(n_217),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1673),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1708),
.B(n_218),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1747),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1682),
.B(n_220),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1798),
.B(n_221),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_SL g2012 ( 
.A1(n_1895),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_2012)
);

AO21x2_ASAP7_75t_L g2013 ( 
.A1(n_1804),
.A2(n_222),
.B(n_224),
.Y(n_2013)
);

AOI21xp33_ASAP7_75t_L g2014 ( 
.A1(n_1860),
.A2(n_1866),
.B(n_1864),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1822),
.B(n_227),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1821),
.B(n_231),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1832),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1758),
.B(n_233),
.Y(n_2018)
);

OA22x2_ASAP7_75t_L g2019 ( 
.A1(n_1743),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1706),
.B(n_234),
.Y(n_2020)
);

AO31x2_ASAP7_75t_L g2021 ( 
.A1(n_1698),
.A2(n_239),
.A3(n_237),
.B(n_238),
.Y(n_2021)
);

AOI21xp33_ASAP7_75t_L g2022 ( 
.A1(n_1853),
.A2(n_238),
.B(n_241),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1674),
.A2(n_243),
.B(n_244),
.Y(n_2023)
);

INVxp67_ASAP7_75t_SL g2024 ( 
.A(n_1734),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1778),
.A2(n_244),
.B(n_245),
.Y(n_2025)
);

OAI21x1_ASAP7_75t_SL g2026 ( 
.A1(n_1726),
.A2(n_1777),
.B(n_1856),
.Y(n_2026)
);

AOI221x1_ASAP7_75t_L g2027 ( 
.A1(n_1883),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.C(n_248),
.Y(n_2027)
);

BUFx3_ASAP7_75t_L g2028 ( 
.A(n_1832),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1701),
.B(n_246),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1718),
.B(n_247),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1820),
.B(n_248),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1897),
.A2(n_253),
.B1(n_250),
.B2(n_251),
.Y(n_2032)
);

OAI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1797),
.A2(n_253),
.B(n_254),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1803),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1809),
.B(n_257),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1765),
.B(n_257),
.Y(n_2036)
);

OAI21x1_ASAP7_75t_L g2037 ( 
.A1(n_1766),
.A2(n_258),
.B(n_260),
.Y(n_2037)
);

OAI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1800),
.A2(n_261),
.B(n_262),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1784),
.A2(n_263),
.B(n_265),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1836),
.B(n_263),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1802),
.A2(n_266),
.B(n_267),
.Y(n_2041)
);

OAI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1780),
.A2(n_266),
.B(n_268),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_1751),
.B(n_268),
.Y(n_2043)
);

OAI21x1_ASAP7_75t_L g2044 ( 
.A1(n_1781),
.A2(n_269),
.B(n_270),
.Y(n_2044)
);

AND2x4_ASAP7_75t_L g2045 ( 
.A(n_1688),
.B(n_1736),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1782),
.A2(n_269),
.B(n_270),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1769),
.B(n_271),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1671),
.B(n_273),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_1839),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1666),
.B(n_276),
.Y(n_2050)
);

OAI21x1_ASAP7_75t_SL g2051 ( 
.A1(n_1777),
.A2(n_276),
.B(n_277),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1865),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1776),
.B(n_278),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1807),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1716),
.B(n_280),
.Y(n_2055)
);

OAI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1828),
.A2(n_1672),
.B(n_1699),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1703),
.B(n_1679),
.Y(n_2057)
);

NOR2xp67_ASAP7_75t_SL g2058 ( 
.A(n_1774),
.B(n_281),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_L g2059 ( 
.A(n_1786),
.B(n_282),
.C(n_283),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1731),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1848),
.Y(n_2061)
);

NAND2x1_ASAP7_75t_L g2062 ( 
.A(n_1736),
.B(n_284),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1722),
.B(n_286),
.Y(n_2063)
);

NAND2x1p5_ASAP7_75t_L g2064 ( 
.A(n_1881),
.B(n_287),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1823),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1881),
.B(n_289),
.Y(n_2066)
);

OAI21x1_ASAP7_75t_SL g2067 ( 
.A1(n_1884),
.A2(n_289),
.B(n_290),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1727),
.B(n_290),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1887),
.A2(n_291),
.B(n_292),
.Y(n_2069)
);

INVx6_ASAP7_75t_L g2070 ( 
.A(n_1837),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1791),
.A2(n_291),
.B(n_293),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1730),
.B(n_294),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1795),
.A2(n_295),
.B(n_296),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1893),
.A2(n_295),
.B(n_296),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_1829),
.B(n_297),
.Y(n_2075)
);

NAND2xp33_ASAP7_75t_L g2076 ( 
.A(n_1734),
.B(n_298),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1793),
.B(n_299),
.Y(n_2077)
);

OAI22x1_ASAP7_75t_L g2078 ( 
.A1(n_1767),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1707),
.B(n_302),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1732),
.Y(n_2080)
);

BUFx8_ASAP7_75t_SL g2081 ( 
.A(n_1847),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1734),
.Y(n_2082)
);

BUFx8_ASAP7_75t_SL g2083 ( 
.A(n_1847),
.Y(n_2083)
);

AO21x1_ASAP7_75t_L g2084 ( 
.A1(n_1894),
.A2(n_303),
.B(n_304),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1740),
.B(n_304),
.Y(n_2085)
);

OAI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_1805),
.A2(n_1806),
.B(n_1867),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1746),
.B(n_305),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1752),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1719),
.B(n_307),
.Y(n_2089)
);

INVx3_ASAP7_75t_L g2090 ( 
.A(n_1886),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1886),
.B(n_307),
.Y(n_2091)
);

NAND2x1p5_ASAP7_75t_L g2092 ( 
.A(n_1752),
.B(n_308),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1789),
.B(n_1693),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1794),
.B(n_310),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1812),
.B(n_311),
.Y(n_2095)
);

OAI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1855),
.A2(n_1882),
.B1(n_1878),
.B2(n_1858),
.Y(n_2096)
);

A2O1A1Ixp33_ASAP7_75t_L g2097 ( 
.A1(n_1854),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1888),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1752),
.Y(n_2099)
);

NOR2xp67_ASAP7_75t_L g2100 ( 
.A(n_1824),
.B(n_317),
.Y(n_2100)
);

INVx8_ASAP7_75t_L g2101 ( 
.A(n_1891),
.Y(n_2101)
);

AOI21xp5_ASAP7_75t_L g2102 ( 
.A1(n_1801),
.A2(n_318),
.B(n_320),
.Y(n_2102)
);

OAI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_1700),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_2103)
);

NAND2x1p5_ASAP7_75t_L g2104 ( 
.A(n_1717),
.B(n_324),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1680),
.Y(n_2105)
);

INVx3_ASAP7_75t_L g2106 ( 
.A(n_1814),
.Y(n_2106)
);

INVx1_ASAP7_75t_SL g2107 ( 
.A(n_1891),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1745),
.B(n_1685),
.Y(n_2108)
);

OAI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_1831),
.A2(n_325),
.B(n_326),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1690),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1819),
.B(n_327),
.Y(n_2111)
);

NOR2xp67_ASAP7_75t_L g2112 ( 
.A(n_1696),
.B(n_329),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_1817),
.A2(n_1705),
.B(n_1825),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1818),
.B(n_332),
.Y(n_2114)
);

OAI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_1838),
.A2(n_333),
.B(n_334),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1891),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_1875),
.B(n_336),
.Y(n_2117)
);

NAND2x1_ASAP7_75t_L g2118 ( 
.A(n_1891),
.B(n_337),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1875),
.B(n_340),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_1775),
.A2(n_341),
.B(n_342),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_1810),
.A2(n_1815),
.B(n_1684),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1663),
.A2(n_345),
.B1(n_341),
.B2(n_344),
.Y(n_2122)
);

AOI221xp5_ASAP7_75t_L g2123 ( 
.A1(n_1685),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.C(n_349),
.Y(n_2123)
);

OR2x6_ASAP7_75t_L g2124 ( 
.A(n_1879),
.B(n_346),
.Y(n_2124)
);

NOR2x1_ASAP7_75t_L g2125 ( 
.A(n_1668),
.B(n_347),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_SL g2126 ( 
.A(n_1898),
.B(n_348),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1744),
.B(n_349),
.Y(n_2127)
);

O2A1O1Ixp5_ASAP7_75t_L g2128 ( 
.A1(n_1827),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1898),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1898),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1830),
.B(n_353),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_1843),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1755),
.B(n_1898),
.Y(n_2133)
);

OAI21xp33_ASAP7_75t_SL g2134 ( 
.A1(n_1875),
.A2(n_355),
.B(n_356),
.Y(n_2134)
);

AO31x2_ASAP7_75t_L g2135 ( 
.A1(n_1846),
.A2(n_358),
.A3(n_356),
.B(n_357),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_1851),
.A2(n_359),
.B(n_361),
.Y(n_2136)
);

NAND2xp33_ASAP7_75t_L g2137 ( 
.A(n_1813),
.B(n_359),
.Y(n_2137)
);

AOI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_1667),
.A2(n_361),
.B(n_362),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1873),
.B(n_362),
.Y(n_2139)
);

NOR2x1_ASAP7_75t_SL g2140 ( 
.A(n_1873),
.B(n_363),
.Y(n_2140)
);

NAND2x1_ASAP7_75t_L g2141 ( 
.A(n_1873),
.B(n_363),
.Y(n_2141)
);

NAND3xp33_ASAP7_75t_L g2142 ( 
.A(n_1749),
.B(n_364),
.C(n_365),
.Y(n_2142)
);

AOI21x1_ASAP7_75t_SL g2143 ( 
.A1(n_1711),
.A2(n_364),
.B(n_366),
.Y(n_2143)
);

OAI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_1667),
.A2(n_366),
.B(n_367),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1667),
.A2(n_367),
.B(n_368),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_1873),
.B(n_370),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1873),
.B(n_370),
.Y(n_2147)
);

OAI21xp5_ASAP7_75t_L g2148 ( 
.A1(n_1667),
.A2(n_371),
.B(n_372),
.Y(n_2148)
);

OAI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_1667),
.A2(n_371),
.B(n_372),
.Y(n_2149)
);

OA21x2_ASAP7_75t_L g2150 ( 
.A1(n_1667),
.A2(n_373),
.B(n_374),
.Y(n_2150)
);

AOI21xp5_ASAP7_75t_L g2151 ( 
.A1(n_1667),
.A2(n_373),
.B(n_374),
.Y(n_2151)
);

O2A1O1Ixp33_ASAP7_75t_L g2152 ( 
.A1(n_1811),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_2152)
);

A2O1A1Ixp33_ASAP7_75t_L g2153 ( 
.A1(n_1702),
.A2(n_381),
.B(n_377),
.C(n_380),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_1873),
.Y(n_2154)
);

AOI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_1667),
.A2(n_380),
.B(n_381),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_1873),
.B(n_382),
.Y(n_2156)
);

OAI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_1667),
.A2(n_383),
.B(n_384),
.Y(n_2157)
);

INVx4_ASAP7_75t_L g2158 ( 
.A(n_1832),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1873),
.B(n_385),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_1873),
.B(n_386),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_1873),
.B(n_388),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_1677),
.B(n_390),
.Y(n_2162)
);

AOI21xp5_ASAP7_75t_L g2163 ( 
.A1(n_1667),
.A2(n_390),
.B(n_392),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1873),
.B(n_393),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1873),
.B(n_393),
.Y(n_2165)
);

O2A1O1Ixp33_ASAP7_75t_L g2166 ( 
.A1(n_1811),
.A2(n_396),
.B(n_394),
.C(n_395),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1873),
.B(n_395),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_SL g2168 ( 
.A1(n_1845),
.A2(n_396),
.B(n_397),
.Y(n_2168)
);

OAI22x1_ASAP7_75t_L g2169 ( 
.A1(n_1816),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_2169)
);

BUFx12f_ASAP7_75t_L g2170 ( 
.A(n_1862),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_1662),
.Y(n_2171)
);

OAI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_1667),
.A2(n_398),
.B(n_399),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_1667),
.A2(n_400),
.B(n_403),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_1677),
.B(n_405),
.Y(n_2174)
);

OAI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_1667),
.A2(n_407),
.B(n_408),
.Y(n_2175)
);

AO21x2_ASAP7_75t_L g2176 ( 
.A1(n_1667),
.A2(n_410),
.B(n_411),
.Y(n_2176)
);

INVx5_ASAP7_75t_L g2177 ( 
.A(n_1891),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1873),
.B(n_411),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_1667),
.A2(n_413),
.B(n_414),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1873),
.B(n_414),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_1678),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1873),
.B(n_417),
.Y(n_2182)
);

BUFx12f_ASAP7_75t_L g2183 ( 
.A(n_1862),
.Y(n_2183)
);

OAI21x1_ASAP7_75t_SL g2184 ( 
.A1(n_1850),
.A2(n_418),
.B(n_419),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_1667),
.A2(n_420),
.B(n_421),
.Y(n_2185)
);

NOR2x1_ASAP7_75t_SL g2186 ( 
.A(n_1873),
.B(n_420),
.Y(n_2186)
);

A2O1A1Ixp33_ASAP7_75t_L g2187 ( 
.A1(n_1702),
.A2(n_424),
.B(n_422),
.C(n_423),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1873),
.B(n_423),
.Y(n_2188)
);

A2O1A1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_1702),
.A2(n_427),
.B(n_425),
.C(n_426),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_1662),
.Y(n_2190)
);

INVx3_ASAP7_75t_SL g2191 ( 
.A(n_1774),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1873),
.B(n_429),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1873),
.B(n_430),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1873),
.B(n_431),
.Y(n_2194)
);

OA22x2_ASAP7_75t_L g2195 ( 
.A1(n_1729),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_SL g2196 ( 
.A1(n_1850),
.A2(n_434),
.B(n_435),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1873),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1873),
.B(n_435),
.Y(n_2198)
);

OAI21x1_ASAP7_75t_SL g2199 ( 
.A1(n_1850),
.A2(n_436),
.B(n_438),
.Y(n_2199)
);

A2O1A1Ixp33_ASAP7_75t_L g2200 ( 
.A1(n_1702),
.A2(n_439),
.B(n_436),
.C(n_438),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_1873),
.A2(n_443),
.B1(n_440),
.B2(n_442),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1873),
.Y(n_2202)
);

AO21x1_ASAP7_75t_L g2203 ( 
.A1(n_1850),
.A2(n_440),
.B(n_443),
.Y(n_2203)
);

OAI21xp33_ASAP7_75t_L g2204 ( 
.A1(n_1728),
.A2(n_444),
.B(n_445),
.Y(n_2204)
);

AOI21xp5_ASAP7_75t_L g2205 ( 
.A1(n_1667),
.A2(n_445),
.B(n_446),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1873),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1873),
.B(n_446),
.Y(n_2207)
);

OAI21xp33_ASAP7_75t_L g2208 ( 
.A1(n_1728),
.A2(n_447),
.B(n_448),
.Y(n_2208)
);

AOI21xp33_ASAP7_75t_L g2209 ( 
.A1(n_1840),
.A2(n_448),
.B(n_450),
.Y(n_2209)
);

BUFx6f_ASAP7_75t_L g2210 ( 
.A(n_1813),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1873),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_1677),
.B(n_450),
.Y(n_2212)
);

AOI21xp33_ASAP7_75t_L g2213 ( 
.A1(n_1840),
.A2(n_451),
.B(n_453),
.Y(n_2213)
);

NAND2xp33_ASAP7_75t_L g2214 ( 
.A(n_1813),
.B(n_451),
.Y(n_2214)
);

NOR2x1_ASAP7_75t_SL g2215 ( 
.A(n_1873),
.B(n_453),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1873),
.B(n_454),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_1725),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_SL g2218 ( 
.A(n_1724),
.B(n_455),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_1677),
.B(n_456),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_1667),
.A2(n_459),
.B(n_460),
.Y(n_2220)
);

OAI22x1_ASAP7_75t_L g2221 ( 
.A1(n_1816),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_2221)
);

AOI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_1667),
.A2(n_461),
.B(n_462),
.Y(n_2222)
);

AO31x2_ASAP7_75t_L g2223 ( 
.A1(n_1890),
.A2(n_465),
.A3(n_463),
.B(n_464),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1873),
.B(n_463),
.Y(n_2224)
);

INVx1_ASAP7_75t_SL g2225 ( 
.A(n_1873),
.Y(n_2225)
);

OAI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_1667),
.A2(n_465),
.B(n_466),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1873),
.B(n_467),
.Y(n_2227)
);

NAND2x1_ASAP7_75t_L g2228 ( 
.A(n_1873),
.B(n_468),
.Y(n_2228)
);

NAND2x1_ASAP7_75t_L g2229 ( 
.A(n_1873),
.B(n_469),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1873),
.B(n_471),
.Y(n_2230)
);

OA22x2_ASAP7_75t_L g2231 ( 
.A1(n_1729),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_1873),
.B(n_472),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1873),
.B(n_475),
.Y(n_2233)
);

INVx2_ASAP7_75t_SL g2234 ( 
.A(n_1832),
.Y(n_2234)
);

AOI21xp5_ASAP7_75t_L g2235 ( 
.A1(n_1667),
.A2(n_476),
.B(n_477),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1873),
.B(n_479),
.Y(n_2236)
);

INVx2_ASAP7_75t_SL g2237 ( 
.A(n_1832),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1873),
.B(n_479),
.Y(n_2238)
);

BUFx3_ASAP7_75t_L g2239 ( 
.A(n_1725),
.Y(n_2239)
);

OAI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_1667),
.A2(n_480),
.B(n_481),
.Y(n_2240)
);

CKINVDCx6p67_ASAP7_75t_R g2241 ( 
.A(n_1862),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1813),
.Y(n_2242)
);

AOI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_1667),
.A2(n_480),
.B(n_482),
.Y(n_2243)
);

AOI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_1667),
.A2(n_482),
.B(n_483),
.Y(n_2244)
);

OAI22x1_ASAP7_75t_L g2245 ( 
.A1(n_1816),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_1832),
.Y(n_2246)
);

AOI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_1835),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1873),
.B(n_491),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1873),
.B(n_492),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_1667),
.A2(n_492),
.B(n_493),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_1662),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1873),
.Y(n_2252)
);

AOI21xp33_ASAP7_75t_L g2253 ( 
.A1(n_1840),
.A2(n_494),
.B(n_495),
.Y(n_2253)
);

INVxp67_ASAP7_75t_SL g2254 ( 
.A(n_1873),
.Y(n_2254)
);

NAND2x1p5_ASAP7_75t_L g2255 ( 
.A(n_1724),
.B(n_497),
.Y(n_2255)
);

OAI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_1873),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_2256)
);

NAND2x1p5_ASAP7_75t_L g2257 ( 
.A(n_1724),
.B(n_498),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1873),
.Y(n_2258)
);

AOI21xp5_ASAP7_75t_L g2259 ( 
.A1(n_1667),
.A2(n_499),
.B(n_500),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_L g2260 ( 
.A(n_1748),
.B(n_501),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1873),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1873),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_1862),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_1667),
.A2(n_505),
.B(n_506),
.Y(n_2264)
);

A2O1A1Ixp33_ASAP7_75t_L g2265 ( 
.A1(n_1702),
.A2(n_508),
.B(n_506),
.C(n_507),
.Y(n_2265)
);

INVx6_ASAP7_75t_SL g2266 ( 
.A(n_1816),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_1748),
.B(n_509),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_1873),
.B(n_511),
.Y(n_2268)
);

A2O1A1Ixp33_ASAP7_75t_L g2269 ( 
.A1(n_1702),
.A2(n_515),
.B(n_511),
.C(n_513),
.Y(n_2269)
);

NOR2x1_ASAP7_75t_SL g2270 ( 
.A(n_1873),
.B(n_517),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1873),
.B(n_518),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_1873),
.B(n_518),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1873),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1873),
.Y(n_2274)
);

AO31x2_ASAP7_75t_L g2275 ( 
.A1(n_1890),
.A2(n_524),
.A3(n_522),
.B(n_523),
.Y(n_2275)
);

AOI21xp5_ASAP7_75t_L g2276 ( 
.A1(n_1667),
.A2(n_526),
.B(n_527),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_1832),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1873),
.B(n_528),
.Y(n_2278)
);

AOI21xp5_ASAP7_75t_L g2279 ( 
.A1(n_1667),
.A2(n_528),
.B(n_529),
.Y(n_2279)
);

OAI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_1873),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_1667),
.A2(n_531),
.B(n_532),
.Y(n_2281)
);

OAI22x1_ASAP7_75t_L g2282 ( 
.A1(n_1816),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_1873),
.B(n_535),
.Y(n_2283)
);

OAI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_1667),
.A2(n_536),
.B(n_538),
.Y(n_2284)
);

NAND3xp33_ASAP7_75t_L g2285 ( 
.A(n_2027),
.B(n_538),
.C(n_539),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_1901),
.Y(n_2286)
);

INVx2_ASAP7_75t_SL g2287 ( 
.A(n_1931),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1900),
.Y(n_2288)
);

NOR2xp33_ASAP7_75t_L g2289 ( 
.A(n_1901),
.B(n_540),
.Y(n_2289)
);

OA21x2_ASAP7_75t_L g2290 ( 
.A1(n_1942),
.A2(n_540),
.B(n_541),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2202),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2154),
.B(n_2225),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_1971),
.A2(n_1969),
.B(n_1991),
.Y(n_2293)
);

INVx2_ASAP7_75t_SL g2294 ( 
.A(n_1913),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2211),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2154),
.B(n_2225),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_1984),
.Y(n_2297)
);

AO21x2_ASAP7_75t_L g2298 ( 
.A1(n_1904),
.A2(n_542),
.B(n_544),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2254),
.B(n_542),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_1937),
.B(n_546),
.Y(n_2300)
);

OAI21x1_ASAP7_75t_L g2301 ( 
.A1(n_2143),
.A2(n_547),
.B(n_549),
.Y(n_2301)
);

CKINVDCx6p67_ASAP7_75t_R g2302 ( 
.A(n_2241),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2197),
.Y(n_2303)
);

HB1xp67_ASAP7_75t_L g2304 ( 
.A(n_2146),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_2126),
.B(n_547),
.Y(n_2305)
);

AOI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_2098),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_2306)
);

INVx1_ASAP7_75t_SL g2307 ( 
.A(n_2049),
.Y(n_2307)
);

AO21x2_ASAP7_75t_L g2308 ( 
.A1(n_2014),
.A2(n_552),
.B(n_553),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_1937),
.B(n_786),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2252),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2049),
.A2(n_557),
.B1(n_554),
.B2(n_555),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_1902),
.Y(n_2312)
);

NAND2x1p5_ASAP7_75t_L g2313 ( 
.A(n_2177),
.B(n_557),
.Y(n_2313)
);

OAI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_1961),
.A2(n_558),
.B(n_559),
.Y(n_2314)
);

OAI21x1_ASAP7_75t_L g2315 ( 
.A1(n_1917),
.A2(n_560),
.B(n_561),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_L g2316 ( 
.A1(n_2124),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2206),
.Y(n_2317)
);

CKINVDCx20_ASAP7_75t_R g2318 ( 
.A(n_1905),
.Y(n_2318)
);

BUFx3_ASAP7_75t_L g2319 ( 
.A(n_2082),
.Y(n_2319)
);

AOI21x1_ASAP7_75t_L g2320 ( 
.A1(n_2129),
.A2(n_563),
.B(n_564),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2261),
.Y(n_2321)
);

NAND2x1p5_ASAP7_75t_L g2322 ( 
.A(n_2177),
.B(n_563),
.Y(n_2322)
);

OAI21xp5_ASAP7_75t_L g2323 ( 
.A1(n_1961),
.A2(n_1993),
.B(n_2014),
.Y(n_2323)
);

AO21x2_ASAP7_75t_L g2324 ( 
.A1(n_2184),
.A2(n_564),
.B(n_565),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2273),
.Y(n_2325)
);

OR2x6_ASAP7_75t_L g2326 ( 
.A(n_2101),
.B(n_2158),
.Y(n_2326)
);

INVx4_ASAP7_75t_L g2327 ( 
.A(n_2170),
.Y(n_2327)
);

CKINVDCx6p67_ASAP7_75t_R g2328 ( 
.A(n_2183),
.Y(n_2328)
);

INVx4_ASAP7_75t_L g2329 ( 
.A(n_2217),
.Y(n_2329)
);

AO31x2_ASAP7_75t_L g2330 ( 
.A1(n_1908),
.A2(n_568),
.A3(n_566),
.B(n_567),
.Y(n_2330)
);

BUFx2_ASAP7_75t_L g2331 ( 
.A(n_1927),
.Y(n_2331)
);

INVx3_ASAP7_75t_L g2332 ( 
.A(n_2101),
.Y(n_2332)
);

BUFx3_ASAP7_75t_L g2333 ( 
.A(n_2082),
.Y(n_2333)
);

INVx3_ASAP7_75t_L g2334 ( 
.A(n_2101),
.Y(n_2334)
);

BUFx2_ASAP7_75t_SL g2335 ( 
.A(n_2239),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2258),
.Y(n_2336)
);

OAI21xp5_ASAP7_75t_SL g2337 ( 
.A1(n_2012),
.A2(n_1986),
.B(n_2015),
.Y(n_2337)
);

AOI21x1_ASAP7_75t_L g2338 ( 
.A1(n_2130),
.A2(n_571),
.B(n_572),
.Y(n_2338)
);

OR2x2_ASAP7_75t_L g2339 ( 
.A(n_2262),
.B(n_573),
.Y(n_2339)
);

OA21x2_ASAP7_75t_L g2340 ( 
.A1(n_1997),
.A2(n_574),
.B(n_575),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2274),
.B(n_576),
.Y(n_2341)
);

OAI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_1958),
.A2(n_577),
.B(n_578),
.Y(n_2342)
);

NAND2x1p5_ASAP7_75t_L g2343 ( 
.A(n_2177),
.B(n_582),
.Y(n_2343)
);

OA21x2_ASAP7_75t_L g2344 ( 
.A1(n_1938),
.A2(n_582),
.B(n_583),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1959),
.B(n_583),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1907),
.Y(n_2346)
);

BUFx12f_ASAP7_75t_L g2347 ( 
.A(n_2263),
.Y(n_2347)
);

INVx4_ASAP7_75t_L g2348 ( 
.A(n_2158),
.Y(n_2348)
);

INVx3_ASAP7_75t_L g2349 ( 
.A(n_2082),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1906),
.Y(n_2350)
);

HB1xp67_ASAP7_75t_L g2351 ( 
.A(n_2146),
.Y(n_2351)
);

OAI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_1958),
.A2(n_589),
.B(n_591),
.Y(n_2352)
);

BUFx3_ASAP7_75t_L g2353 ( 
.A(n_2088),
.Y(n_2353)
);

AO21x2_ASAP7_75t_L g2354 ( 
.A1(n_2196),
.A2(n_591),
.B(n_592),
.Y(n_2354)
);

AO21x2_ASAP7_75t_L g2355 ( 
.A1(n_2199),
.A2(n_592),
.B(n_593),
.Y(n_2355)
);

OA21x2_ASAP7_75t_L g2356 ( 
.A1(n_1938),
.A2(n_594),
.B(n_595),
.Y(n_2356)
);

AO21x2_ASAP7_75t_L g2357 ( 
.A1(n_1910),
.A2(n_598),
.B(n_599),
.Y(n_2357)
);

OAI21x1_ASAP7_75t_SL g2358 ( 
.A1(n_1910),
.A2(n_599),
.B(n_600),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1906),
.Y(n_2359)
);

BUFx3_ASAP7_75t_L g2360 ( 
.A(n_2088),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_1957),
.Y(n_2361)
);

AND2x4_ASAP7_75t_L g2362 ( 
.A(n_2080),
.B(n_784),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_2088),
.Y(n_2363)
);

OA21x2_ASAP7_75t_L g2364 ( 
.A1(n_1971),
.A2(n_600),
.B(n_601),
.Y(n_2364)
);

AO21x2_ASAP7_75t_L g2365 ( 
.A1(n_2144),
.A2(n_604),
.B(n_605),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2159),
.Y(n_2366)
);

OAI21xp33_ASAP7_75t_SL g2367 ( 
.A1(n_2107),
.A2(n_606),
.B(n_607),
.Y(n_2367)
);

BUFx3_ASAP7_75t_L g2368 ( 
.A(n_2099),
.Y(n_2368)
);

AOI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_1991),
.A2(n_2086),
.B(n_2113),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2159),
.Y(n_2370)
);

AO31x2_ASAP7_75t_L g2371 ( 
.A1(n_1929),
.A2(n_606),
.A3(n_607),
.B(n_608),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2178),
.Y(n_2372)
);

AO31x2_ASAP7_75t_L g2373 ( 
.A1(n_2203),
.A2(n_608),
.A3(n_609),
.B(n_610),
.Y(n_2373)
);

INVx3_ASAP7_75t_L g2374 ( 
.A(n_2099),
.Y(n_2374)
);

BUFx2_ASAP7_75t_R g2375 ( 
.A(n_2061),
.Y(n_2375)
);

NOR2xp33_ASAP7_75t_L g2376 ( 
.A(n_1994),
.B(n_612),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_2191),
.Y(n_2377)
);

AOI21x1_ASAP7_75t_L g2378 ( 
.A1(n_1949),
.A2(n_614),
.B(n_615),
.Y(n_2378)
);

BUFx2_ASAP7_75t_SL g2379 ( 
.A(n_2028),
.Y(n_2379)
);

INVx4_ASAP7_75t_L g2380 ( 
.A(n_2132),
.Y(n_2380)
);

BUFx12f_ASAP7_75t_L g2381 ( 
.A(n_2017),
.Y(n_2381)
);

AO21x2_ASAP7_75t_L g2382 ( 
.A1(n_2148),
.A2(n_616),
.B(n_617),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2178),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2002),
.B(n_616),
.Y(n_2384)
);

NAND2x1p5_ASAP7_75t_L g2385 ( 
.A(n_2116),
.B(n_617),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2182),
.Y(n_2386)
);

OA21x2_ASAP7_75t_L g2387 ( 
.A1(n_2148),
.A2(n_618),
.B(n_619),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_1983),
.B(n_620),
.Y(n_2388)
);

AO21x2_ASAP7_75t_L g2389 ( 
.A1(n_2149),
.A2(n_621),
.B(n_622),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2182),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2093),
.B(n_621),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_1926),
.B(n_622),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2188),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2188),
.Y(n_2394)
);

BUFx2_ASAP7_75t_SL g2395 ( 
.A(n_2234),
.Y(n_2395)
);

OAI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_1966),
.A2(n_624),
.B(n_625),
.Y(n_2396)
);

CKINVDCx6p67_ASAP7_75t_R g2397 ( 
.A(n_1951),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_1944),
.A2(n_626),
.B(n_627),
.Y(n_2398)
);

OA21x2_ASAP7_75t_L g2399 ( 
.A1(n_2149),
.A2(n_626),
.B(n_627),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_R g2400 ( 
.A(n_2116),
.B(n_629),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2192),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_2099),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_1944),
.A2(n_630),
.B(n_631),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2210),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_2210),
.Y(n_2405)
);

OA21x2_ASAP7_75t_L g2406 ( 
.A1(n_2157),
.A2(n_634),
.B(n_635),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2192),
.Y(n_2407)
);

AOI221xp5_ASAP7_75t_L g2408 ( 
.A1(n_1948),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.C(n_637),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2194),
.Y(n_2409)
);

OAI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_1966),
.A2(n_638),
.B(n_639),
.Y(n_2410)
);

BUFx2_ASAP7_75t_R g2411 ( 
.A(n_2081),
.Y(n_2411)
);

NAND2x1p5_ASAP7_75t_L g2412 ( 
.A(n_2116),
.B(n_1960),
.Y(n_2412)
);

AO21x2_ASAP7_75t_L g2413 ( 
.A1(n_2157),
.A2(n_641),
.B(n_642),
.Y(n_2413)
);

OAI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2096),
.A2(n_641),
.B(n_642),
.Y(n_2414)
);

BUFx8_ASAP7_75t_L g2415 ( 
.A(n_2237),
.Y(n_2415)
);

OA21x2_ASAP7_75t_L g2416 ( 
.A1(n_2172),
.A2(n_643),
.B(n_644),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2194),
.Y(n_2417)
);

NAND3xp33_ASAP7_75t_L g2418 ( 
.A(n_1987),
.B(n_644),
.C(n_645),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_1943),
.B(n_646),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_1936),
.B(n_648),
.Y(n_2420)
);

INVx1_ASAP7_75t_SL g2421 ( 
.A(n_1932),
.Y(n_2421)
);

BUFx2_ASAP7_75t_L g2422 ( 
.A(n_2266),
.Y(n_2422)
);

OA21x2_ASAP7_75t_L g2423 ( 
.A1(n_2172),
.A2(n_648),
.B(n_649),
.Y(n_2423)
);

NOR2xp67_ASAP7_75t_L g2424 ( 
.A(n_2246),
.B(n_650),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2198),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2198),
.Y(n_2426)
);

AO21x2_ASAP7_75t_L g2427 ( 
.A1(n_2175),
.A2(n_650),
.B(n_651),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2207),
.Y(n_2428)
);

NOR2x1_ASAP7_75t_R g2429 ( 
.A(n_2117),
.B(n_651),
.Y(n_2429)
);

OR2x2_ASAP7_75t_L g2430 ( 
.A(n_1903),
.B(n_652),
.Y(n_2430)
);

AO21x2_ASAP7_75t_L g2431 ( 
.A1(n_2175),
.A2(n_655),
.B(n_657),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2207),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2216),
.Y(n_2433)
);

AO222x2_ASAP7_75t_L g2434 ( 
.A1(n_2030),
.A2(n_655),
.B1(n_658),
.B2(n_659),
.C1(n_660),
.C2(n_661),
.Y(n_2434)
);

CKINVDCx20_ASAP7_75t_R g2435 ( 
.A(n_2083),
.Y(n_2435)
);

OAI21x1_ASAP7_75t_SL g2436 ( 
.A1(n_2284),
.A2(n_658),
.B(n_659),
.Y(n_2436)
);

OAI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2096),
.A2(n_660),
.B(n_662),
.Y(n_2437)
);

AO31x2_ASAP7_75t_L g2438 ( 
.A1(n_2084),
.A2(n_662),
.A3(n_663),
.B(n_664),
.Y(n_2438)
);

OAI21x1_ASAP7_75t_SL g2439 ( 
.A1(n_2179),
.A2(n_665),
.B(n_666),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2216),
.Y(n_2440)
);

NAND2x1p5_ASAP7_75t_L g2441 ( 
.A(n_1960),
.B(n_667),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_2162),
.B(n_2174),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2156),
.A2(n_668),
.B1(n_669),
.B2(n_670),
.Y(n_2443)
);

OAI21x1_ASAP7_75t_SL g2444 ( 
.A1(n_2284),
.A2(n_669),
.B(n_671),
.Y(n_2444)
);

OAI21x1_ASAP7_75t_L g2445 ( 
.A1(n_2026),
.A2(n_671),
.B(n_672),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2283),
.A2(n_673),
.B1(n_674),
.B2(n_675),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2045),
.Y(n_2447)
);

AO21x2_ASAP7_75t_L g2448 ( 
.A1(n_2179),
.A2(n_674),
.B(n_675),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2224),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2224),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_1934),
.B(n_676),
.Y(n_2451)
);

AO21x2_ASAP7_75t_L g2452 ( 
.A1(n_2226),
.A2(n_677),
.B(n_679),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2248),
.Y(n_2453)
);

AO21x2_ASAP7_75t_L g2454 ( 
.A1(n_2226),
.A2(n_680),
.B(n_681),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2248),
.Y(n_2455)
);

NAND2x1p5_ASAP7_75t_L g2456 ( 
.A(n_1967),
.B(n_683),
.Y(n_2456)
);

OR2x2_ASAP7_75t_L g2457 ( 
.A(n_2212),
.B(n_684),
.Y(n_2457)
);

INVx2_ASAP7_75t_SL g2458 ( 
.A(n_2070),
.Y(n_2458)
);

AO21x2_ASAP7_75t_L g2459 ( 
.A1(n_2240),
.A2(n_687),
.B(n_688),
.Y(n_2459)
);

HB1xp67_ASAP7_75t_L g2460 ( 
.A(n_2156),
.Y(n_2460)
);

HB1xp67_ASAP7_75t_L g2461 ( 
.A(n_2164),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2249),
.Y(n_2462)
);

BUFx12f_ASAP7_75t_L g2463 ( 
.A(n_2277),
.Y(n_2463)
);

OAI21x1_ASAP7_75t_L g2464 ( 
.A1(n_1990),
.A2(n_689),
.B(n_691),
.Y(n_2464)
);

OAI21x1_ASAP7_75t_L g2465 ( 
.A1(n_1946),
.A2(n_693),
.B(n_694),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2249),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2278),
.Y(n_2467)
);

BUFx3_ASAP7_75t_L g2468 ( 
.A(n_2070),
.Y(n_2468)
);

OAI21x1_ASAP7_75t_SL g2469 ( 
.A1(n_2240),
.A2(n_695),
.B(n_696),
.Y(n_2469)
);

OAI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_1914),
.A2(n_696),
.B(n_697),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_2266),
.Y(n_2471)
);

INVx3_ASAP7_75t_L g2472 ( 
.A(n_2045),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_1976),
.B(n_697),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2219),
.B(n_699),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2242),
.Y(n_2475)
);

INVx3_ASAP7_75t_L g2476 ( 
.A(n_2117),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_1943),
.B(n_700),
.Y(n_2477)
);

BUFx2_ASAP7_75t_SL g2478 ( 
.A(n_2119),
.Y(n_2478)
);

CKINVDCx6p67_ASAP7_75t_R g2479 ( 
.A(n_2124),
.Y(n_2479)
);

OA21x2_ASAP7_75t_L g2480 ( 
.A1(n_2250),
.A2(n_701),
.B(n_702),
.Y(n_2480)
);

A2O1A1Ixp33_ASAP7_75t_L g2481 ( 
.A1(n_2069),
.A2(n_701),
.B(n_702),
.C(n_704),
.Y(n_2481)
);

OAI21xp5_ASAP7_75t_L g2482 ( 
.A1(n_1914),
.A2(n_705),
.B(n_706),
.Y(n_2482)
);

BUFx12f_ASAP7_75t_L g2483 ( 
.A(n_1952),
.Y(n_2483)
);

INVxp67_ASAP7_75t_L g2484 ( 
.A(n_2218),
.Y(n_2484)
);

BUFx2_ASAP7_75t_L g2485 ( 
.A(n_1967),
.Y(n_2485)
);

OAI21x1_ASAP7_75t_L g2486 ( 
.A1(n_2250),
.A2(n_707),
.B(n_708),
.Y(n_2486)
);

OAI21xp5_ASAP7_75t_L g2487 ( 
.A1(n_2016),
.A2(n_709),
.B(n_711),
.Y(n_2487)
);

NOR2xp67_ASAP7_75t_SL g2488 ( 
.A(n_2168),
.B(n_712),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_1945),
.B(n_713),
.Y(n_2489)
);

OAI21x1_ASAP7_75t_L g2490 ( 
.A1(n_2136),
.A2(n_716),
.B(n_717),
.Y(n_2490)
);

BUFx6f_ASAP7_75t_L g2491 ( 
.A(n_2118),
.Y(n_2491)
);

OA21x2_ASAP7_75t_L g2492 ( 
.A1(n_2115),
.A2(n_717),
.B(n_718),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2164),
.B(n_718),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_1909),
.B(n_2007),
.Y(n_2494)
);

BUFx2_ASAP7_75t_L g2495 ( 
.A(n_1973),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2056),
.B(n_719),
.Y(n_2496)
);

CKINVDCx20_ASAP7_75t_R g2497 ( 
.A(n_1956),
.Y(n_2497)
);

NAND2x1p5_ASAP7_75t_L g2498 ( 
.A(n_1973),
.B(n_720),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_1955),
.Y(n_2499)
);

NAND2x1p5_ASAP7_75t_L g2500 ( 
.A(n_2283),
.B(n_2119),
.Y(n_2500)
);

NAND2x1p5_ASAP7_75t_L g2501 ( 
.A(n_2107),
.B(n_721),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_1979),
.B(n_722),
.Y(n_2502)
);

OAI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2016),
.A2(n_723),
.B(n_725),
.Y(n_2503)
);

OAI21x1_ASAP7_75t_L g2504 ( 
.A1(n_2150),
.A2(n_1950),
.B(n_1922),
.Y(n_2504)
);

NAND3xp33_ASAP7_75t_L g2505 ( 
.A(n_2142),
.B(n_727),
.C(n_728),
.Y(n_2505)
);

INVxp67_ASAP7_75t_SL g2506 ( 
.A(n_1923),
.Y(n_2506)
);

AOI21xp33_ASAP7_75t_L g2507 ( 
.A1(n_2089),
.A2(n_729),
.B(n_730),
.Y(n_2507)
);

BUFx3_ASAP7_75t_L g2508 ( 
.A(n_1955),
.Y(n_2508)
);

OAI21x1_ASAP7_75t_SL g2509 ( 
.A1(n_2069),
.A2(n_1921),
.B(n_1988),
.Y(n_2509)
);

AND2x4_ASAP7_75t_L g2510 ( 
.A(n_2034),
.B(n_731),
.Y(n_2510)
);

NAND2x1p5_ASAP7_75t_L g2511 ( 
.A(n_2066),
.B(n_731),
.Y(n_2511)
);

OAI21x1_ASAP7_75t_L g2512 ( 
.A1(n_1924),
.A2(n_733),
.B(n_734),
.Y(n_2512)
);

BUFx12f_ASAP7_75t_L g2513 ( 
.A(n_1952),
.Y(n_2513)
);

AOI22xp33_ASAP7_75t_L g2514 ( 
.A1(n_2124),
.A2(n_734),
.B1(n_735),
.B2(n_736),
.Y(n_2514)
);

OR2x2_ASAP7_75t_L g2515 ( 
.A(n_2075),
.B(n_736),
.Y(n_2515)
);

OAI21x1_ASAP7_75t_SL g2516 ( 
.A1(n_1921),
.A2(n_737),
.B(n_738),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2278),
.Y(n_2517)
);

AO31x2_ASAP7_75t_L g2518 ( 
.A1(n_2153),
.A2(n_737),
.A3(n_738),
.B(n_739),
.Y(n_2518)
);

INVx1_ASAP7_75t_SL g2519 ( 
.A(n_2066),
.Y(n_2519)
);

AOI21x1_ASAP7_75t_L g2520 ( 
.A1(n_1999),
.A2(n_741),
.B(n_742),
.Y(n_2520)
);

BUFx3_ASAP7_75t_L g2521 ( 
.A(n_2090),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_1954),
.Y(n_2522)
);

OA21x2_ASAP7_75t_L g2523 ( 
.A1(n_1912),
.A2(n_743),
.B(n_744),
.Y(n_2523)
);

AND2x2_ASAP7_75t_SL g2524 ( 
.A(n_2218),
.B(n_2076),
.Y(n_2524)
);

HB1xp67_ASAP7_75t_L g2525 ( 
.A(n_2064),
.Y(n_2525)
);

NOR2x1_ASAP7_75t_SL g2526 ( 
.A(n_1923),
.B(n_1940),
.Y(n_2526)
);

AOI21x1_ASAP7_75t_L g2527 ( 
.A1(n_2133),
.A2(n_745),
.B(n_746),
.Y(n_2527)
);

BUFx3_ASAP7_75t_L g2528 ( 
.A(n_2090),
.Y(n_2528)
);

HB1xp67_ASAP7_75t_L g2529 ( 
.A(n_2064),
.Y(n_2529)
);

OAI21x1_ASAP7_75t_SL g2530 ( 
.A1(n_2140),
.A2(n_746),
.B(n_747),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2056),
.B(n_747),
.Y(n_2531)
);

NOR2xp67_ASAP7_75t_L g2532 ( 
.A(n_2169),
.B(n_748),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2139),
.B(n_2161),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2054),
.Y(n_2534)
);

AOI22x1_ASAP7_75t_L g2535 ( 
.A1(n_2121),
.A2(n_750),
.B1(n_751),
.B2(n_752),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2029),
.Y(n_2536)
);

OAI21x1_ASAP7_75t_L g2537 ( 
.A1(n_2037),
.A2(n_753),
.B(n_754),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2029),
.Y(n_2538)
);

AOI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2057),
.A2(n_754),
.B(n_755),
.Y(n_2539)
);

OAI21x1_ASAP7_75t_L g2540 ( 
.A1(n_2044),
.A2(n_2074),
.B(n_1972),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2167),
.Y(n_2541)
);

BUFx2_ASAP7_75t_L g2542 ( 
.A(n_1911),
.Y(n_2542)
);

INVx6_ASAP7_75t_L g2543 ( 
.A(n_2127),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2180),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_L g2545 ( 
.A(n_1962),
.Y(n_2545)
);

BUFx2_ASAP7_75t_L g2546 ( 
.A(n_1911),
.Y(n_2546)
);

OA21x2_ASAP7_75t_L g2547 ( 
.A1(n_2074),
.A2(n_755),
.B(n_757),
.Y(n_2547)
);

NAND3xp33_ASAP7_75t_L g2548 ( 
.A(n_2187),
.B(n_2200),
.C(n_2189),
.Y(n_2548)
);

INVx6_ASAP7_75t_L g2549 ( 
.A(n_2227),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2085),
.B(n_757),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2232),
.B(n_758),
.Y(n_2551)
);

AOI22x1_ASAP7_75t_L g2552 ( 
.A1(n_2109),
.A2(n_758),
.B1(n_759),
.B2(n_760),
.Y(n_2552)
);

AOI22xp33_ASAP7_75t_L g2553 ( 
.A1(n_2019),
.A2(n_759),
.B1(n_760),
.B2(n_761),
.Y(n_2553)
);

INVx2_ASAP7_75t_SL g2554 ( 
.A(n_1930),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_1920),
.Y(n_2555)
);

OA21x2_ASAP7_75t_L g2556 ( 
.A1(n_1963),
.A2(n_762),
.B(n_763),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2268),
.Y(n_2557)
);

BUFx6f_ASAP7_75t_L g2558 ( 
.A(n_1978),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2272),
.Y(n_2559)
);

AO21x2_ASAP7_75t_L g2560 ( 
.A1(n_2176),
.A2(n_764),
.B(n_765),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_1940),
.Y(n_2561)
);

AO21x2_ASAP7_75t_L g2562 ( 
.A1(n_2176),
.A2(n_764),
.B(n_765),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2147),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2230),
.Y(n_2564)
);

NAND2x1p5_ASAP7_75t_L g2565 ( 
.A(n_2171),
.B(n_766),
.Y(n_2565)
);

BUFx3_ASAP7_75t_L g2566 ( 
.A(n_2171),
.Y(n_2566)
);

INVxp67_ASAP7_75t_SL g2567 ( 
.A(n_1916),
.Y(n_2567)
);

OAI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2040),
.A2(n_2079),
.B(n_2068),
.Y(n_2568)
);

BUFx3_ASAP7_75t_L g2569 ( 
.A(n_2190),
.Y(n_2569)
);

AOI221xp5_ASAP7_75t_SL g2570 ( 
.A1(n_1989),
.A2(n_768),
.B1(n_769),
.B2(n_770),
.C(n_771),
.Y(n_2570)
);

AO21x2_ASAP7_75t_L g2571 ( 
.A1(n_1985),
.A2(n_769),
.B(n_770),
.Y(n_2571)
);

NAND2x1p5_ASAP7_75t_L g2572 ( 
.A(n_2190),
.B(n_771),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2032),
.Y(n_2573)
);

OAI21x1_ASAP7_75t_L g2574 ( 
.A1(n_2141),
.A2(n_773),
.B(n_775),
.Y(n_2574)
);

HB1xp67_ASAP7_75t_L g2575 ( 
.A(n_2092),
.Y(n_2575)
);

BUFx2_ASAP7_75t_L g2576 ( 
.A(n_1930),
.Y(n_2576)
);

A2O1A1Ixp33_ASAP7_75t_L g2577 ( 
.A1(n_1995),
.A2(n_773),
.B(n_775),
.C(n_777),
.Y(n_2577)
);

OAI21x1_ASAP7_75t_L g2578 ( 
.A1(n_2228),
.A2(n_779),
.B(n_780),
.Y(n_2578)
);

OAI21x1_ASAP7_75t_L g2579 ( 
.A1(n_2229),
.A2(n_781),
.B(n_783),
.Y(n_2579)
);

INVx2_ASAP7_75t_SL g2580 ( 
.A(n_1939),
.Y(n_2580)
);

OAI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2040),
.A2(n_781),
.B(n_2079),
.Y(n_2581)
);

BUFx12f_ASAP7_75t_L g2582 ( 
.A(n_1939),
.Y(n_2582)
);

INVx4_ASAP7_75t_L g2583 ( 
.A(n_2001),
.Y(n_2583)
);

BUFx2_ASAP7_75t_L g2584 ( 
.A(n_2001),
.Y(n_2584)
);

AO21x2_ASAP7_75t_L g2585 ( 
.A1(n_2109),
.A2(n_2038),
.B(n_2033),
.Y(n_2585)
);

BUFx3_ASAP7_75t_L g2586 ( 
.A(n_2251),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_2032),
.Y(n_2587)
);

BUFx6f_ASAP7_75t_L g2588 ( 
.A(n_2251),
.Y(n_2588)
);

OAI21x1_ASAP7_75t_L g2589 ( 
.A1(n_2138),
.A2(n_2151),
.B(n_2145),
.Y(n_2589)
);

BUFx2_ASAP7_75t_L g2590 ( 
.A(n_2255),
.Y(n_2590)
);

OAI21x1_ASAP7_75t_L g2591 ( 
.A1(n_2155),
.A2(n_2173),
.B(n_2163),
.Y(n_2591)
);

OAI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2063),
.A2(n_2072),
.B(n_2068),
.Y(n_2592)
);

OAI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_1916),
.A2(n_1965),
.B1(n_1974),
.B2(n_1968),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2036),
.B(n_2050),
.Y(n_2594)
);

NAND3xp33_ASAP7_75t_L g2595 ( 
.A(n_2265),
.B(n_2269),
.C(n_2128),
.Y(n_2595)
);

OR2x6_ASAP7_75t_L g2596 ( 
.A(n_2255),
.B(n_2257),
.Y(n_2596)
);

OAI21x1_ASAP7_75t_L g2597 ( 
.A1(n_2185),
.A2(n_2220),
.B(n_2205),
.Y(n_2597)
);

OAI21x1_ASAP7_75t_L g2598 ( 
.A1(n_2222),
.A2(n_2243),
.B(n_2235),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2233),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_1915),
.Y(n_2600)
);

OAI21x1_ASAP7_75t_L g2601 ( 
.A1(n_2244),
.A2(n_2264),
.B(n_2259),
.Y(n_2601)
);

INVx3_ASAP7_75t_L g2602 ( 
.A(n_2257),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2060),
.Y(n_2603)
);

OAI21x1_ASAP7_75t_L g2604 ( 
.A1(n_2276),
.A2(n_2281),
.B(n_2279),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2260),
.B(n_2267),
.Y(n_2605)
);

BUFx6f_ASAP7_75t_L g2606 ( 
.A(n_1935),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2055),
.B(n_2077),
.Y(n_2607)
);

BUFx2_ASAP7_75t_R g2608 ( 
.A(n_2108),
.Y(n_2608)
);

AO31x2_ASAP7_75t_L g2609 ( 
.A1(n_2097),
.A2(n_1968),
.A3(n_1965),
.B(n_2052),
.Y(n_2609)
);

AO21x2_ASAP7_75t_L g2610 ( 
.A1(n_2033),
.A2(n_2041),
.B(n_2038),
.Y(n_2610)
);

AO21x2_ASAP7_75t_L g2611 ( 
.A1(n_2041),
.A2(n_2067),
.B(n_1964),
.Y(n_2611)
);

AO21x2_ASAP7_75t_L g2612 ( 
.A1(n_1963),
.A2(n_1975),
.B(n_1964),
.Y(n_2612)
);

HB1xp67_ASAP7_75t_L g2613 ( 
.A(n_2104),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2043),
.B(n_2094),
.Y(n_2614)
);

NAND2x1_ASAP7_75t_L g2615 ( 
.A(n_2065),
.B(n_2106),
.Y(n_2615)
);

NAND2x1p5_ASAP7_75t_L g2616 ( 
.A(n_2062),
.B(n_2125),
.Y(n_2616)
);

HB1xp67_ASAP7_75t_L g2617 ( 
.A(n_2104),
.Y(n_2617)
);

NAND2x1_ASAP7_75t_L g2618 ( 
.A(n_2106),
.B(n_2105),
.Y(n_2618)
);

OA21x2_ASAP7_75t_L g2619 ( 
.A1(n_2204),
.A2(n_2208),
.B(n_1953),
.Y(n_2619)
);

OAI21x1_ASAP7_75t_L g2620 ( 
.A1(n_2051),
.A2(n_1996),
.B(n_2004),
.Y(n_2620)
);

INVx2_ASAP7_75t_SL g2621 ( 
.A(n_2053),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2236),
.Y(n_2622)
);

INVx4_ASAP7_75t_L g2623 ( 
.A(n_2019),
.Y(n_2623)
);

BUFx3_ASAP7_75t_L g2624 ( 
.A(n_2110),
.Y(n_2624)
);

OAI21xp5_ASAP7_75t_L g2625 ( 
.A1(n_2063),
.A2(n_2072),
.B(n_1977),
.Y(n_2625)
);

AO21x2_ASAP7_75t_L g2626 ( 
.A1(n_2013),
.A2(n_1992),
.B(n_2046),
.Y(n_2626)
);

AO21x1_ASAP7_75t_L g2627 ( 
.A1(n_2201),
.A2(n_2280),
.B(n_2256),
.Y(n_2627)
);

OA21x2_ASAP7_75t_L g2628 ( 
.A1(n_1992),
.A2(n_2046),
.B(n_2042),
.Y(n_2628)
);

OAI21x1_ASAP7_75t_SL g2629 ( 
.A1(n_2186),
.A2(n_2215),
.B(n_2270),
.Y(n_2629)
);

OR2x6_ASAP7_75t_L g2630 ( 
.A(n_2221),
.B(n_2245),
.Y(n_2630)
);

BUFx12f_ASAP7_75t_L g2631 ( 
.A(n_2114),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_SL g2632 ( 
.A(n_2058),
.B(n_2201),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2582),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2291),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2295),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2286),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2310),
.Y(n_2637)
);

NAND2x1p5_ASAP7_75t_L g2638 ( 
.A(n_2292),
.B(n_2112),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2321),
.Y(n_2639)
);

OAI21x1_ASAP7_75t_SL g2640 ( 
.A1(n_2526),
.A2(n_2003),
.B(n_2280),
.Y(n_2640)
);

OAI22xp5_ASAP7_75t_L g2641 ( 
.A1(n_2573),
.A2(n_2256),
.B1(n_2195),
.B2(n_2231),
.Y(n_2641)
);

BUFx3_ASAP7_75t_L g2642 ( 
.A(n_2415),
.Y(n_2642)
);

OAI21x1_ASAP7_75t_SL g2643 ( 
.A1(n_2627),
.A2(n_2042),
.B(n_2103),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2325),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2534),
.Y(n_2645)
);

AOI22xp33_ASAP7_75t_L g2646 ( 
.A1(n_2573),
.A2(n_2231),
.B1(n_2195),
.B2(n_2282),
.Y(n_2646)
);

BUFx2_ASAP7_75t_L g2647 ( 
.A(n_2582),
.Y(n_2647)
);

BUFx3_ASAP7_75t_L g2648 ( 
.A(n_2415),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2534),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_SL g2650 ( 
.A1(n_2587),
.A2(n_2103),
.B1(n_2031),
.B2(n_2134),
.Y(n_2650)
);

AOI22xp33_ASAP7_75t_SL g2651 ( 
.A1(n_2587),
.A2(n_2059),
.B1(n_2008),
.B2(n_2010),
.Y(n_2651)
);

BUFx3_ASAP7_75t_L g2652 ( 
.A(n_2415),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2286),
.Y(n_2653)
);

OA21x2_ASAP7_75t_L g2654 ( 
.A1(n_2369),
.A2(n_2022),
.B(n_2253),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2288),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2296),
.Y(n_2656)
);

BUFx3_ASAP7_75t_L g2657 ( 
.A(n_2468),
.Y(n_2657)
);

BUFx2_ASAP7_75t_L g2658 ( 
.A(n_2483),
.Y(n_2658)
);

INVx6_ASAP7_75t_L g2659 ( 
.A(n_2329),
.Y(n_2659)
);

INVx3_ASAP7_75t_L g2660 ( 
.A(n_2583),
.Y(n_2660)
);

AOI22xp33_ASAP7_75t_L g2661 ( 
.A1(n_2630),
.A2(n_2506),
.B1(n_2479),
.B2(n_2631),
.Y(n_2661)
);

OA21x2_ASAP7_75t_L g2662 ( 
.A1(n_2293),
.A2(n_2022),
.B(n_2253),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2303),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2317),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2336),
.Y(n_2665)
);

BUFx10_ASAP7_75t_L g2666 ( 
.A(n_2312),
.Y(n_2666)
);

AND2x2_ASAP7_75t_L g2667 ( 
.A(n_2391),
.B(n_2300),
.Y(n_2667)
);

BUFx3_ASAP7_75t_L g2668 ( 
.A(n_2468),
.Y(n_2668)
);

NAND2x1p5_ASAP7_75t_L g2669 ( 
.A(n_2292),
.B(n_2091),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2555),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2555),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2603),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_2292),
.Y(n_2673)
);

BUFx2_ASAP7_75t_L g2674 ( 
.A(n_2483),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2339),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2561),
.B(n_2087),
.Y(n_2676)
);

INVx1_ASAP7_75t_SL g2677 ( 
.A(n_2478),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2391),
.B(n_2078),
.Y(n_2678)
);

AND2x4_ASAP7_75t_L g2679 ( 
.A(n_2596),
.B(n_2583),
.Y(n_2679)
);

AOI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2605),
.A2(n_1941),
.B1(n_1980),
.B2(n_1982),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2300),
.B(n_2011),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_2326),
.Y(n_2682)
);

OR2x2_ASAP7_75t_L g2683 ( 
.A(n_2307),
.B(n_2238),
.Y(n_2683)
);

INVx1_ASAP7_75t_SL g2684 ( 
.A(n_2500),
.Y(n_2684)
);

INVx2_ASAP7_75t_SL g2685 ( 
.A(n_2302),
.Y(n_2685)
);

OAI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_2500),
.A2(n_2122),
.B1(n_1970),
.B2(n_2181),
.Y(n_2686)
);

AOI22xp33_ASAP7_75t_L g2687 ( 
.A1(n_2630),
.A2(n_1933),
.B1(n_2209),
.B2(n_1918),
.Y(n_2687)
);

BUFx6f_ASAP7_75t_SL g2688 ( 
.A(n_2327),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2309),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_L g2690 ( 
.A1(n_2630),
.A2(n_1918),
.B1(n_2209),
.B2(n_2213),
.Y(n_2690)
);

INVx4_ASAP7_75t_SL g2691 ( 
.A(n_2596),
.Y(n_2691)
);

INVx3_ASAP7_75t_L g2692 ( 
.A(n_2326),
.Y(n_2692)
);

AOI22xp33_ASAP7_75t_SL g2693 ( 
.A1(n_2506),
.A2(n_2095),
.B1(n_2131),
.B2(n_2000),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2510),
.Y(n_2694)
);

AOI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_2631),
.A2(n_2213),
.B1(n_2006),
.B2(n_2247),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2510),
.Y(n_2696)
);

BUFx2_ASAP7_75t_SL g2697 ( 
.A(n_2327),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2525),
.Y(n_2698)
);

HB1xp67_ASAP7_75t_L g2699 ( 
.A(n_2525),
.Y(n_2699)
);

AOI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2605),
.A2(n_2047),
.B1(n_1998),
.B2(n_1925),
.Y(n_2700)
);

INVx3_ASAP7_75t_L g2701 ( 
.A(n_2326),
.Y(n_2701)
);

OR2x2_ASAP7_75t_L g2702 ( 
.A(n_2331),
.B(n_2271),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2493),
.B(n_2100),
.Y(n_2703)
);

OR2x2_ASAP7_75t_L g2704 ( 
.A(n_2421),
.B(n_2087),
.Y(n_2704)
);

AOI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2337),
.A2(n_2160),
.B1(n_2165),
.B2(n_2193),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2623),
.A2(n_2123),
.B1(n_1981),
.B2(n_2018),
.Y(n_2706)
);

BUFx3_ASAP7_75t_L g2707 ( 
.A(n_2381),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2537),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2345),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2537),
.Y(n_2710)
);

INVx2_ASAP7_75t_SL g2711 ( 
.A(n_2328),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2323),
.B(n_2035),
.Y(n_2712)
);

HB1xp67_ASAP7_75t_L g2713 ( 
.A(n_2529),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2511),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2511),
.Y(n_2715)
);

BUFx3_ASAP7_75t_L g2716 ( 
.A(n_2381),
.Y(n_2716)
);

BUFx3_ASAP7_75t_L g2717 ( 
.A(n_2463),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2485),
.B(n_2048),
.Y(n_2718)
);

OAI21xp5_ASAP7_75t_L g2719 ( 
.A1(n_2593),
.A2(n_2018),
.B(n_2023),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_2513),
.Y(n_2720)
);

AOI22xp33_ASAP7_75t_SL g2721 ( 
.A1(n_2304),
.A2(n_2020),
.B1(n_2214),
.B2(n_2137),
.Y(n_2721)
);

BUFx3_ASAP7_75t_L g2722 ( 
.A(n_2463),
.Y(n_2722)
);

INVx2_ASAP7_75t_SL g2723 ( 
.A(n_2329),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2441),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2495),
.B(n_2009),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2441),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_SL g2727 ( 
.A(n_2524),
.Y(n_2727)
);

AND2x4_ASAP7_75t_L g2728 ( 
.A(n_2596),
.B(n_2024),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2456),
.Y(n_2729)
);

BUFx2_ASAP7_75t_L g2730 ( 
.A(n_2513),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2456),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2498),
.Y(n_2732)
);

NAND2x1p5_ASAP7_75t_L g2733 ( 
.A(n_2348),
.B(n_1947),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2567),
.B(n_1919),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2567),
.B(n_1919),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2522),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2498),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2348),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2565),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2565),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2522),
.Y(n_2741)
);

HB1xp67_ASAP7_75t_L g2742 ( 
.A(n_2529),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2572),
.Y(n_2743)
);

NAND2x1p5_ASAP7_75t_L g2744 ( 
.A(n_2332),
.B(n_2020),
.Y(n_2744)
);

BUFx3_ASAP7_75t_L g2745 ( 
.A(n_2319),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2350),
.B(n_1919),
.Y(n_2746)
);

INVxp67_ASAP7_75t_L g2747 ( 
.A(n_2289),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2572),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2362),
.Y(n_2749)
);

OAI221xp5_ASAP7_75t_L g2750 ( 
.A1(n_2414),
.A2(n_2437),
.B1(n_2614),
.B2(n_2607),
.C(n_2632),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2522),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_SL g2752 ( 
.A1(n_2304),
.A2(n_2102),
.B1(n_2025),
.B2(n_2039),
.Y(n_2752)
);

BUFx2_ASAP7_75t_L g2753 ( 
.A(n_2542),
.Y(n_2753)
);

AOI22xp33_ASAP7_75t_L g2754 ( 
.A1(n_2623),
.A2(n_2071),
.B1(n_2073),
.B2(n_2111),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2489),
.B(n_2005),
.Y(n_2755)
);

NOR2x1_ASAP7_75t_R g2756 ( 
.A(n_2297),
.B(n_1928),
.Y(n_2756)
);

INVx3_ASAP7_75t_L g2757 ( 
.A(n_2332),
.Y(n_2757)
);

BUFx4f_ASAP7_75t_SL g2758 ( 
.A(n_2347),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2362),
.Y(n_2759)
);

BUFx4f_ASAP7_75t_L g2760 ( 
.A(n_2347),
.Y(n_2760)
);

AO21x2_ASAP7_75t_L g2761 ( 
.A1(n_2509),
.A2(n_2120),
.B(n_2152),
.Y(n_2761)
);

INVx2_ASAP7_75t_SL g2762 ( 
.A(n_2377),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2341),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2359),
.B(n_1928),
.Y(n_2764)
);

INVx3_ASAP7_75t_L g2765 ( 
.A(n_2334),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2430),
.Y(n_2766)
);

BUFx3_ASAP7_75t_L g2767 ( 
.A(n_2319),
.Y(n_2767)
);

INVx1_ASAP7_75t_SL g2768 ( 
.A(n_2519),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2334),
.Y(n_2769)
);

BUFx3_ASAP7_75t_L g2770 ( 
.A(n_2333),
.Y(n_2770)
);

HB1xp67_ASAP7_75t_L g2771 ( 
.A(n_2351),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2457),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2289),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2315),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2388),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2366),
.B(n_2223),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2299),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2442),
.A2(n_2166),
.B1(n_2223),
.B2(n_2275),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2474),
.B(n_2275),
.Y(n_2779)
);

NAND2x1_ASAP7_75t_L g2780 ( 
.A(n_2491),
.B(n_2275),
.Y(n_2780)
);

BUFx12f_ASAP7_75t_L g2781 ( 
.A(n_2312),
.Y(n_2781)
);

AO21x1_ASAP7_75t_SL g2782 ( 
.A1(n_2613),
.A2(n_2135),
.B(n_2021),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2420),
.B(n_2021),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2613),
.Y(n_2784)
);

OAI21x1_ASAP7_75t_L g2785 ( 
.A1(n_2540),
.A2(n_2135),
.B(n_2021),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2617),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2617),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2546),
.Y(n_2788)
);

OA21x2_ASAP7_75t_L g2789 ( 
.A1(n_2504),
.A2(n_2135),
.B(n_2301),
.Y(n_2789)
);

INVx2_ASAP7_75t_SL g2790 ( 
.A(n_2377),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2576),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2584),
.Y(n_2792)
);

INVx4_ASAP7_75t_L g2793 ( 
.A(n_2297),
.Y(n_2793)
);

HB1xp67_ASAP7_75t_L g2794 ( 
.A(n_2351),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2590),
.Y(n_2795)
);

AOI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_2594),
.A2(n_2497),
.B1(n_2550),
.B2(n_2460),
.Y(n_2796)
);

INVx1_ASAP7_75t_SL g2797 ( 
.A(n_2624),
.Y(n_2797)
);

INVxp67_ASAP7_75t_L g2798 ( 
.A(n_2460),
.Y(n_2798)
);

CKINVDCx6p67_ASAP7_75t_R g2799 ( 
.A(n_2335),
.Y(n_2799)
);

INVx4_ASAP7_75t_SL g2800 ( 
.A(n_2333),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2461),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2461),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2473),
.B(n_2502),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2624),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2438),
.Y(n_2805)
);

CKINVDCx11_ASAP7_75t_R g2806 ( 
.A(n_2318),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2438),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2438),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2424),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2545),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2541),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_2318),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2544),
.Y(n_2813)
);

NAND2x1p5_ASAP7_75t_L g2814 ( 
.A(n_2602),
.B(n_2476),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2557),
.Y(n_2815)
);

BUFx2_ASAP7_75t_L g2816 ( 
.A(n_2400),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2558),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2559),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2494),
.Y(n_2819)
);

INVx4_ASAP7_75t_L g2820 ( 
.A(n_2380),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2376),
.B(n_2515),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2558),
.Y(n_2822)
);

CKINVDCx5p33_ASAP7_75t_R g2823 ( 
.A(n_2361),
.Y(n_2823)
);

INVx1_ASAP7_75t_SL g2824 ( 
.A(n_2412),
.Y(n_2824)
);

INVx1_ASAP7_75t_SL g2825 ( 
.A(n_2412),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2532),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2574),
.Y(n_2827)
);

INVxp67_ASAP7_75t_L g2828 ( 
.A(n_2305),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2578),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2558),
.Y(n_2830)
);

AND2x4_ASAP7_75t_L g2831 ( 
.A(n_2602),
.B(n_2476),
.Y(n_2831)
);

HB1xp67_ASAP7_75t_L g2832 ( 
.A(n_2575),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2579),
.Y(n_2833)
);

AO21x2_ASAP7_75t_L g2834 ( 
.A1(n_2436),
.A2(n_2444),
.B(n_2439),
.Y(n_2834)
);

NAND2x1p5_ASAP7_75t_L g2835 ( 
.A(n_2554),
.B(n_2580),
.Y(n_2835)
);

INVx4_ASAP7_75t_L g2836 ( 
.A(n_2380),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2384),
.Y(n_2837)
);

HB1xp67_ASAP7_75t_L g2838 ( 
.A(n_2575),
.Y(n_2838)
);

BUFx3_ASAP7_75t_L g2839 ( 
.A(n_2353),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2376),
.Y(n_2840)
);

BUFx2_ASAP7_75t_L g2841 ( 
.A(n_2400),
.Y(n_2841)
);

HB1xp67_ASAP7_75t_L g2842 ( 
.A(n_2484),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_2484),
.Y(n_2843)
);

HB1xp67_ASAP7_75t_L g2844 ( 
.A(n_2404),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2290),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2550),
.B(n_2621),
.Y(n_2846)
);

AOI22xp33_ASAP7_75t_SL g2847 ( 
.A1(n_2552),
.A2(n_2497),
.B1(n_2524),
.B2(n_2516),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2443),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2535),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2446),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2353),
.Y(n_2851)
);

OR2x6_ASAP7_75t_L g2852 ( 
.A(n_2313),
.B(n_2322),
.Y(n_2852)
);

OAI21x1_ASAP7_75t_L g2853 ( 
.A1(n_2589),
.A2(n_2598),
.B(n_2597),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2499),
.B(n_2508),
.Y(n_2854)
);

CKINVDCx11_ASAP7_75t_R g2855 ( 
.A(n_2435),
.Y(n_2855)
);

BUFx2_ASAP7_75t_L g2856 ( 
.A(n_2397),
.Y(n_2856)
);

AOI22xp33_ASAP7_75t_SL g2857 ( 
.A1(n_2358),
.A2(n_2469),
.B1(n_2628),
.B2(n_2434),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2330),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2371),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2371),
.Y(n_2860)
);

BUFx2_ASAP7_75t_L g2861 ( 
.A(n_2429),
.Y(n_2861)
);

INVxp67_ASAP7_75t_SL g2862 ( 
.A(n_2501),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2360),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2371),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2434),
.B(n_2594),
.Y(n_2865)
);

OAI21x1_ASAP7_75t_L g2866 ( 
.A1(n_2589),
.A2(n_2598),
.B(n_2597),
.Y(n_2866)
);

INVx1_ASAP7_75t_SL g2867 ( 
.A(n_2360),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2370),
.B(n_2372),
.Y(n_2868)
);

CKINVDCx6p67_ASAP7_75t_R g2869 ( 
.A(n_2435),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2316),
.B(n_2514),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2316),
.B(n_2514),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2373),
.Y(n_2872)
);

CKINVDCx6p67_ASAP7_75t_R g2873 ( 
.A(n_2379),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2290),
.Y(n_2874)
);

INVx3_ASAP7_75t_L g2875 ( 
.A(n_2363),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2373),
.Y(n_2876)
);

OAI21x1_ASAP7_75t_L g2877 ( 
.A1(n_2601),
.A2(n_2604),
.B(n_2591),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2383),
.B(n_2386),
.Y(n_2878)
);

OAI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2481),
.A2(n_2553),
.B1(n_2501),
.B2(n_2322),
.Y(n_2879)
);

BUFx12f_ASAP7_75t_L g2880 ( 
.A(n_2361),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2390),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2393),
.Y(n_2882)
);

OAI21x1_ASAP7_75t_L g2883 ( 
.A1(n_2601),
.A2(n_2620),
.B(n_2346),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2394),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2499),
.B(n_2508),
.Y(n_2885)
);

HB1xp67_ASAP7_75t_L g2886 ( 
.A(n_2404),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2401),
.Y(n_2887)
);

INVx3_ASAP7_75t_L g2888 ( 
.A(n_2363),
.Y(n_2888)
);

BUFx10_ASAP7_75t_L g2889 ( 
.A(n_2287),
.Y(n_2889)
);

OAI33xp33_ASAP7_75t_L g2890 ( 
.A1(n_2496),
.A2(n_2531),
.A3(n_2477),
.B1(n_2419),
.B2(n_2285),
.B3(n_2392),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2407),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2368),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2409),
.B(n_2417),
.Y(n_2893)
);

BUFx8_ASAP7_75t_L g2894 ( 
.A(n_2294),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2425),
.Y(n_2895)
);

NAND2x1p5_ASAP7_75t_L g2896 ( 
.A(n_2368),
.B(n_2475),
.Y(n_2896)
);

AOI22xp5_ASAP7_75t_L g2897 ( 
.A1(n_2549),
.A2(n_2451),
.B1(n_2543),
.B2(n_2488),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2676),
.B(n_2536),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2655),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2803),
.B(n_2306),
.Y(n_2900)
);

NAND4xp25_ASAP7_75t_L g2901 ( 
.A(n_2865),
.B(n_2553),
.C(n_2408),
.D(n_2306),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2634),
.Y(n_2902)
);

INVx3_ASAP7_75t_L g2903 ( 
.A(n_2738),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_2865),
.A2(n_2612),
.B1(n_2462),
.B2(n_2449),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2821),
.B(n_2342),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2635),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2637),
.Y(n_2907)
);

AND2x4_ASAP7_75t_SL g2908 ( 
.A(n_2799),
.B(n_2447),
.Y(n_2908)
);

BUFx2_ASAP7_75t_L g2909 ( 
.A(n_2642),
.Y(n_2909)
);

AOI22xp33_ASAP7_75t_L g2910 ( 
.A1(n_2857),
.A2(n_2612),
.B1(n_2433),
.B2(n_2467),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2766),
.B(n_2352),
.Y(n_2911)
);

AOI22xp33_ASAP7_75t_L g2912 ( 
.A1(n_2857),
.A2(n_2517),
.B1(n_2440),
.B2(n_2453),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2747),
.B(n_2549),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2772),
.B(n_2396),
.Y(n_2914)
);

HB1xp67_ASAP7_75t_L g2915 ( 
.A(n_2636),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2639),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2676),
.B(n_2779),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2846),
.B(n_2410),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2644),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2811),
.Y(n_2920)
);

AOI22xp33_ASAP7_75t_L g2921 ( 
.A1(n_2870),
.A2(n_2432),
.B1(n_2450),
.B2(n_2466),
.Y(n_2921)
);

INVxp67_ASAP7_75t_L g2922 ( 
.A(n_2698),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2813),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2783),
.B(n_2538),
.Y(n_2924)
);

AOI22xp33_ASAP7_75t_SL g2925 ( 
.A1(n_2750),
.A2(n_2416),
.B1(n_2387),
.B2(n_2423),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2667),
.B(n_2447),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2775),
.B(n_2472),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2819),
.B(n_2698),
.Y(n_2928)
);

HB1xp67_ASAP7_75t_L g2929 ( 
.A(n_2673),
.Y(n_2929)
);

INVx3_ASAP7_75t_L g2930 ( 
.A(n_2738),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2699),
.B(n_2311),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2815),
.Y(n_2932)
);

BUFx3_ASAP7_75t_L g2933 ( 
.A(n_2642),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2713),
.B(n_2742),
.Y(n_2934)
);

AND2x4_ASAP7_75t_L g2935 ( 
.A(n_2691),
.B(n_2349),
.Y(n_2935)
);

BUFx3_ASAP7_75t_L g2936 ( 
.A(n_2648),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2871),
.A2(n_2455),
.B1(n_2428),
.B2(n_2426),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2713),
.B(n_2742),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2818),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2723),
.B(n_2543),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2797),
.B(n_2659),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2881),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2882),
.B(n_2609),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2884),
.Y(n_2944)
);

OAI22xp33_ASAP7_75t_L g2945 ( 
.A1(n_2750),
.A2(n_2581),
.B1(n_2314),
.B2(n_2470),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2797),
.B(n_2543),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2659),
.B(n_2482),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2887),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2891),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2659),
.B(n_2533),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2895),
.Y(n_2951)
);

BUFx3_ASAP7_75t_L g2952 ( 
.A(n_2648),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2645),
.Y(n_2953)
);

BUFx2_ASAP7_75t_SL g2954 ( 
.A(n_2652),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2657),
.B(n_2487),
.Y(n_2955)
);

AND2x2_ASAP7_75t_L g2956 ( 
.A(n_2657),
.B(n_2503),
.Y(n_2956)
);

AND2x4_ASAP7_75t_L g2957 ( 
.A(n_2691),
.B(n_2349),
.Y(n_2957)
);

OR2x2_ASAP7_75t_L g2958 ( 
.A(n_2649),
.B(n_2481),
.Y(n_2958)
);

BUFx2_ASAP7_75t_L g2959 ( 
.A(n_2652),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2653),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2668),
.B(n_2753),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_SL g2962 ( 
.A1(n_2879),
.A2(n_2678),
.B1(n_2641),
.B2(n_2640),
.Y(n_2962)
);

AND2x4_ASAP7_75t_L g2963 ( 
.A(n_2691),
.B(n_2374),
.Y(n_2963)
);

AOI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2850),
.A2(n_2599),
.B1(n_2622),
.B2(n_2563),
.Y(n_2964)
);

INVx2_ASAP7_75t_SL g2965 ( 
.A(n_2894),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2670),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2746),
.B(n_2609),
.Y(n_2967)
);

CKINVDCx5p33_ASAP7_75t_R g2968 ( 
.A(n_2806),
.Y(n_2968)
);

BUFx3_ASAP7_75t_L g2969 ( 
.A(n_2894),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2668),
.B(n_2451),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2671),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2704),
.B(n_2549),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2832),
.B(n_2571),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2832),
.B(n_2571),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2746),
.B(n_2609),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2838),
.B(n_2564),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2838),
.B(n_2551),
.Y(n_2977)
);

OR2x2_ASAP7_75t_L g2978 ( 
.A(n_2656),
.B(n_2560),
.Y(n_2978)
);

NOR2x1_ASAP7_75t_SL g2979 ( 
.A(n_2852),
.B(n_2305),
.Y(n_2979)
);

AOI22xp33_ASAP7_75t_L g2980 ( 
.A1(n_2641),
.A2(n_2625),
.B1(n_2592),
.B2(n_2568),
.Y(n_2980)
);

HB1xp67_ASAP7_75t_L g2981 ( 
.A(n_2673),
.Y(n_2981)
);

CKINVDCx14_ASAP7_75t_R g2982 ( 
.A(n_2806),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2661),
.B(n_2521),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2661),
.B(n_2521),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2672),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2868),
.Y(n_2986)
);

BUFx3_ASAP7_75t_L g2987 ( 
.A(n_2633),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2840),
.B(n_2528),
.Y(n_2988)
);

AND2x2_ASAP7_75t_SL g2989 ( 
.A(n_2816),
.B(n_2387),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2747),
.B(n_2528),
.Y(n_2990)
);

AOI222xp33_ASAP7_75t_L g2991 ( 
.A1(n_2861),
.A2(n_2758),
.B1(n_2760),
.B2(n_2647),
.C1(n_2646),
.C2(n_2687),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2868),
.Y(n_2992)
);

NOR2x1_ASAP7_75t_SL g2993 ( 
.A(n_2852),
.B(n_2491),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2878),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2718),
.B(n_2566),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2788),
.B(n_2569),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2791),
.B(n_2569),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2878),
.Y(n_2998)
);

OAI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2727),
.A2(n_2628),
.B1(n_2343),
.B2(n_2313),
.Y(n_2999)
);

NAND2x1_ASAP7_75t_L g3000 ( 
.A(n_2852),
.B(n_2629),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2727),
.A2(n_2343),
.B1(n_2556),
.B2(n_2547),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2893),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2792),
.B(n_2586),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2663),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2664),
.Y(n_3005)
);

CKINVDCx20_ASAP7_75t_R g3006 ( 
.A(n_2758),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2679),
.B(n_2374),
.Y(n_3007)
);

OAI21xp5_ASAP7_75t_SL g3008 ( 
.A1(n_2841),
.A2(n_2616),
.B(n_2385),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2795),
.B(n_2586),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2703),
.B(n_2395),
.Y(n_3010)
);

HB1xp67_ASAP7_75t_L g3011 ( 
.A(n_2771),
.Y(n_3011)
);

BUFx2_ASAP7_75t_L g3012 ( 
.A(n_2660),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2675),
.B(n_2507),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2764),
.B(n_2609),
.Y(n_3014)
);

INVx3_ASAP7_75t_L g3015 ( 
.A(n_2660),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2768),
.B(n_2560),
.Y(n_3016)
);

AND2x2_ASAP7_75t_L g3017 ( 
.A(n_2768),
.B(n_2562),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2665),
.Y(n_3018)
);

OR2x2_ASAP7_75t_L g3019 ( 
.A(n_2784),
.B(n_2562),
.Y(n_3019)
);

OR2x2_ASAP7_75t_L g3020 ( 
.A(n_2786),
.B(n_2518),
.Y(n_3020)
);

INVx3_ASAP7_75t_L g3021 ( 
.A(n_2682),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2845),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2787),
.B(n_2324),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2801),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2802),
.Y(n_3025)
);

INVx2_ASAP7_75t_SL g3026 ( 
.A(n_2889),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2771),
.B(n_2518),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2826),
.Y(n_3028)
);

HB1xp67_ASAP7_75t_L g3029 ( 
.A(n_2794),
.Y(n_3029)
);

HB1xp67_ASAP7_75t_L g3030 ( 
.A(n_2794),
.Y(n_3030)
);

OR2x2_ASAP7_75t_L g3031 ( 
.A(n_2804),
.B(n_2518),
.Y(n_3031)
);

BUFx3_ASAP7_75t_L g3032 ( 
.A(n_2873),
.Y(n_3032)
);

AND2x2_ASAP7_75t_L g3033 ( 
.A(n_2677),
.B(n_2796),
.Y(n_3033)
);

OAI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_2680),
.A2(n_2556),
.B1(n_2547),
.B2(n_2387),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2776),
.B(n_2610),
.Y(n_3035)
);

NOR2xp67_ASAP7_75t_SL g3036 ( 
.A(n_2697),
.B(n_2471),
.Y(n_3036)
);

AND2x2_ASAP7_75t_L g3037 ( 
.A(n_2677),
.B(n_2324),
.Y(n_3037)
);

INVx2_ASAP7_75t_SL g3038 ( 
.A(n_2889),
.Y(n_3038)
);

OAI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2690),
.A2(n_2556),
.B1(n_2547),
.B2(n_2406),
.Y(n_3039)
);

CKINVDCx20_ASAP7_75t_R g3040 ( 
.A(n_2855),
.Y(n_3040)
);

AND2x2_ASAP7_75t_L g3041 ( 
.A(n_2681),
.B(n_2777),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2724),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2844),
.Y(n_3043)
);

OR2x2_ASAP7_75t_L g3044 ( 
.A(n_2798),
.B(n_2518),
.Y(n_3044)
);

AND2x4_ASAP7_75t_L g3045 ( 
.A(n_2854),
.B(n_2402),
.Y(n_3045)
);

OAI22xp5_ASAP7_75t_L g3046 ( 
.A1(n_2690),
.A2(n_2399),
.B1(n_2480),
.B2(n_2423),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2773),
.B(n_2354),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2726),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2755),
.B(n_2725),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2837),
.B(n_2610),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2658),
.B(n_2354),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2729),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2674),
.B(n_2355),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2749),
.B(n_2626),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2874),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2759),
.B(n_2626),
.Y(n_3056)
);

HB1xp67_ASAP7_75t_L g3057 ( 
.A(n_2844),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2720),
.B(n_2355),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_SL g3059 ( 
.A1(n_2879),
.A2(n_2399),
.B1(n_2406),
.B2(n_2416),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2707),
.Y(n_3060)
);

OAI21xp33_ASAP7_75t_L g3061 ( 
.A1(n_2646),
.A2(n_2608),
.B(n_2577),
.Y(n_3061)
);

INVx4_ASAP7_75t_L g3062 ( 
.A(n_2820),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2731),
.Y(n_3063)
);

OAI21xp5_ASAP7_75t_SL g3064 ( 
.A1(n_2847),
.A2(n_2616),
.B(n_2385),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2730),
.B(n_2458),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2702),
.B(n_2422),
.Y(n_3066)
);

AOI22xp33_ASAP7_75t_L g3067 ( 
.A1(n_2848),
.A2(n_2548),
.B1(n_2611),
.B2(n_2585),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2732),
.Y(n_3068)
);

BUFx4f_ASAP7_75t_SL g3069 ( 
.A(n_2781),
.Y(n_3069)
);

HB1xp67_ASAP7_75t_L g3070 ( 
.A(n_2886),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2737),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2886),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2714),
.Y(n_3073)
);

BUFx3_ASAP7_75t_L g3074 ( 
.A(n_2707),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2715),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2694),
.B(n_2611),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2683),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2684),
.B(n_2398),
.Y(n_3078)
);

OAI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2687),
.A2(n_2423),
.B1(n_2399),
.B2(n_2406),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2842),
.Y(n_3080)
);

AND2x4_ASAP7_75t_L g3081 ( 
.A(n_2854),
.B(n_2402),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2763),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2842),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2843),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2696),
.B(n_2585),
.Y(n_3085)
);

BUFx2_ASAP7_75t_L g3086 ( 
.A(n_2885),
.Y(n_3086)
);

BUFx2_ASAP7_75t_L g3087 ( 
.A(n_2885),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_2684),
.B(n_2403),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2897),
.B(n_2418),
.Y(n_3089)
);

AND2x2_ASAP7_75t_L g3090 ( 
.A(n_2798),
.B(n_2588),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2843),
.Y(n_3091)
);

AND2x4_ASAP7_75t_L g3092 ( 
.A(n_2682),
.B(n_2475),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2809),
.Y(n_3093)
);

BUFx3_ASAP7_75t_L g3094 ( 
.A(n_2716),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2728),
.B(n_2820),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2728),
.B(n_2836),
.Y(n_3096)
);

OAI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_2705),
.A2(n_2480),
.B1(n_2416),
.B2(n_2344),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_L g3098 ( 
.A1(n_2643),
.A2(n_2357),
.B1(n_2389),
.B2(n_2452),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2836),
.B(n_2588),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2835),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2835),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2709),
.Y(n_3102)
);

INVx3_ASAP7_75t_L g3103 ( 
.A(n_2692),
.Y(n_3103)
);

HB1xp67_ASAP7_75t_L g3104 ( 
.A(n_2862),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2689),
.B(n_2298),
.Y(n_3105)
);

INVxp67_ASAP7_75t_L g3106 ( 
.A(n_2782),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_2855),
.Y(n_3107)
);

AND2x4_ASAP7_75t_L g3108 ( 
.A(n_2701),
.B(n_2800),
.Y(n_3108)
);

BUFx2_ASAP7_75t_L g3109 ( 
.A(n_2745),
.Y(n_3109)
);

BUFx3_ASAP7_75t_L g3110 ( 
.A(n_2716),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_SL g3111 ( 
.A(n_2862),
.B(n_2411),
.Y(n_3111)
);

BUFx2_ASAP7_75t_L g3112 ( 
.A(n_2745),
.Y(n_3112)
);

BUFx2_ASAP7_75t_L g3113 ( 
.A(n_2767),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2739),
.Y(n_3114)
);

OAI22xp5_ASAP7_75t_L g3115 ( 
.A1(n_2650),
.A2(n_2480),
.B1(n_2344),
.B2(n_2356),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2740),
.Y(n_3116)
);

CKINVDCx6p67_ASAP7_75t_R g3117 ( 
.A(n_2688),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2831),
.B(n_2298),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2743),
.Y(n_3119)
);

INVx3_ASAP7_75t_L g3120 ( 
.A(n_2701),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2831),
.B(n_2365),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2748),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2756),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2805),
.Y(n_3124)
);

BUFx2_ASAP7_75t_L g3125 ( 
.A(n_2767),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2717),
.B(n_2382),
.Y(n_3126)
);

AND2x4_ASAP7_75t_SL g3127 ( 
.A(n_2666),
.B(n_2491),
.Y(n_3127)
);

BUFx2_ASAP7_75t_L g3128 ( 
.A(n_2770),
.Y(n_3128)
);

INVx1_ASAP7_75t_SL g3129 ( 
.A(n_2867),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_2717),
.B(n_2382),
.Y(n_3130)
);

AOI22xp33_ASAP7_75t_SL g3131 ( 
.A1(n_2834),
.A2(n_2356),
.B1(n_2344),
.B2(n_2492),
.Y(n_3131)
);

NOR2x1_ASAP7_75t_L g3132 ( 
.A(n_2722),
.B(n_2389),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2722),
.B(n_2413),
.Y(n_3133)
);

HB1xp67_ASAP7_75t_L g3134 ( 
.A(n_2708),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2807),
.Y(n_3135)
);

BUFx2_ASAP7_75t_L g3136 ( 
.A(n_2770),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_2839),
.B(n_2413),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2808),
.Y(n_3138)
);

HB1xp67_ASAP7_75t_L g3139 ( 
.A(n_2710),
.Y(n_3139)
);

AND2x4_ASAP7_75t_L g3140 ( 
.A(n_2800),
.B(n_2405),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2839),
.B(n_2856),
.Y(n_3141)
);

INVx3_ASAP7_75t_L g3142 ( 
.A(n_2814),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2693),
.B(n_2427),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_3077),
.B(n_2734),
.Y(n_3144)
);

INVxp67_ASAP7_75t_L g3145 ( 
.A(n_2954),
.Y(n_3145)
);

AOI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_2991),
.A2(n_2695),
.B1(n_2686),
.B2(n_2700),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2928),
.B(n_2693),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2986),
.B(n_2712),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_3124),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_3135),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_3049),
.B(n_2867),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2992),
.B(n_2712),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3138),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2943),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_3106),
.B(n_3104),
.Y(n_3155)
);

OR2x2_ASAP7_75t_L g3156 ( 
.A(n_2917),
.B(n_2734),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_3041),
.B(n_2828),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2943),
.Y(n_3158)
);

HB1xp67_ASAP7_75t_L g3159 ( 
.A(n_2922),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_2972),
.B(n_2828),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_3106),
.B(n_2800),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_2926),
.B(n_2824),
.Y(n_3162)
);

CKINVDCx6p67_ASAP7_75t_R g3163 ( 
.A(n_2969),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_2995),
.B(n_2824),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2950),
.B(n_2825),
.Y(n_3165)
);

BUFx2_ASAP7_75t_SL g3166 ( 
.A(n_3006),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2902),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2994),
.B(n_2858),
.Y(n_3168)
);

HB1xp67_ASAP7_75t_L g3169 ( 
.A(n_2922),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2906),
.Y(n_3170)
);

AND2x2_ASAP7_75t_L g3171 ( 
.A(n_2976),
.B(n_2825),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2907),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2916),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2998),
.B(n_2859),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2919),
.Y(n_3175)
);

INVx3_ASAP7_75t_SL g3176 ( 
.A(n_3117),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_3033),
.B(n_2851),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_3062),
.B(n_2847),
.Y(n_3178)
);

AND2x4_ASAP7_75t_L g3179 ( 
.A(n_2934),
.B(n_2860),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2899),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_2941),
.B(n_2851),
.Y(n_3181)
);

AND2x4_ASAP7_75t_L g3182 ( 
.A(n_2938),
.B(n_2864),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2942),
.Y(n_3183)
);

AND2x2_ASAP7_75t_L g3184 ( 
.A(n_2961),
.B(n_2863),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2944),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2948),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_3109),
.B(n_2863),
.Y(n_3187)
);

AND2x2_ASAP7_75t_L g3188 ( 
.A(n_3112),
.B(n_2875),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2953),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3113),
.B(n_2875),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_3125),
.B(n_2888),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2949),
.Y(n_3192)
);

INVx3_ASAP7_75t_L g3193 ( 
.A(n_3062),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_3002),
.B(n_3102),
.Y(n_3194)
);

OR2x2_ASAP7_75t_L g3195 ( 
.A(n_2917),
.B(n_2735),
.Y(n_3195)
);

INVxp67_ASAP7_75t_SL g3196 ( 
.A(n_3057),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_3082),
.B(n_2872),
.Y(n_3197)
);

OR2x2_ASAP7_75t_L g3198 ( 
.A(n_2924),
.B(n_2735),
.Y(n_3198)
);

INVx3_ASAP7_75t_L g3199 ( 
.A(n_2903),
.Y(n_3199)
);

AND2x4_ASAP7_75t_SL g3200 ( 
.A(n_3006),
.B(n_2666),
.Y(n_3200)
);

NOR2x1_ASAP7_75t_SL g3201 ( 
.A(n_3008),
.B(n_2685),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2951),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2920),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2923),
.Y(n_3204)
);

OR2x6_ASAP7_75t_L g3205 ( 
.A(n_2969),
.B(n_2711),
.Y(n_3205)
);

INVxp67_ASAP7_75t_L g3206 ( 
.A(n_2987),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_3128),
.B(n_2888),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2921),
.B(n_2876),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2932),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_3136),
.B(n_2892),
.Y(n_3210)
);

OAI211xp5_ASAP7_75t_SL g3211 ( 
.A1(n_2991),
.A2(n_3028),
.B(n_3093),
.C(n_2904),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2966),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2971),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2985),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_3111),
.B(n_3012),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_3086),
.B(n_2892),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_SL g3217 ( 
.A(n_3111),
.B(n_2812),
.Y(n_3217)
);

AOI22xp33_ASAP7_75t_L g3218 ( 
.A1(n_3061),
.A2(n_2650),
.B1(n_2695),
.B2(n_2651),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3087),
.B(n_2834),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_2990),
.B(n_2736),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3004),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_2946),
.B(n_2741),
.Y(n_3222)
);

OAI21xp5_ASAP7_75t_L g3223 ( 
.A1(n_3089),
.A2(n_2651),
.B(n_2367),
.Y(n_3223)
);

AND2x4_ASAP7_75t_L g3224 ( 
.A(n_3080),
.B(n_3083),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2921),
.B(n_2778),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_3066),
.B(n_2751),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_2927),
.B(n_2977),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_2937),
.B(n_2778),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3005),
.Y(n_3229)
);

NOR2x1_ASAP7_75t_L g3230 ( 
.A(n_2933),
.B(n_2793),
.Y(n_3230)
);

INVx4_ASAP7_75t_L g3231 ( 
.A(n_2987),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2939),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2960),
.Y(n_3233)
);

AND2x4_ASAP7_75t_L g3234 ( 
.A(n_3084),
.B(n_2883),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2937),
.B(n_2719),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3024),
.Y(n_3236)
);

OR2x2_ASAP7_75t_L g3237 ( 
.A(n_2924),
.B(n_2869),
.Y(n_3237)
);

OR2x2_ASAP7_75t_L g3238 ( 
.A(n_2915),
.B(n_2785),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_3095),
.B(n_2810),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_3096),
.B(n_2817),
.Y(n_3240)
);

INVxp67_ASAP7_75t_SL g3241 ( 
.A(n_3057),
.Y(n_3241)
);

AOI22xp33_ASAP7_75t_L g3242 ( 
.A1(n_2962),
.A2(n_2686),
.B1(n_2890),
.B2(n_2530),
.Y(n_3242)
);

OR2x2_ASAP7_75t_L g3243 ( 
.A(n_2915),
.B(n_2744),
.Y(n_3243)
);

INVx4_ASAP7_75t_SL g3244 ( 
.A(n_3032),
.Y(n_3244)
);

NOR2xp67_ASAP7_75t_L g3245 ( 
.A(n_2965),
.B(n_2793),
.Y(n_3245)
);

OR2x2_ASAP7_75t_L g3246 ( 
.A(n_3011),
.B(n_2744),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3025),
.Y(n_3247)
);

NOR2x1_ASAP7_75t_SL g3248 ( 
.A(n_2933),
.B(n_2491),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3018),
.Y(n_3249)
);

HB1xp67_ASAP7_75t_L g3250 ( 
.A(n_3011),
.Y(n_3250)
);

AND2x2_ASAP7_75t_L g3251 ( 
.A(n_2988),
.B(n_2822),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_3051),
.B(n_2830),
.Y(n_3252)
);

NOR2xp33_ASAP7_75t_L g3253 ( 
.A(n_2909),
.B(n_2812),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_3053),
.B(n_2896),
.Y(n_3254)
);

OR2x2_ASAP7_75t_L g3255 ( 
.A(n_3029),
.B(n_2774),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3058),
.B(n_2896),
.Y(n_3256)
);

AND2x2_ASAP7_75t_L g3257 ( 
.A(n_3141),
.B(n_2719),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3091),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3029),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_2970),
.B(n_2814),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3022),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_2996),
.B(n_2654),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3022),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2911),
.B(n_2706),
.Y(n_3264)
);

OR2x2_ASAP7_75t_L g3265 ( 
.A(n_3030),
.B(n_2762),
.Y(n_3265)
);

BUFx6f_ASAP7_75t_L g3266 ( 
.A(n_2936),
.Y(n_3266)
);

OR2x2_ASAP7_75t_L g3267 ( 
.A(n_3030),
.B(n_2790),
.Y(n_3267)
);

AND2x4_ASAP7_75t_L g3268 ( 
.A(n_3126),
.B(n_2853),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2914),
.B(n_2905),
.Y(n_3269)
);

INVx1_ASAP7_75t_SL g3270 ( 
.A(n_3060),
.Y(n_3270)
);

OAI21xp5_ASAP7_75t_SL g3271 ( 
.A1(n_2962),
.A2(n_2638),
.B(n_2721),
.Y(n_3271)
);

BUFx2_ASAP7_75t_L g3272 ( 
.A(n_2936),
.Y(n_3272)
);

OR2x2_ASAP7_75t_L g3273 ( 
.A(n_3129),
.B(n_2638),
.Y(n_3273)
);

HB1xp67_ASAP7_75t_L g3274 ( 
.A(n_3070),
.Y(n_3274)
);

OR2x2_ASAP7_75t_L g3275 ( 
.A(n_3129),
.B(n_2789),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3114),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_L g3277 ( 
.A1(n_2901),
.A2(n_2890),
.B1(n_2721),
.B2(n_2752),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3116),
.Y(n_3278)
);

INVx2_ASAP7_75t_SL g3279 ( 
.A(n_3032),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3119),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3122),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_2959),
.B(n_2789),
.Y(n_3282)
);

HB1xp67_ASAP7_75t_L g3283 ( 
.A(n_3070),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2980),
.B(n_2706),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_2997),
.B(n_3003),
.Y(n_3285)
);

AND2x4_ASAP7_75t_L g3286 ( 
.A(n_3130),
.B(n_2866),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2980),
.B(n_2654),
.Y(n_3287)
);

AND2x2_ASAP7_75t_L g3288 ( 
.A(n_3009),
.B(n_3010),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_2904),
.B(n_2662),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3042),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2918),
.B(n_2662),
.Y(n_3291)
);

AND2x4_ASAP7_75t_L g3292 ( 
.A(n_3133),
.B(n_2877),
.Y(n_3292)
);

AOI22xp33_ASAP7_75t_SL g3293 ( 
.A1(n_2979),
.A2(n_2688),
.B1(n_2364),
.B2(n_2760),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3048),
.Y(n_3294)
);

OR2x2_ASAP7_75t_L g3295 ( 
.A(n_3043),
.B(n_3072),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2900),
.B(n_2570),
.Y(n_3296)
);

OAI222xp33_ASAP7_75t_L g3297 ( 
.A1(n_2912),
.A2(n_3000),
.B1(n_2910),
.B2(n_3123),
.C1(n_2982),
.C2(n_2999),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3052),
.Y(n_3298)
);

AND2x4_ASAP7_75t_L g3299 ( 
.A(n_3118),
.B(n_3037),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3063),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3068),
.B(n_2761),
.Y(n_3301)
);

AND2x2_ASAP7_75t_L g3302 ( 
.A(n_3071),
.B(n_2761),
.Y(n_3302)
);

NAND3xp33_ASAP7_75t_L g3303 ( 
.A(n_3089),
.B(n_2752),
.C(n_2754),
.Y(n_3303)
);

NOR2x1_ASAP7_75t_R g3304 ( 
.A(n_2968),
.B(n_2880),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3073),
.B(n_2780),
.Y(n_3305)
);

INVxp67_ASAP7_75t_SL g3306 ( 
.A(n_2929),
.Y(n_3306)
);

AND2x2_ASAP7_75t_L g3307 ( 
.A(n_3075),
.B(n_2827),
.Y(n_3307)
);

NOR2x1_ASAP7_75t_L g3308 ( 
.A(n_2952),
.B(n_2427),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3055),
.Y(n_3309)
);

AOI222xp33_ASAP7_75t_L g3310 ( 
.A1(n_2912),
.A2(n_2505),
.B1(n_2754),
.B2(n_2595),
.C1(n_2471),
.C2(n_2486),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3090),
.B(n_2829),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_2955),
.B(n_2833),
.Y(n_3312)
);

AND2x2_ASAP7_75t_L g3313 ( 
.A(n_2956),
.B(n_2952),
.Y(n_3313)
);

AND2x2_ASAP7_75t_L g3314 ( 
.A(n_2913),
.B(n_2364),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_3262),
.B(n_3016),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_3299),
.B(n_3017),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_3299),
.B(n_3047),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3167),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_L g3319 ( 
.A(n_3211),
.B(n_3013),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_3261),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3261),
.Y(n_3321)
);

AND2x2_ASAP7_75t_L g3322 ( 
.A(n_3312),
.B(n_3105),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3269),
.B(n_3023),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3257),
.B(n_3067),
.Y(n_3324)
);

NAND3xp33_ASAP7_75t_L g3325 ( 
.A(n_3303),
.B(n_2910),
.C(n_3067),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3170),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_3264),
.B(n_2973),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3301),
.B(n_2974),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_3146),
.B(n_2913),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3263),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3172),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_3302),
.B(n_3121),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3291),
.B(n_3031),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3173),
.Y(n_3334)
);

INVx2_ASAP7_75t_L g3335 ( 
.A(n_3263),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3252),
.B(n_2967),
.Y(n_3336)
);

AND2x4_ASAP7_75t_L g3337 ( 
.A(n_3268),
.B(n_3137),
.Y(n_3337)
);

OAI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3218),
.A2(n_2982),
.B1(n_3064),
.B2(n_2964),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3157),
.B(n_2964),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_3314),
.B(n_2967),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_3268),
.B(n_2975),
.Y(n_3341)
);

OR2x2_ASAP7_75t_L g3342 ( 
.A(n_3156),
.B(n_2929),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3175),
.Y(n_3343)
);

OR2x2_ASAP7_75t_L g3344 ( 
.A(n_3195),
.B(n_2981),
.Y(n_3344)
);

INVx1_ASAP7_75t_SL g3345 ( 
.A(n_3163),
.Y(n_3345)
);

BUFx2_ASAP7_75t_L g3346 ( 
.A(n_3231),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3180),
.Y(n_3347)
);

BUFx2_ASAP7_75t_L g3348 ( 
.A(n_3231),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3183),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3286),
.B(n_2975),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3185),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3186),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_3286),
.B(n_3014),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3192),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3202),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3154),
.B(n_3014),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3203),
.Y(n_3357)
);

OR2x2_ASAP7_75t_L g3358 ( 
.A(n_3144),
.B(n_3027),
.Y(n_3358)
);

BUFx3_ASAP7_75t_L g3359 ( 
.A(n_3193),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3154),
.B(n_3158),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3158),
.B(n_3311),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_3284),
.B(n_3060),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3292),
.B(n_3076),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3292),
.B(n_3076),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_3227),
.B(n_3134),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3179),
.B(n_3134),
.Y(n_3366)
);

OR2x2_ASAP7_75t_L g3367 ( 
.A(n_3198),
.B(n_3085),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3179),
.B(n_3139),
.Y(n_3368)
);

NOR2x1_ASAP7_75t_L g3369 ( 
.A(n_3193),
.B(n_3245),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3204),
.Y(n_3370)
);

AND2x2_ASAP7_75t_L g3371 ( 
.A(n_3182),
.B(n_3139),
.Y(n_3371)
);

AND2x2_ASAP7_75t_L g3372 ( 
.A(n_3182),
.B(n_3035),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3209),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3232),
.Y(n_3374)
);

BUFx2_ASAP7_75t_L g3375 ( 
.A(n_3272),
.Y(n_3375)
);

NAND2x1_ASAP7_75t_SL g3376 ( 
.A(n_3176),
.B(n_2903),
.Y(n_3376)
);

HB1xp67_ASAP7_75t_L g3377 ( 
.A(n_3274),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3224),
.B(n_2978),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3219),
.B(n_3035),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3233),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3307),
.B(n_3054),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_3313),
.B(n_3054),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_3234),
.B(n_3056),
.Y(n_3383)
);

INVx2_ASAP7_75t_SL g3384 ( 
.A(n_3155),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3236),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3234),
.B(n_3056),
.Y(n_3386)
);

AND2x2_ASAP7_75t_L g3387 ( 
.A(n_3309),
.B(n_3085),
.Y(n_3387)
);

OAI221xp5_ASAP7_75t_SL g3388 ( 
.A1(n_3271),
.A2(n_3277),
.B1(n_3242),
.B2(n_3235),
.C(n_3287),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3247),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3276),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3224),
.B(n_3019),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3278),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3280),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3281),
.Y(n_3394)
);

NAND2x1_ASAP7_75t_L g3395 ( 
.A(n_3161),
.B(n_3036),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3290),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3258),
.B(n_3020),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3294),
.Y(n_3398)
);

NOR3xp33_ASAP7_75t_L g3399 ( 
.A(n_3297),
.B(n_2945),
.C(n_3026),
.Y(n_3399)
);

HB1xp67_ASAP7_75t_L g3400 ( 
.A(n_3283),
.Y(n_3400)
);

INVx4_ASAP7_75t_L g3401 ( 
.A(n_3161),
.Y(n_3401)
);

AND2x2_ASAP7_75t_L g3402 ( 
.A(n_3316),
.B(n_3285),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3318),
.Y(n_3403)
);

INVx3_ASAP7_75t_L g3404 ( 
.A(n_3401),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3316),
.B(n_3177),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3326),
.Y(n_3406)
);

INVxp33_ASAP7_75t_L g3407 ( 
.A(n_3395),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3360),
.B(n_3333),
.Y(n_3408)
);

NAND4xp75_ASAP7_75t_L g3409 ( 
.A(n_3369),
.B(n_3217),
.C(n_3230),
.D(n_3178),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3331),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3320),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_3388),
.B(n_3237),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3334),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3320),
.Y(n_3414)
);

OR2x2_ASAP7_75t_L g3415 ( 
.A(n_3365),
.B(n_3250),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_3321),
.Y(n_3416)
);

OAI22xp33_ASAP7_75t_L g3417 ( 
.A1(n_3338),
.A2(n_3215),
.B1(n_3270),
.B2(n_3223),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3321),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3343),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3360),
.B(n_3259),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3347),
.Y(n_3421)
);

NAND2xp33_ASAP7_75t_R g3422 ( 
.A(n_3346),
.B(n_3348),
.Y(n_3422)
);

NOR2x1p5_ASAP7_75t_L g3423 ( 
.A(n_3401),
.B(n_3359),
.Y(n_3423)
);

INVx1_ASAP7_75t_SL g3424 ( 
.A(n_3345),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3317),
.B(n_3288),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3349),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_3330),
.Y(n_3427)
);

OAI21xp33_ASAP7_75t_L g3428 ( 
.A1(n_3319),
.A2(n_3399),
.B(n_3325),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3317),
.B(n_3151),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3351),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3365),
.B(n_3254),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3315),
.B(n_3256),
.Y(n_3432)
);

OR2x2_ASAP7_75t_L g3433 ( 
.A(n_3358),
.B(n_3379),
.Y(n_3433)
);

INVx3_ASAP7_75t_L g3434 ( 
.A(n_3401),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3352),
.Y(n_3435)
);

OR2x2_ASAP7_75t_L g3436 ( 
.A(n_3358),
.B(n_3159),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3354),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3355),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3330),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_3315),
.B(n_3155),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3357),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3382),
.B(n_3184),
.Y(n_3442)
);

OR2x2_ASAP7_75t_L g3443 ( 
.A(n_3379),
.B(n_3169),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3370),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3382),
.B(n_3332),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3373),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3374),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3380),
.Y(n_3448)
);

OR2x2_ASAP7_75t_L g3449 ( 
.A(n_3342),
.B(n_3295),
.Y(n_3449)
);

OR2x2_ASAP7_75t_L g3450 ( 
.A(n_3344),
.B(n_3196),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3332),
.B(n_3171),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_3335),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3372),
.B(n_3181),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3385),
.Y(n_3454)
);

OR2x2_ASAP7_75t_L g3455 ( 
.A(n_3367),
.B(n_3241),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3333),
.B(n_3249),
.Y(n_3456)
);

HB1xp67_ASAP7_75t_L g3457 ( 
.A(n_3377),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3319),
.B(n_3206),
.Y(n_3458)
);

INVxp33_ASAP7_75t_L g3459 ( 
.A(n_3376),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3389),
.Y(n_3460)
);

INVx1_ASAP7_75t_SL g3461 ( 
.A(n_3375),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3390),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_3372),
.B(n_3160),
.Y(n_3463)
);

OR2x2_ASAP7_75t_L g3464 ( 
.A(n_3367),
.B(n_3306),
.Y(n_3464)
);

OR2x2_ASAP7_75t_L g3465 ( 
.A(n_3323),
.B(n_3255),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3322),
.B(n_3165),
.Y(n_3466)
);

HB1xp67_ASAP7_75t_L g3467 ( 
.A(n_3400),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3324),
.B(n_3189),
.Y(n_3468)
);

INVx1_ASAP7_75t_SL g3469 ( 
.A(n_3359),
.Y(n_3469)
);

NOR2x1_ASAP7_75t_SL g3470 ( 
.A(n_3384),
.B(n_3205),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3324),
.B(n_3189),
.Y(n_3471)
);

INVx2_ASAP7_75t_SL g3472 ( 
.A(n_3384),
.Y(n_3472)
);

OR2x2_ASAP7_75t_L g3473 ( 
.A(n_3336),
.B(n_3282),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3366),
.Y(n_3474)
);

INVx3_ASAP7_75t_L g3475 ( 
.A(n_3337),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3457),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3457),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3467),
.Y(n_3478)
);

OR2x2_ASAP7_75t_L g3479 ( 
.A(n_3433),
.B(n_3328),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3467),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3436),
.Y(n_3481)
);

OAI221xp5_ASAP7_75t_L g3482 ( 
.A1(n_3428),
.A2(n_3145),
.B1(n_3293),
.B2(n_3329),
.C(n_3205),
.Y(n_3482)
);

AOI221xp5_ASAP7_75t_L g3483 ( 
.A1(n_3417),
.A2(n_3329),
.B1(n_3362),
.B2(n_3339),
.C(n_3327),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_L g3484 ( 
.A(n_3424),
.B(n_3040),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3440),
.B(n_3337),
.Y(n_3485)
);

OR2x2_ASAP7_75t_L g3486 ( 
.A(n_3408),
.B(n_3328),
.Y(n_3486)
);

OAI22xp33_ASAP7_75t_L g3487 ( 
.A1(n_3422),
.A2(n_3266),
.B1(n_3147),
.B2(n_3246),
.Y(n_3487)
);

INVx3_ASAP7_75t_L g3488 ( 
.A(n_3404),
.Y(n_3488)
);

A2O1A1Ixp33_ASAP7_75t_L g3489 ( 
.A1(n_3407),
.A2(n_3253),
.B(n_3279),
.C(n_3200),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3475),
.B(n_3337),
.Y(n_3490)
);

AOI22xp5_ASAP7_75t_L g3491 ( 
.A1(n_3417),
.A2(n_3362),
.B1(n_3341),
.B2(n_3353),
.Y(n_3491)
);

INVx1_ASAP7_75t_SL g3492 ( 
.A(n_3469),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3411),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3408),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3420),
.Y(n_3495)
);

OAI22xp33_ASAP7_75t_L g3496 ( 
.A1(n_3422),
.A2(n_3266),
.B1(n_3199),
.B2(n_3074),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3420),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3468),
.B(n_3340),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3475),
.B(n_3341),
.Y(n_3499)
);

OAI22xp33_ASAP7_75t_SL g3500 ( 
.A1(n_3461),
.A2(n_3074),
.B1(n_3110),
.B2(n_3094),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3456),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3456),
.Y(n_3502)
);

BUFx3_ASAP7_75t_L g3503 ( 
.A(n_3404),
.Y(n_3503)
);

AND2x4_ASAP7_75t_L g3504 ( 
.A(n_3423),
.B(n_3350),
.Y(n_3504)
);

OAI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3407),
.A2(n_2945),
.B(n_3308),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3455),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3445),
.B(n_3350),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3432),
.B(n_3353),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3464),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3403),
.Y(n_3510)
);

HB1xp67_ASAP7_75t_L g3511 ( 
.A(n_3411),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3406),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3410),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3413),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3419),
.Y(n_3515)
);

OR2x2_ASAP7_75t_L g3516 ( 
.A(n_3473),
.B(n_3361),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3421),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3451),
.B(n_3405),
.Y(n_3518)
);

OAI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_3459),
.A2(n_3265),
.B1(n_3267),
.B2(n_3366),
.Y(n_3519)
);

AOI22xp5_ASAP7_75t_L g3520 ( 
.A1(n_3412),
.A2(n_3364),
.B1(n_3363),
.B2(n_3383),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3414),
.Y(n_3521)
);

NAND3xp33_ASAP7_75t_L g3522 ( 
.A(n_3412),
.B(n_3310),
.C(n_3038),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3414),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3416),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3426),
.Y(n_3525)
);

INVx2_ASAP7_75t_SL g3526 ( 
.A(n_3434),
.Y(n_3526)
);

AOI32xp33_ASAP7_75t_L g3527 ( 
.A1(n_3459),
.A2(n_3458),
.A3(n_3434),
.B1(n_3425),
.B2(n_3472),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3468),
.B(n_3471),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3416),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3471),
.B(n_3340),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3418),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3418),
.Y(n_3532)
);

OAI211xp5_ASAP7_75t_L g3533 ( 
.A1(n_3458),
.A2(n_3110),
.B(n_3094),
.C(n_3040),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3430),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3427),
.Y(n_3535)
);

AND2x2_ASAP7_75t_L g3536 ( 
.A(n_3466),
.B(n_3363),
.Y(n_3536)
);

AOI22xp5_ASAP7_75t_L g3537 ( 
.A1(n_3409),
.A2(n_3364),
.B1(n_3386),
.B2(n_3383),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3429),
.B(n_3368),
.Y(n_3538)
);

INVx1_ASAP7_75t_SL g3539 ( 
.A(n_3450),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3504),
.B(n_3490),
.Y(n_3540)
);

AND2x2_ASAP7_75t_SL g3541 ( 
.A(n_3483),
.B(n_3470),
.Y(n_3541)
);

OAI211xp5_ASAP7_75t_SL g3542 ( 
.A1(n_3483),
.A2(n_3435),
.B(n_3438),
.C(n_3437),
.Y(n_3542)
);

OAI22xp33_ASAP7_75t_L g3543 ( 
.A1(n_3491),
.A2(n_3415),
.B1(n_3443),
.B2(n_3266),
.Y(n_3543)
);

OR2x2_ASAP7_75t_L g3544 ( 
.A(n_3498),
.B(n_3465),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3476),
.B(n_3361),
.Y(n_3545)
);

AOI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3522),
.A2(n_3463),
.B1(n_3386),
.B2(n_3356),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3477),
.Y(n_3547)
);

NOR3xp33_ASAP7_75t_L g3548 ( 
.A(n_3482),
.B(n_3304),
.C(n_3065),
.Y(n_3548)
);

INVxp67_ASAP7_75t_SL g3549 ( 
.A(n_3500),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3511),
.Y(n_3550)
);

AND2x4_ASAP7_75t_L g3551 ( 
.A(n_3504),
.B(n_3201),
.Y(n_3551)
);

AOI22xp5_ASAP7_75t_L g3552 ( 
.A1(n_3522),
.A2(n_3356),
.B1(n_3371),
.B2(n_3368),
.Y(n_3552)
);

AOI221xp5_ASAP7_75t_L g3553 ( 
.A1(n_3482),
.A2(n_3446),
.B1(n_3447),
.B2(n_3444),
.C(n_3441),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3495),
.Y(n_3554)
);

OAI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3489),
.A2(n_2999),
.B(n_3289),
.Y(n_3555)
);

O2A1O1Ixp33_ASAP7_75t_SL g3556 ( 
.A1(n_3487),
.A2(n_3496),
.B(n_3533),
.C(n_3492),
.Y(n_3556)
);

OAI31xp33_ASAP7_75t_SL g3557 ( 
.A1(n_3533),
.A2(n_3402),
.A3(n_3431),
.B(n_3442),
.Y(n_3557)
);

OAI22xp5_ASAP7_75t_L g3558 ( 
.A1(n_3520),
.A2(n_3449),
.B1(n_3474),
.B2(n_3453),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3497),
.Y(n_3559)
);

AOI21xp33_ASAP7_75t_L g3560 ( 
.A1(n_3487),
.A2(n_3107),
.B(n_3273),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3511),
.Y(n_3561)
);

NAND2xp33_ASAP7_75t_L g3562 ( 
.A(n_3527),
.B(n_2823),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3510),
.Y(n_3563)
);

OAI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3519),
.A2(n_3166),
.B1(n_3371),
.B2(n_3391),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3512),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3513),
.Y(n_3566)
);

OAI22xp33_ASAP7_75t_L g3567 ( 
.A1(n_3519),
.A2(n_3199),
.B1(n_3378),
.B2(n_3228),
.Y(n_3567)
);

OAI21xp33_ASAP7_75t_L g3568 ( 
.A1(n_3537),
.A2(n_3454),
.B(n_3448),
.Y(n_3568)
);

AOI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3505),
.A2(n_3248),
.B(n_2908),
.Y(n_3569)
);

NAND4xp25_ASAP7_75t_SL g3570 ( 
.A(n_3492),
.B(n_3244),
.C(n_3225),
.D(n_3069),
.Y(n_3570)
);

OAI22xp5_ASAP7_75t_L g3571 ( 
.A1(n_3488),
.A2(n_3336),
.B1(n_3462),
.B2(n_3460),
.Y(n_3571)
);

AOI22xp5_ASAP7_75t_L g3572 ( 
.A1(n_3501),
.A2(n_3381),
.B1(n_3244),
.B2(n_3322),
.Y(n_3572)
);

AOI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3502),
.A2(n_3381),
.B1(n_3188),
.B2(n_3190),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_R g3574 ( 
.A(n_3484),
.B(n_3069),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_3505),
.A2(n_2908),
.B(n_2993),
.Y(n_3575)
);

AOI33xp33_ASAP7_75t_L g3576 ( 
.A1(n_3539),
.A2(n_3481),
.A3(n_3509),
.B1(n_3506),
.B2(n_3494),
.B3(n_3514),
.Y(n_3576)
);

NAND3xp33_ASAP7_75t_L g3577 ( 
.A(n_3478),
.B(n_3393),
.C(n_3392),
.Y(n_3577)
);

AOI32xp33_ASAP7_75t_L g3578 ( 
.A1(n_3539),
.A2(n_3127),
.A3(n_3187),
.B1(n_3207),
.B2(n_3191),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_3488),
.A2(n_2989),
.B1(n_3296),
.B2(n_3059),
.Y(n_3579)
);

OAI22xp5_ASAP7_75t_L g3580 ( 
.A1(n_3503),
.A2(n_2989),
.B1(n_3059),
.B2(n_3243),
.Y(n_3580)
);

AOI21xp33_ASAP7_75t_L g3581 ( 
.A1(n_3480),
.A2(n_3152),
.B(n_3148),
.Y(n_3581)
);

OAI21xp33_ASAP7_75t_L g3582 ( 
.A1(n_3557),
.A2(n_3528),
.B(n_3526),
.Y(n_3582)
);

INVx3_ASAP7_75t_L g3583 ( 
.A(n_3551),
.Y(n_3583)
);

AOI221xp5_ASAP7_75t_L g3584 ( 
.A1(n_3556),
.A2(n_3517),
.B1(n_3534),
.B2(n_3525),
.C(n_3515),
.Y(n_3584)
);

OAI22xp33_ASAP7_75t_SL g3585 ( 
.A1(n_3549),
.A2(n_3479),
.B1(n_3516),
.B2(n_3528),
.Y(n_3585)
);

OAI22xp5_ASAP7_75t_L g3586 ( 
.A1(n_3541),
.A2(n_3486),
.B1(n_3530),
.B2(n_3498),
.Y(n_3586)
);

AOI211xp5_ASAP7_75t_SL g3587 ( 
.A1(n_3562),
.A2(n_3034),
.B(n_3079),
.C(n_3046),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3546),
.B(n_3530),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_3540),
.B(n_3551),
.Y(n_3589)
);

NOR2xp33_ASAP7_75t_L g3590 ( 
.A(n_3568),
.B(n_3485),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3550),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3577),
.Y(n_3592)
);

NOR2xp33_ASAP7_75t_SL g3593 ( 
.A(n_3570),
.B(n_2375),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3577),
.Y(n_3594)
);

NAND4xp25_ASAP7_75t_L g3595 ( 
.A(n_3548),
.B(n_2983),
.C(n_2984),
.D(n_3098),
.Y(n_3595)
);

OAI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_3553),
.A2(n_3518),
.B(n_3079),
.Y(n_3596)
);

NOR4xp25_ASAP7_75t_SL g3597 ( 
.A(n_3542),
.B(n_2823),
.C(n_3396),
.D(n_3394),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3545),
.Y(n_3598)
);

AOI221xp5_ASAP7_75t_L g3599 ( 
.A1(n_3567),
.A2(n_3398),
.B1(n_3499),
.B2(n_3507),
.C(n_3536),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3576),
.B(n_3508),
.Y(n_3600)
);

NAND3xp33_ASAP7_75t_SL g3601 ( 
.A(n_3578),
.B(n_2925),
.C(n_3098),
.Y(n_3601)
);

OA22x2_ASAP7_75t_L g3602 ( 
.A1(n_3552),
.A2(n_3564),
.B1(n_3572),
.B2(n_3579),
.Y(n_3602)
);

AOI221x1_ASAP7_75t_L g3603 ( 
.A1(n_3560),
.A2(n_2930),
.B1(n_3101),
.B2(n_3100),
.C(n_3015),
.Y(n_3603)
);

AOI211xp5_ASAP7_75t_L g3604 ( 
.A1(n_3543),
.A2(n_3034),
.B(n_3115),
.C(n_3046),
.Y(n_3604)
);

XNOR2x2_ASAP7_75t_L g3605 ( 
.A(n_3575),
.B(n_3132),
.Y(n_3605)
);

AOI32xp33_ASAP7_75t_L g3606 ( 
.A1(n_3580),
.A2(n_3538),
.A3(n_3127),
.B1(n_3210),
.B2(n_2947),
.Y(n_3606)
);

AOI22xp5_ASAP7_75t_L g3607 ( 
.A1(n_3558),
.A2(n_3216),
.B1(n_3521),
.B2(n_3493),
.Y(n_3607)
);

NAND3xp33_ASAP7_75t_SL g3608 ( 
.A(n_3569),
.B(n_2925),
.C(n_3143),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3581),
.A2(n_3524),
.B(n_3523),
.Y(n_3609)
);

AOI221xp5_ASAP7_75t_L g3610 ( 
.A1(n_3571),
.A2(n_3529),
.B1(n_3535),
.B2(n_3532),
.C(n_3531),
.Y(n_3610)
);

AOI32xp33_ASAP7_75t_L g3611 ( 
.A1(n_3561),
.A2(n_3559),
.A3(n_3554),
.B1(n_3547),
.B2(n_3563),
.Y(n_3611)
);

OR2x2_ASAP7_75t_L g3612 ( 
.A(n_3544),
.B(n_3427),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3565),
.B(n_3439),
.Y(n_3613)
);

OAI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_3573),
.A2(n_3397),
.B1(n_2930),
.B2(n_3015),
.Y(n_3614)
);

OAI22xp33_ASAP7_75t_SL g3615 ( 
.A1(n_3555),
.A2(n_3300),
.B1(n_3298),
.B2(n_3194),
.Y(n_3615)
);

AOI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_3566),
.A2(n_3240),
.B1(n_3239),
.B2(n_3162),
.Y(n_3616)
);

XOR2x2_ASAP7_75t_L g3617 ( 
.A(n_3574),
.B(n_3260),
.Y(n_3617)
);

OAI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3541),
.A2(n_3143),
.B1(n_3164),
.B2(n_3439),
.Y(n_3618)
);

NAND3xp33_ASAP7_75t_SL g3619 ( 
.A(n_3548),
.B(n_3001),
.C(n_3131),
.Y(n_3619)
);

AOI222xp33_ASAP7_75t_L g3620 ( 
.A1(n_3541),
.A2(n_3115),
.B1(n_3039),
.B2(n_3387),
.C1(n_3212),
.C2(n_3229),
.Y(n_3620)
);

OAI21xp33_ASAP7_75t_L g3621 ( 
.A1(n_3557),
.A2(n_3387),
.B(n_3452),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_3541),
.A2(n_3001),
.B(n_3039),
.Y(n_3622)
);

OAI31xp33_ASAP7_75t_L g3623 ( 
.A1(n_3556),
.A2(n_3097),
.A3(n_2931),
.B(n_3108),
.Y(n_3623)
);

OAI21xp5_ASAP7_75t_SL g3624 ( 
.A1(n_3557),
.A2(n_3108),
.B(n_2940),
.Y(n_3624)
);

AOI21xp5_ASAP7_75t_SL g3625 ( 
.A1(n_3549),
.A2(n_2957),
.B(n_2935),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3550),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3598),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3592),
.B(n_3452),
.Y(n_3628)
);

OAI211xp5_ASAP7_75t_L g3629 ( 
.A1(n_3623),
.A2(n_3131),
.B(n_3099),
.C(n_2539),
.Y(n_3629)
);

AOI21xp5_ASAP7_75t_L g3630 ( 
.A1(n_3602),
.A2(n_3097),
.B(n_3208),
.Y(n_3630)
);

NAND2x1_ASAP7_75t_L g3631 ( 
.A(n_3583),
.B(n_3140),
.Y(n_3631)
);

OAI321xp33_ASAP7_75t_L g3632 ( 
.A1(n_3584),
.A2(n_3044),
.A3(n_3238),
.B1(n_3305),
.B2(n_2733),
.C(n_3050),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3613),
.Y(n_3633)
);

INVx2_ASAP7_75t_SL g3634 ( 
.A(n_3617),
.Y(n_3634)
);

NAND3xp33_ASAP7_75t_L g3635 ( 
.A(n_3620),
.B(n_2364),
.C(n_2356),
.Y(n_3635)
);

OAI211xp5_ASAP7_75t_L g3636 ( 
.A1(n_3625),
.A2(n_3619),
.B(n_3606),
.C(n_3587),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3593),
.A2(n_3197),
.B(n_3174),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3594),
.B(n_3226),
.Y(n_3638)
);

NAND3xp33_ASAP7_75t_SL g3639 ( 
.A(n_3597),
.B(n_2733),
.C(n_2669),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3588),
.B(n_3212),
.Y(n_3640)
);

NAND3xp33_ASAP7_75t_L g3641 ( 
.A(n_3611),
.B(n_2492),
.C(n_3050),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_SL g3642 ( 
.A1(n_3585),
.A2(n_3007),
.B1(n_3251),
.B2(n_3220),
.Y(n_3642)
);

INVxp67_ASAP7_75t_SL g3643 ( 
.A(n_3615),
.Y(n_3643)
);

NOR3xp33_ASAP7_75t_L g3644 ( 
.A(n_3608),
.B(n_2765),
.C(n_2757),
.Y(n_3644)
);

NAND3xp33_ASAP7_75t_L g3645 ( 
.A(n_3586),
.B(n_2606),
.C(n_2600),
.Y(n_3645)
);

AOI211x1_ASAP7_75t_L g3646 ( 
.A1(n_3582),
.A2(n_3214),
.B(n_3221),
.C(n_3213),
.Y(n_3646)
);

OAI21xp5_ASAP7_75t_SL g3647 ( 
.A1(n_3603),
.A2(n_2957),
.B(n_2935),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3612),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3591),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3626),
.Y(n_3650)
);

NAND2x1_ASAP7_75t_L g3651 ( 
.A(n_3583),
.B(n_3140),
.Y(n_3651)
);

NOR2x1_ASAP7_75t_L g3652 ( 
.A(n_3624),
.B(n_2431),
.Y(n_3652)
);

OAI21xp5_ASAP7_75t_SL g3653 ( 
.A1(n_3622),
.A2(n_2963),
.B(n_3078),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3600),
.B(n_3213),
.Y(n_3654)
);

AOI211x1_ASAP7_75t_L g3655 ( 
.A1(n_3596),
.A2(n_3221),
.B(n_3229),
.C(n_3214),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3589),
.B(n_3222),
.Y(n_3656)
);

AOI211xp5_ASAP7_75t_L g3657 ( 
.A1(n_3618),
.A2(n_2963),
.B(n_2958),
.C(n_3088),
.Y(n_3657)
);

NAND3xp33_ASAP7_75t_L g3658 ( 
.A(n_3636),
.B(n_3599),
.C(n_3595),
.Y(n_3658)
);

NOR3xp33_ASAP7_75t_L g3659 ( 
.A(n_3629),
.B(n_3601),
.C(n_3590),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3643),
.B(n_3621),
.Y(n_3660)
);

NAND3xp33_ASAP7_75t_L g3661 ( 
.A(n_3634),
.B(n_3604),
.C(n_3610),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3642),
.B(n_3607),
.Y(n_3662)
);

AND2x2_ASAP7_75t_L g3663 ( 
.A(n_3648),
.B(n_3616),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_3627),
.B(n_3609),
.Y(n_3664)
);

AOI21xp5_ASAP7_75t_L g3665 ( 
.A1(n_3630),
.A2(n_3614),
.B(n_3605),
.Y(n_3665)
);

NOR3xp33_ASAP7_75t_L g3666 ( 
.A(n_3632),
.B(n_2527),
.C(n_2378),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3656),
.B(n_3633),
.Y(n_3667)
);

NOR2x1_ASAP7_75t_L g3668 ( 
.A(n_3647),
.B(n_3631),
.Y(n_3668)
);

NOR3xp33_ASAP7_75t_L g3669 ( 
.A(n_3641),
.B(n_2338),
.C(n_2320),
.Y(n_3669)
);

NOR2x1_ASAP7_75t_L g3670 ( 
.A(n_3651),
.B(n_2431),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3654),
.B(n_3149),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3638),
.Y(n_3672)
);

NOR2x1_ASAP7_75t_L g3673 ( 
.A(n_3645),
.B(n_2448),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3649),
.Y(n_3674)
);

AOI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3637),
.A2(n_2898),
.B(n_3168),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3655),
.B(n_3149),
.Y(n_3676)
);

NOR3xp33_ASAP7_75t_L g3677 ( 
.A(n_3645),
.B(n_2765),
.C(n_2757),
.Y(n_3677)
);

NOR3x1_ASAP7_75t_L g3678 ( 
.A(n_3653),
.B(n_3635),
.C(n_3639),
.Y(n_3678)
);

NOR3xp33_ASAP7_75t_L g3679 ( 
.A(n_3652),
.B(n_2769),
.C(n_2512),
.Y(n_3679)
);

NAND3xp33_ASAP7_75t_L g3680 ( 
.A(n_3646),
.B(n_2492),
.C(n_2600),
.Y(n_3680)
);

OAI211xp5_ASAP7_75t_SL g3681 ( 
.A1(n_3644),
.A2(n_3142),
.B(n_2898),
.C(n_2769),
.Y(n_3681)
);

NOR3x1_ASAP7_75t_L g3682 ( 
.A(n_3628),
.B(n_2490),
.C(n_2512),
.Y(n_3682)
);

XOR2x2_ASAP7_75t_L g3683 ( 
.A(n_3661),
.B(n_3640),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3674),
.Y(n_3684)
);

NOR3xp33_ASAP7_75t_L g3685 ( 
.A(n_3658),
.B(n_3650),
.C(n_3657),
.Y(n_3685)
);

NAND4xp75_ASAP7_75t_L g3686 ( 
.A(n_3678),
.B(n_3668),
.C(n_3660),
.D(n_3665),
.Y(n_3686)
);

NAND3xp33_ASAP7_75t_L g3687 ( 
.A(n_3659),
.B(n_2606),
.C(n_2600),
.Y(n_3687)
);

AOI22xp5_ASAP7_75t_L g3688 ( 
.A1(n_3664),
.A2(n_3007),
.B1(n_2448),
.B2(n_2454),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3667),
.Y(n_3689)
);

NOR2x1_ASAP7_75t_SL g3690 ( 
.A(n_3672),
.B(n_2452),
.Y(n_3690)
);

AOI21xp33_ASAP7_75t_SL g3691 ( 
.A1(n_3662),
.A2(n_2459),
.B(n_2454),
.Y(n_3691)
);

NAND4xp75_ASAP7_75t_L g3692 ( 
.A(n_3673),
.B(n_2523),
.C(n_2340),
.D(n_2619),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3663),
.Y(n_3693)
);

NAND3xp33_ASAP7_75t_L g3694 ( 
.A(n_3679),
.B(n_2606),
.C(n_2600),
.Y(n_3694)
);

NAND3xp33_ASAP7_75t_L g3695 ( 
.A(n_3669),
.B(n_2606),
.C(n_2618),
.Y(n_3695)
);

NAND3xp33_ASAP7_75t_SL g3696 ( 
.A(n_3666),
.B(n_2669),
.C(n_2615),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3676),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3675),
.B(n_3150),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3671),
.B(n_3150),
.Y(n_3699)
);

NOR2xp33_ASAP7_75t_L g3700 ( 
.A(n_3671),
.B(n_3153),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3670),
.Y(n_3701)
);

NAND3xp33_ASAP7_75t_SL g3702 ( 
.A(n_3677),
.B(n_2849),
.C(n_3275),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3682),
.Y(n_3703)
);

NOR3xp33_ASAP7_75t_L g3704 ( 
.A(n_3681),
.B(n_2520),
.C(n_2464),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3684),
.Y(n_3705)
);

OAI211xp5_ASAP7_75t_L g3706 ( 
.A1(n_3685),
.A2(n_3680),
.B(n_3142),
.C(n_2445),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3689),
.Y(n_3707)
);

INVxp67_ASAP7_75t_L g3708 ( 
.A(n_3686),
.Y(n_3708)
);

NOR2xp67_ASAP7_75t_L g3709 ( 
.A(n_3703),
.B(n_3021),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3690),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3701),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3693),
.Y(n_3712)
);

INVx2_ASAP7_75t_SL g3713 ( 
.A(n_3683),
.Y(n_3713)
);

NOR2x1_ASAP7_75t_L g3714 ( 
.A(n_3696),
.B(n_3687),
.Y(n_3714)
);

NOR2x1_ASAP7_75t_L g3715 ( 
.A(n_3697),
.B(n_2308),
.Y(n_3715)
);

NAND2x1p5_ASAP7_75t_L g3716 ( 
.A(n_3698),
.B(n_3045),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3699),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3700),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3708),
.B(n_3713),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3711),
.A2(n_3712),
.B(n_3705),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3712),
.Y(n_3721)
);

CKINVDCx20_ASAP7_75t_R g3722 ( 
.A(n_3707),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3716),
.Y(n_3723)
);

AOI22xp5_ASAP7_75t_L g3724 ( 
.A1(n_3709),
.A2(n_3702),
.B1(n_3704),
.B2(n_3688),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3717),
.Y(n_3725)
);

OAI22xp5_ASAP7_75t_L g3726 ( 
.A1(n_3714),
.A2(n_3691),
.B1(n_3688),
.B2(n_3694),
.Y(n_3726)
);

INVx1_ASAP7_75t_SL g3727 ( 
.A(n_3710),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3717),
.Y(n_3728)
);

OR2x2_ASAP7_75t_L g3729 ( 
.A(n_3718),
.B(n_3695),
.Y(n_3729)
);

AO21x1_ASAP7_75t_L g3730 ( 
.A1(n_3719),
.A2(n_3706),
.B(n_3715),
.Y(n_3730)
);

OAI22xp5_ASAP7_75t_L g3731 ( 
.A1(n_3727),
.A2(n_3692),
.B1(n_3021),
.B2(n_3120),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3723),
.Y(n_3732)
);

OAI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_3720),
.A2(n_2490),
.B(n_2465),
.Y(n_3733)
);

OAI21xp5_ASAP7_75t_SL g3734 ( 
.A1(n_3729),
.A2(n_3120),
.B(n_3103),
.Y(n_3734)
);

CKINVDCx5p33_ASAP7_75t_R g3735 ( 
.A(n_3722),
.Y(n_3735)
);

OAI22xp5_ASAP7_75t_L g3736 ( 
.A1(n_3724),
.A2(n_3103),
.B1(n_3081),
.B2(n_3045),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3732),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3735),
.Y(n_3738)
);

AOI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_3730),
.A2(n_3726),
.B1(n_3728),
.B2(n_3725),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3736),
.Y(n_3740)
);

INVx3_ASAP7_75t_L g3741 ( 
.A(n_3734),
.Y(n_3741)
);

OA22x2_ASAP7_75t_L g3742 ( 
.A1(n_3737),
.A2(n_3721),
.B1(n_3731),
.B2(n_3733),
.Y(n_3742)
);

OAI22xp5_ASAP7_75t_L g3743 ( 
.A1(n_3738),
.A2(n_3092),
.B1(n_3081),
.B2(n_3153),
.Y(n_3743)
);

OAI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3742),
.A2(n_3739),
.B(n_3740),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3743),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3744),
.A2(n_3741),
.B(n_2464),
.Y(n_3746)
);

OR2x6_ASAP7_75t_L g3747 ( 
.A(n_3746),
.B(n_3745),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3747),
.Y(n_3748)
);

AOI22xp33_ASAP7_75t_L g3749 ( 
.A1(n_3748),
.A2(n_3092),
.B1(n_2459),
.B2(n_2308),
.Y(n_3749)
);


endmodule