module fake_netlist_1_7861_n_30 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_30);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_0), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_0), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
A2O1A1Ixp33_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_1), .B(n_2), .C(n_3), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
AND2x6_ASAP7_75t_L g18 ( .A(n_15), .B(n_7), .Y(n_18) );
CKINVDCx14_ASAP7_75t_R g19 ( .A(n_11), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_16), .B(n_14), .C(n_13), .Y(n_20) );
INVx5_ASAP7_75t_SL g21 ( .A(n_19), .Y(n_21) );
AND2x4_ASAP7_75t_L g22 ( .A(n_20), .B(n_17), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_15), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_25), .Y(n_26) );
XOR2xp5_ASAP7_75t_L g27 ( .A(n_25), .B(n_22), .Y(n_27) );
AO22x2_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_22), .B1(n_23), .B2(n_6), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_26), .B(n_22), .Y(n_29) );
AOI222xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_3), .B1(n_5), .B2(n_8), .C1(n_18), .C2(n_29), .Y(n_30) );
endmodule