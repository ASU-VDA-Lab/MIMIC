module fake_jpeg_17420_n_111 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_27),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_33),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_30),
.B1(n_37),
.B2(n_15),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_11),
.B1(n_20),
.B2(n_17),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_19),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_18),
.C(n_27),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_21),
.A2(n_0),
.B1(n_18),
.B2(n_2),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_45),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_23),
.B1(n_27),
.B2(n_18),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_34),
.B1(n_35),
.B2(n_31),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_10),
.B(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_46),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_37),
.B1(n_13),
.B2(n_12),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_0),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_61),
.B1(n_29),
.B2(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_13),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_42),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_44),
.B(n_47),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2x1_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_45),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_69),
.B(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_39),
.B1(n_35),
.B2(n_12),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_71),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_39),
.B(n_0),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_57),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_73),
.Y(n_88)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_56),
.B(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_57),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_80),
.C(n_83),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_60),
.C(n_54),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_51),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_83),
.C(n_67),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_87),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_82),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_69),
.B(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_88),
.B(n_78),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_58),
.C(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_90),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_64),
.C(n_68),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_63),
.B(n_61),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_3),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_96),
.B(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_101),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_94),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_4),
.B(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_5),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_107),
.B(n_103),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_7),
.B(n_9),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_110),
.Y(n_111)
);


endmodule