module fake_netlist_1_6275_n_957 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_957);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_957;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_949;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_951;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_947;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g233 ( .A(n_172), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_98), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_44), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_185), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_82), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_133), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_212), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_178), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_189), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_183), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_13), .Y(n_243) );
BUFx10_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_121), .Y(n_245) );
INVx1_ASAP7_75t_SL g246 ( .A(n_53), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_139), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_166), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_107), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_145), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_102), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_3), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_59), .Y(n_253) );
INVxp67_ASAP7_75t_L g254 ( .A(n_206), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_42), .Y(n_255) );
CKINVDCx14_ASAP7_75t_R g256 ( .A(n_12), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_12), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_138), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_215), .Y(n_259) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_83), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_186), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_163), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_52), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_130), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_149), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_170), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_77), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_79), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_56), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_94), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_112), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_37), .Y(n_272) );
INVxp33_ASAP7_75t_L g273 ( .A(n_86), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_177), .Y(n_274) );
CKINVDCx14_ASAP7_75t_R g275 ( .A(n_131), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_74), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_53), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_39), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_16), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_75), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_86), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_187), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_62), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_60), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_64), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_64), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_34), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_188), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_208), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_191), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_157), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_201), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_132), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_228), .Y(n_294) );
BUFx10_ASAP7_75t_L g295 ( .A(n_26), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_95), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_125), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_49), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_171), .Y(n_299) );
INVxp67_ASAP7_75t_SL g300 ( .A(n_42), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_74), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_128), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_14), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_104), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_114), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_147), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_15), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_18), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_20), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_221), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_36), .Y(n_311) );
CKINVDCx16_ASAP7_75t_R g312 ( .A(n_110), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_46), .Y(n_313) );
INVxp33_ASAP7_75t_L g314 ( .A(n_174), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_205), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_158), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_127), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_90), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_24), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_118), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_150), .Y(n_321) );
BUFx10_ASAP7_75t_L g322 ( .A(n_154), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_79), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_0), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_85), .Y(n_325) );
CKINVDCx14_ASAP7_75t_R g326 ( .A(n_109), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_200), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_84), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_78), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_176), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_126), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_28), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_160), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_162), .Y(n_334) );
BUFx10_ASAP7_75t_L g335 ( .A(n_224), .Y(n_335) );
INVxp33_ASAP7_75t_L g336 ( .A(n_60), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_54), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_140), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_231), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_59), .B(n_153), .Y(n_340) );
BUFx3_ASAP7_75t_L g341 ( .A(n_75), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_198), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_81), .Y(n_343) );
INVxp67_ASAP7_75t_L g344 ( .A(n_227), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_124), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_129), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_167), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_5), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_103), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_57), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_41), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_192), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_211), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_29), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_43), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_93), .Y(n_356) );
INVxp33_ASAP7_75t_SL g357 ( .A(n_58), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_4), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_182), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_108), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_66), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_117), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_70), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_175), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_20), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_268), .B(n_0), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_268), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_273), .B(n_1), .Y(n_368) );
AND2x6_ASAP7_75t_L g369 ( .A(n_291), .B(n_96), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_256), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_256), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_265), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_341), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_265), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_271), .B(n_2), .Y(n_375) );
INVx4_ASAP7_75t_L g376 ( .A(n_244), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_234), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_238), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_311), .Y(n_379) );
CKINVDCx6p67_ASAP7_75t_R g380 ( .A(n_261), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_239), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_252), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_240), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_241), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_237), .B(n_6), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_265), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_245), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_293), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g389 ( .A1(n_263), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_282), .B(n_7), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_273), .B(n_8), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_336), .B(n_10), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_293), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_336), .B(n_10), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_291), .B(n_11), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_247), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_248), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_233), .B(n_11), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_317), .B(n_14), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_250), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_244), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_293), .Y(n_402) );
BUFx12f_ASAP7_75t_L g403 ( .A(n_244), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_376), .B(n_312), .Y(n_404) );
INVx4_ASAP7_75t_L g405 ( .A(n_395), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_366), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
INVx3_ASAP7_75t_L g408 ( .A(n_366), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_371), .B(n_233), .Y(n_409) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_382), .B(n_260), .C(n_286), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_376), .Y(n_411) );
XNOR2xp5_ASAP7_75t_L g412 ( .A(n_371), .B(n_263), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_386), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_370), .A2(n_323), .B1(n_324), .B2(n_303), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_395), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_386), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_386), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_377), .B(n_314), .Y(n_419) );
AOI22xp5_ASAP7_75t_SL g420 ( .A1(n_382), .A2(n_323), .B1(n_324), .B2(n_303), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
BUFx4f_ASAP7_75t_L g422 ( .A(n_369), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_386), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_376), .B(n_314), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_377), .B(n_236), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_395), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_399), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_401), .B(n_254), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_399), .Y(n_430) );
INVx5_ASAP7_75t_L g431 ( .A(n_369), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_399), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_368), .A2(n_257), .B1(n_270), .B2(n_235), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_401), .B(n_351), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_386), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_401), .B(n_339), .Y(n_437) );
NAND2xp33_ASAP7_75t_L g438 ( .A(n_369), .B(n_242), .Y(n_438) );
BUFx4f_ASAP7_75t_L g439 ( .A(n_369), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_401), .B(n_351), .Y(n_440) );
BUFx4f_ASAP7_75t_L g441 ( .A(n_369), .Y(n_441) );
INVx4_ASAP7_75t_L g442 ( .A(n_369), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_372), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_403), .B(n_322), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_378), .B(n_236), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g446 ( .A1(n_370), .A2(n_283), .B1(n_287), .B2(n_255), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_378), .B(n_258), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_372), .Y(n_448) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_368), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_422), .Y(n_450) );
AND2x6_ASAP7_75t_SL g451 ( .A(n_420), .B(n_392), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_405), .B(n_398), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_409), .B(n_403), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_443), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_449), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_425), .B(n_391), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_419), .B(n_379), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_405), .A2(n_375), .B1(n_390), .B2(n_383), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_409), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_411), .B(n_403), .Y(n_460) );
NOR2x2_ASAP7_75t_L g461 ( .A(n_412), .B(n_380), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_412), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_435), .B(n_380), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_422), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_406), .Y(n_465) );
NOR2x2_ASAP7_75t_L g466 ( .A(n_420), .B(n_325), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_405), .A2(n_375), .B1(n_390), .B2(n_383), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_422), .A2(n_390), .B(n_375), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_440), .B(n_381), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_429), .B(n_381), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_443), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_442), .B(n_375), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_437), .B(n_384), .Y(n_473) );
AND2x4_ASAP7_75t_SL g474 ( .A(n_410), .B(n_306), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_448), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_406), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_404), .B(n_390), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_407), .B(n_384), .Y(n_478) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_422), .B(n_392), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_408), .A2(n_387), .B1(n_397), .B2(n_396), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_415), .B(n_394), .Y(n_482) );
INVx3_ASAP7_75t_L g483 ( .A(n_408), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_442), .B(n_397), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_413), .B(n_400), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_413), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_416), .B(n_400), .Y(n_487) );
BUFx2_ASAP7_75t_L g488 ( .A(n_415), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_416), .B(n_385), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_446), .A2(n_357), .B1(n_316), .B2(n_331), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_434), .A2(n_316), .B1(n_331), .B2(n_306), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_421), .B(n_367), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_408), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_421), .B(n_367), .Y(n_495) );
INVx5_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
NOR2x2_ASAP7_75t_L g497 ( .A(n_444), .B(n_325), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_441), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_427), .A2(n_253), .B1(n_269), .B2(n_243), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_433), .A2(n_373), .B1(n_369), .B2(n_326), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_427), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_441), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_428), .B(n_249), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_428), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_433), .A2(n_369), .B1(n_326), .B2(n_275), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_430), .B(n_300), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_430), .A2(n_275), .B1(n_277), .B2(n_276), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_432), .B(n_352), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_441), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_432), .B(n_352), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_426), .Y(n_511) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_426), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_445), .A2(n_279), .B1(n_280), .B2(n_278), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_445), .B(n_295), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_447), .A2(n_284), .B1(n_285), .B2(n_281), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_438), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_441), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_431), .A2(n_308), .B1(n_309), .B2(n_307), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_414), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_414), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_414), .Y(n_521) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_431), .B(n_313), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_431), .Y(n_523) );
NOR2x2_ASAP7_75t_L g524 ( .A(n_417), .B(n_332), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_418), .B(n_318), .Y(n_525) );
OR2x6_ASAP7_75t_L g526 ( .A(n_418), .B(n_319), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_418), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_423), .B(n_251), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_436), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_512), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_511), .Y(n_531) );
BUFx8_ASAP7_75t_L g532 ( .A(n_488), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_514), .B(n_389), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_SL g534 ( .A1(n_453), .A2(n_340), .B(n_374), .C(n_372), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_472), .A2(n_424), .B(n_423), .Y(n_535) );
NOR3xp33_ASAP7_75t_SL g536 ( .A(n_462), .B(n_492), .C(n_301), .Y(n_536) );
NOR2xp33_ASAP7_75t_R g537 ( .A(n_462), .B(n_332), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_459), .B(n_343), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_524), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_458), .A2(n_467), .B1(n_485), .B2(n_478), .Y(n_540) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_450), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_457), .B(n_343), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_456), .A2(n_329), .B(n_337), .C(n_328), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_455), .B(n_355), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_482), .B(n_295), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_483), .Y(n_546) );
INVx4_ASAP7_75t_L g547 ( .A(n_452), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_482), .A2(n_298), .B1(n_348), .B2(n_246), .Y(n_549) );
BUFx2_ASAP7_75t_L g550 ( .A(n_524), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_494), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_487), .A2(n_354), .B1(n_356), .B2(n_350), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_494), .Y(n_553) );
INVx5_ASAP7_75t_L g554 ( .A(n_526), .Y(n_554) );
NOR2x1_ASAP7_75t_L g555 ( .A(n_463), .B(n_358), .Y(n_555) );
INVx3_ASAP7_75t_SL g556 ( .A(n_461), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_465), .A2(n_363), .B1(n_361), .B2(n_259), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_474), .B(n_295), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g559 ( .A1(n_466), .A2(n_365), .B1(n_344), .B2(n_292), .Y(n_559) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_450), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_476), .A2(n_262), .B1(n_266), .B2(n_264), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_474), .A2(n_335), .B1(n_322), .B2(n_267), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_464), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_496), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_496), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_496), .Y(n_566) );
INVx3_ASAP7_75t_L g567 ( .A(n_496), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_493), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_464), .Y(n_569) );
INVxp67_ASAP7_75t_SL g570 ( .A(n_517), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_486), .A2(n_504), .B1(n_501), .B2(n_489), .Y(n_571) );
NOR2xp33_ASAP7_75t_R g572 ( .A(n_451), .B(n_322), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_469), .A2(n_289), .B1(n_290), .B2(n_288), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_526), .Y(n_574) );
INVx4_ASAP7_75t_L g575 ( .A(n_526), .Y(n_575) );
A2O1A1Ixp33_ASAP7_75t_L g576 ( .A1(n_468), .A2(n_294), .B(n_299), .C(n_297), .Y(n_576) );
O2A1O1Ixp5_ASAP7_75t_L g577 ( .A1(n_470), .A2(n_302), .B(n_310), .C(n_258), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_481), .B(n_304), .Y(n_578) );
BUFx2_ASAP7_75t_L g579 ( .A(n_466), .Y(n_579) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_517), .Y(n_580) );
INVx4_ASAP7_75t_L g581 ( .A(n_526), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_454), .Y(n_582) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_480), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_506), .B(n_335), .Y(n_584) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_480), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_473), .A2(n_320), .B1(n_333), .B2(n_315), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_L g587 ( .A1(n_495), .A2(n_338), .B(n_345), .C(n_334), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_477), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_513), .A2(n_347), .B1(n_349), .B2(n_346), .Y(n_589) );
NOR2xp33_ASAP7_75t_SL g590 ( .A(n_502), .B(n_305), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_477), .B(n_360), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_460), .B(n_364), .Y(n_592) );
BUFx2_ASAP7_75t_L g593 ( .A(n_497), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_516), .A2(n_353), .B(n_310), .C(n_330), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_471), .Y(n_595) );
NAND3xp33_ASAP7_75t_SL g596 ( .A(n_507), .B(n_274), .C(n_321), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_499), .B(n_267), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_503), .B(n_327), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_479), .A2(n_342), .B1(n_272), .B2(n_267), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_508), .B(n_510), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_484), .A2(n_353), .B(n_330), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_515), .A2(n_272), .B1(n_267), .B2(n_317), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_475), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_497), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_525), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_479), .B(n_272), .Y(n_606) );
BUFx3_ASAP7_75t_L g607 ( .A(n_525), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_528), .A2(n_388), .B(n_436), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_522), .Y(n_609) );
BUFx2_ASAP7_75t_L g610 ( .A(n_525), .Y(n_610) );
NOR2xp33_ASAP7_75t_R g611 ( .A(n_505), .B(n_15), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_500), .B(n_16), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_518), .A2(n_296), .B1(n_359), .B2(n_293), .Y(n_613) );
AND2x6_ASAP7_75t_L g614 ( .A(n_498), .B(n_296), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_490), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_519), .A2(n_436), .B(n_362), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_490), .B(n_17), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_490), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_509), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_527), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_527), .B(n_18), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_519), .A2(n_436), .B(n_362), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_520), .A2(n_362), .B(n_359), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_523), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_509), .B(n_19), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_520), .A2(n_362), .B(n_402), .C(n_393), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_509), .A2(n_402), .B1(n_393), .B2(n_22), .Y(n_627) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_521), .B(n_19), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_529), .B(n_21), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_529), .B(n_393), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_529), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_472), .A2(n_402), .B(n_393), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_511), .A2(n_402), .B1(n_393), .B2(n_23), .Y(n_633) );
BUFx3_ASAP7_75t_L g634 ( .A(n_514), .Y(n_634) );
AOI21x1_ASAP7_75t_L g635 ( .A1(n_472), .A2(n_99), .B(n_97), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_496), .Y(n_636) );
BUFx12f_ASAP7_75t_L g637 ( .A(n_451), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_472), .A2(n_101), .B(n_100), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_531), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_530), .B(n_21), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_595), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_571), .A2(n_608), .B(n_535), .Y(n_642) );
AO31x2_ASAP7_75t_L g643 ( .A1(n_571), .A2(n_24), .A3(n_22), .B(n_23), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_542), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_644) );
BUFx3_ASAP7_75t_L g645 ( .A(n_609), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_533), .B(n_29), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_634), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_545), .B(n_30), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_568), .A2(n_543), .B(n_606), .C(n_577), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_603), .Y(n_650) );
AOI221xp5_ASAP7_75t_SL g651 ( .A1(n_576), .A2(n_31), .B1(n_32), .B2(n_33), .C(n_34), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_574), .A2(n_33), .B1(n_35), .B2(n_36), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_538), .B(n_35), .Y(n_653) );
INVx3_ASAP7_75t_L g654 ( .A(n_547), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_603), .Y(n_655) );
BUFx3_ASAP7_75t_L g656 ( .A(n_556), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_540), .A2(n_106), .B(n_105), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_536), .B(n_38), .C(n_40), .Y(n_658) );
AO31x2_ASAP7_75t_L g659 ( .A1(n_633), .A2(n_44), .A3(n_45), .B(n_46), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_582), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_539), .A2(n_47), .B1(n_48), .B2(n_49), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_588), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_574), .A2(n_50), .B1(n_51), .B2(n_52), .Y(n_663) );
BUFx12f_ASAP7_75t_L g664 ( .A(n_579), .Y(n_664) );
CKINVDCx6p67_ASAP7_75t_R g665 ( .A(n_554), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_550), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_532), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_667) );
AO32x2_ASAP7_75t_L g668 ( .A1(n_602), .A2(n_561), .A3(n_573), .B1(n_586), .B2(n_613), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_544), .Y(n_669) );
INVx8_ASAP7_75t_L g670 ( .A(n_554), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_558), .B(n_61), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_591), .Y(n_672) );
BUFx2_ASAP7_75t_L g673 ( .A(n_537), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_597), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_554), .A2(n_63), .B1(n_65), .B2(n_66), .Y(n_675) );
NAND2x1p5_ASAP7_75t_L g676 ( .A(n_575), .B(n_67), .Y(n_676) );
AO31x2_ASAP7_75t_L g677 ( .A1(n_594), .A2(n_68), .A3(n_69), .B(n_70), .Y(n_677) );
AO32x2_ASAP7_75t_L g678 ( .A1(n_602), .A2(n_68), .A3(n_69), .B1(n_71), .B2(n_72), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_632), .A2(n_113), .B(n_111), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_549), .B(n_71), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_559), .A2(n_73), .B1(n_76), .B2(n_77), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_572), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_575), .A2(n_581), .B1(n_610), .B2(n_605), .Y(n_683) );
AO32x2_ASAP7_75t_L g684 ( .A1(n_561), .A2(n_78), .A3(n_80), .B1(n_81), .B2(n_82), .Y(n_684) );
BUFx3_ASAP7_75t_L g685 ( .A(n_637), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_621), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_555), .B(n_84), .Y(n_687) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_541), .Y(n_688) );
AO31x2_ASAP7_75t_L g689 ( .A1(n_626), .A2(n_85), .A3(n_87), .B(n_88), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_584), .Y(n_690) );
AO31x2_ASAP7_75t_L g691 ( .A1(n_613), .A2(n_629), .A3(n_573), .B(n_586), .Y(n_691) );
BUFx2_ASAP7_75t_L g692 ( .A(n_570), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_578), .Y(n_693) );
AO21x2_ASAP7_75t_L g694 ( .A1(n_534), .A2(n_156), .B(n_230), .Y(n_694) );
OAI21xp5_ASAP7_75t_L g695 ( .A1(n_601), .A2(n_155), .B(n_229), .Y(n_695) );
AO32x2_ASAP7_75t_L g696 ( .A1(n_557), .A2(n_88), .A3(n_89), .B1(n_90), .B2(n_91), .Y(n_696) );
OAI21x1_ASAP7_75t_L g697 ( .A1(n_630), .A2(n_159), .B(n_226), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_532), .A2(n_91), .B1(n_92), .B2(n_93), .Y(n_698) );
NAND2x1p5_ASAP7_75t_L g699 ( .A(n_607), .B(n_115), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_546), .A2(n_116), .B(n_119), .Y(n_700) );
OAI22x1_ASAP7_75t_L g701 ( .A1(n_604), .A2(n_120), .B1(n_122), .B2(n_123), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_592), .Y(n_702) );
BUFx10_ASAP7_75t_L g703 ( .A(n_592), .Y(n_703) );
BUFx12f_ASAP7_75t_L g704 ( .A(n_614), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_552), .Y(n_705) );
BUFx3_ASAP7_75t_L g706 ( .A(n_564), .Y(n_706) );
BUFx3_ASAP7_75t_L g707 ( .A(n_565), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_551), .A2(n_134), .B(n_135), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_552), .B(n_589), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_541), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_562), .B(n_136), .C(n_137), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_596), .A2(n_611), .B1(n_612), .B2(n_580), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_625), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_589), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_599), .A2(n_141), .B(n_142), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_617), .A2(n_598), .B(n_628), .C(n_638), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_590), .A2(n_143), .B1(n_144), .B2(n_146), .Y(n_717) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_548), .Y(n_718) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_560), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_548), .B(n_148), .Y(n_720) );
BUFx10_ASAP7_75t_L g721 ( .A(n_614), .Y(n_721) );
OAI21x1_ASAP7_75t_L g722 ( .A1(n_630), .A2(n_151), .B(n_152), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_553), .Y(n_723) );
AO31x2_ASAP7_75t_L g724 ( .A1(n_623), .A2(n_161), .A3(n_164), .B(n_165), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_618), .A2(n_168), .B1(n_169), .B2(n_173), .Y(n_725) );
OAI22x1_ASAP7_75t_L g726 ( .A1(n_627), .A2(n_180), .B1(n_181), .B2(n_184), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_566), .Y(n_727) );
OR2x6_ASAP7_75t_L g728 ( .A(n_567), .B(n_190), .Y(n_728) );
INVx3_ASAP7_75t_L g729 ( .A(n_567), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_636), .A2(n_193), .B1(n_194), .B2(n_195), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_636), .B(n_196), .Y(n_731) );
O2A1O1Ixp33_ASAP7_75t_SL g732 ( .A1(n_619), .A2(n_197), .B(n_199), .C(n_202), .Y(n_732) );
INVx5_ASAP7_75t_L g733 ( .A(n_614), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_624), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_616), .A2(n_203), .B(n_204), .Y(n_735) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_560), .Y(n_736) );
INVx4_ASAP7_75t_L g737 ( .A(n_560), .Y(n_737) );
AO31x2_ASAP7_75t_L g738 ( .A1(n_622), .A2(n_207), .A3(n_209), .B(n_210), .Y(n_738) );
INVx5_ASAP7_75t_SL g739 ( .A(n_563), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g740 ( .A1(n_615), .A2(n_213), .B(n_214), .C(n_216), .Y(n_740) );
AO22x1_ASAP7_75t_SL g741 ( .A1(n_635), .A2(n_217), .B1(n_218), .B2(n_219), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_620), .A2(n_220), .B1(n_222), .B2(n_223), .Y(n_742) );
O2A1O1Ixp33_ASAP7_75t_L g743 ( .A1(n_615), .A2(n_225), .B(n_232), .C(n_631), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_563), .B(n_569), .Y(n_744) );
BUFx5_ASAP7_75t_L g745 ( .A(n_583), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_585), .A2(n_600), .B(n_587), .C(n_571), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_600), .A2(n_472), .B(n_439), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_571), .A2(n_574), .B1(n_554), .B2(n_531), .Y(n_748) );
OR2x6_ASAP7_75t_L g749 ( .A(n_670), .B(n_728), .Y(n_749) );
OAI21xp33_ASAP7_75t_L g750 ( .A1(n_746), .A2(n_709), .B(n_649), .Y(n_750) );
OAI211xp5_ASAP7_75t_L g751 ( .A1(n_681), .A2(n_667), .B(n_698), .C(n_644), .Y(n_751) );
OAI21xp5_ASAP7_75t_L g752 ( .A1(n_747), .A2(n_642), .B(n_657), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_714), .B(n_693), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_680), .B(n_703), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_640), .Y(n_755) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_688), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_676), .Y(n_757) );
INVx1_ASAP7_75t_SL g758 ( .A(n_645), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_690), .B(n_702), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_646), .B(n_648), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_687), .A2(n_671), .B1(n_673), .B2(n_712), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_686), .B(n_662), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_692), .B(n_654), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_674), .B(n_660), .Y(n_764) );
BUFx2_ASAP7_75t_L g765 ( .A(n_665), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_694), .A2(n_732), .B(n_695), .Y(n_766) );
OAI22x1_ASAP7_75t_L g767 ( .A1(n_687), .A2(n_658), .B1(n_666), .B2(n_653), .Y(n_767) );
INVx6_ASAP7_75t_L g768 ( .A(n_734), .Y(n_768) );
OA21x2_ASAP7_75t_L g769 ( .A1(n_651), .A2(n_722), .B(n_697), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_647), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_691), .B(n_723), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_728), .B(n_720), .Y(n_772) );
AO21x2_ASAP7_75t_L g773 ( .A1(n_743), .A2(n_740), .B(n_700), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_691), .B(n_713), .Y(n_774) );
AO21x2_ASAP7_75t_L g775 ( .A1(n_708), .A2(n_742), .B(n_679), .Y(n_775) );
OA21x2_ASAP7_75t_L g776 ( .A1(n_735), .A2(n_731), .B(n_730), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_699), .A2(n_668), .B1(n_683), .B2(n_661), .Y(n_777) );
AO31x2_ASAP7_75t_L g778 ( .A1(n_726), .A2(n_701), .A3(n_725), .B(n_663), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_664), .A2(n_656), .B1(n_675), .B2(n_707), .Y(n_779) );
OA21x2_ASAP7_75t_L g780 ( .A1(n_727), .A2(n_711), .B(n_641), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_739), .Y(n_781) );
AND2x4_ASAP7_75t_L g782 ( .A(n_729), .B(n_706), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_744), .B(n_718), .Y(n_783) );
BUFx3_ASAP7_75t_L g784 ( .A(n_704), .Y(n_784) );
AO31x2_ASAP7_75t_L g785 ( .A1(n_652), .A2(n_650), .A3(n_655), .B(n_741), .Y(n_785) );
AO31x2_ASAP7_75t_L g786 ( .A1(n_668), .A2(n_737), .A3(n_643), .B(n_738), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_659), .Y(n_787) );
AND2x4_ASAP7_75t_L g788 ( .A(n_733), .B(n_710), .Y(n_788) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_739), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_745), .B(n_736), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_659), .Y(n_791) );
BUFx12f_ASAP7_75t_L g792 ( .A(n_721), .Y(n_792) );
OAI21x1_ASAP7_75t_L g793 ( .A1(n_745), .A2(n_736), .B(n_719), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_643), .B(n_745), .Y(n_794) );
AND2x4_ASAP7_75t_L g795 ( .A(n_733), .B(n_736), .Y(n_795) );
AO21x2_ASAP7_75t_L g796 ( .A1(n_677), .A2(n_689), .B(n_724), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_717), .A2(n_710), .B1(n_678), .B2(n_684), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_689), .A2(n_678), .B(n_684), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_696), .B(n_672), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_696), .B(n_530), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_L g801 ( .A1(n_746), .A2(n_649), .B(n_672), .C(n_669), .Y(n_801) );
AO21x2_ASAP7_75t_L g802 ( .A1(n_746), .A2(n_642), .B(n_715), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_716), .A2(n_642), .B(n_571), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_716), .A2(n_642), .B(n_571), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_639), .Y(n_805) );
A2O1A1Ixp33_ASAP7_75t_L g806 ( .A1(n_746), .A2(n_649), .B(n_672), .C(n_669), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_645), .B(n_530), .Y(n_807) );
OAI21x1_ASAP7_75t_SL g808 ( .A1(n_748), .A2(n_715), .B(n_581), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_672), .B(n_531), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_705), .A2(n_604), .B1(n_593), .B2(n_488), .Y(n_810) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_645), .Y(n_811) );
INVx3_ASAP7_75t_L g812 ( .A(n_670), .Y(n_812) );
BUFx2_ASAP7_75t_SL g813 ( .A(n_682), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_639), .Y(n_814) );
AO31x2_ASAP7_75t_L g815 ( .A1(n_642), .A2(n_746), .A3(n_716), .B(n_748), .Y(n_815) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_670), .Y(n_816) );
OR2x2_ASAP7_75t_L g817 ( .A(n_645), .B(n_530), .Y(n_817) );
BUFx12f_ASAP7_75t_L g818 ( .A(n_685), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_680), .B(n_530), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_680), .B(n_530), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_705), .A2(n_604), .B1(n_593), .B2(n_488), .Y(n_821) );
AO21x2_ASAP7_75t_L g822 ( .A1(n_746), .A2(n_642), .B(n_715), .Y(n_822) );
OAI221xp5_ASAP7_75t_SL g823 ( .A1(n_644), .A2(n_491), .B1(n_410), .B2(n_488), .C(n_446), .Y(n_823) );
OR2x2_ASAP7_75t_L g824 ( .A(n_645), .B(n_530), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_705), .A2(n_604), .B1(n_593), .B2(n_488), .Y(n_825) );
O2A1O1Ixp33_ASAP7_75t_L g826 ( .A1(n_709), .A2(n_746), .B(n_534), .C(n_705), .Y(n_826) );
AOI21xp5_ASAP7_75t_L g827 ( .A1(n_716), .A2(n_642), .B(n_571), .Y(n_827) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_817), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_824), .Y(n_829) );
INVx5_ASAP7_75t_L g830 ( .A(n_749), .Y(n_830) );
OA21x2_ASAP7_75t_L g831 ( .A1(n_798), .A2(n_804), .B(n_803), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_805), .B(n_814), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_749), .A2(n_761), .B1(n_760), .B2(n_809), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_818), .Y(n_834) );
OR2x6_ASAP7_75t_L g835 ( .A(n_749), .B(n_808), .Y(n_835) );
OAI222xp33_ASAP7_75t_L g836 ( .A1(n_777), .A2(n_823), .B1(n_797), .B2(n_757), .C1(n_763), .C2(n_758), .Y(n_836) );
AO21x2_ASAP7_75t_L g837 ( .A1(n_827), .A2(n_752), .B(n_766), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_774), .B(n_753), .Y(n_838) );
OA21x2_ASAP7_75t_L g839 ( .A1(n_750), .A2(n_752), .B(n_794), .Y(n_839) );
INVxp67_ASAP7_75t_L g840 ( .A(n_811), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_751), .A2(n_754), .B1(n_819), .B2(n_820), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_787), .Y(n_842) );
INVx3_ASAP7_75t_L g843 ( .A(n_756), .Y(n_843) );
NAND2x1_ASAP7_75t_L g844 ( .A(n_769), .B(n_791), .Y(n_844) );
INVx3_ASAP7_75t_L g845 ( .A(n_756), .Y(n_845) );
NAND3xp33_ASAP7_75t_L g846 ( .A(n_826), .B(n_801), .C(n_806), .Y(n_846) );
AO21x2_ASAP7_75t_L g847 ( .A1(n_796), .A2(n_822), .B(n_802), .Y(n_847) );
OAI211xp5_ASAP7_75t_L g848 ( .A1(n_810), .A2(n_825), .B(n_821), .C(n_779), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_799), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_764), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_764), .Y(n_851) );
BUFx2_ASAP7_75t_L g852 ( .A(n_790), .Y(n_852) );
NAND4xp25_ASAP7_75t_L g853 ( .A(n_755), .B(n_762), .C(n_759), .D(n_800), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_786), .B(n_783), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_770), .B(n_816), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_786), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_767), .A2(n_784), .B1(n_765), .B2(n_792), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_778), .B(n_815), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_785), .B(n_782), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_815), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_793), .Y(n_861) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_812), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_812), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_782), .B(n_778), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_768), .A2(n_773), .B1(n_813), .B2(n_781), .Y(n_865) );
OA21x2_ASAP7_75t_L g866 ( .A1(n_780), .A2(n_795), .B(n_788), .Y(n_866) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_789), .Y(n_867) );
OA21x2_ASAP7_75t_L g868 ( .A1(n_775), .A2(n_776), .B(n_768), .Y(n_868) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_807), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_774), .B(n_772), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_771), .Y(n_871) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_807), .Y(n_872) );
BUFx2_ASAP7_75t_L g873 ( .A(n_835), .Y(n_873) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_852), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_842), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_842), .Y(n_876) );
BUFx2_ASAP7_75t_L g877 ( .A(n_835), .Y(n_877) );
INVx3_ASAP7_75t_L g878 ( .A(n_868), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_864), .B(n_854), .Y(n_879) );
OR2x2_ASAP7_75t_L g880 ( .A(n_870), .B(n_838), .Y(n_880) );
INVx2_ASAP7_75t_SL g881 ( .A(n_830), .Y(n_881) );
BUFx3_ASAP7_75t_L g882 ( .A(n_830), .Y(n_882) );
AND2x4_ASAP7_75t_L g883 ( .A(n_835), .B(n_859), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_858), .B(n_871), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_850), .B(n_851), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_859), .B(n_832), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_866), .Y(n_887) );
OR2x2_ASAP7_75t_L g888 ( .A(n_853), .B(n_849), .Y(n_888) );
BUFx2_ASAP7_75t_L g889 ( .A(n_835), .Y(n_889) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_866), .Y(n_890) );
NOR3xp33_ASAP7_75t_SL g891 ( .A(n_834), .B(n_848), .C(n_836), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_856), .B(n_860), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_831), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_844), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_875), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_875), .Y(n_896) );
BUFx2_ASAP7_75t_L g897 ( .A(n_874), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_886), .B(n_839), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_876), .Y(n_899) );
INVx3_ASAP7_75t_L g900 ( .A(n_878), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_886), .B(n_839), .Y(n_901) );
OR2x2_ASAP7_75t_L g902 ( .A(n_880), .B(n_839), .Y(n_902) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_891), .A2(n_841), .B1(n_865), .B2(n_857), .C(n_833), .Y(n_903) );
AND2x4_ASAP7_75t_L g904 ( .A(n_883), .B(n_865), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_879), .B(n_847), .Y(n_905) );
AND2x2_ASAP7_75t_SL g906 ( .A(n_873), .B(n_868), .Y(n_906) );
AND2x4_ASAP7_75t_L g907 ( .A(n_883), .B(n_861), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_884), .B(n_831), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_884), .B(n_831), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_888), .B(n_837), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_895), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_896), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_905), .B(n_887), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_896), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_899), .Y(n_915) );
AND2x4_ASAP7_75t_L g916 ( .A(n_907), .B(n_894), .Y(n_916) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_897), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_898), .B(n_890), .Y(n_918) );
NOR2x1p5_ASAP7_75t_SL g919 ( .A(n_910), .B(n_893), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_898), .B(n_892), .Y(n_920) );
OAI22xp33_ASAP7_75t_L g921 ( .A1(n_903), .A2(n_873), .B1(n_889), .B2(n_877), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_901), .B(n_892), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_901), .B(n_892), .Y(n_923) );
INVx3_ASAP7_75t_L g924 ( .A(n_900), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_918), .B(n_908), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_918), .B(n_908), .Y(n_926) );
OR2x2_ASAP7_75t_L g927 ( .A(n_913), .B(n_902), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_911), .Y(n_928) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_917), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_920), .B(n_909), .Y(n_930) );
AND2x4_ASAP7_75t_L g931 ( .A(n_919), .B(n_904), .Y(n_931) );
O2A1O1Ixp33_ASAP7_75t_L g932 ( .A1(n_921), .A2(n_840), .B(n_867), .C(n_872), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_912), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_914), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_929), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_933), .Y(n_936) );
O2A1O1Ixp33_ASAP7_75t_L g937 ( .A1(n_932), .A2(n_828), .B(n_829), .C(n_869), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_927), .B(n_922), .Y(n_938) );
OA21x2_ASAP7_75t_L g939 ( .A1(n_931), .A2(n_893), .B(n_915), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_928), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_930), .B(n_923), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_934), .Y(n_942) );
INVx3_ASAP7_75t_L g943 ( .A(n_939), .Y(n_943) );
INVxp67_ASAP7_75t_L g944 ( .A(n_935), .Y(n_944) );
O2A1O1Ixp33_ASAP7_75t_L g945 ( .A1(n_937), .A2(n_863), .B(n_862), .C(n_855), .Y(n_945) );
A2O1A1Ixp33_ASAP7_75t_L g946 ( .A1(n_938), .A2(n_919), .B(n_925), .C(n_926), .Y(n_946) );
OAI211xp5_ASAP7_75t_L g947 ( .A1(n_946), .A2(n_846), .B(n_940), .C(n_941), .Y(n_947) );
NAND3xp33_ASAP7_75t_L g948 ( .A(n_944), .B(n_942), .C(n_936), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_947), .B(n_943), .C(n_945), .Y(n_949) );
AND2x4_ASAP7_75t_L g950 ( .A(n_949), .B(n_948), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_950), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_951), .Y(n_952) );
BUFx6f_ASAP7_75t_L g953 ( .A(n_952), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_953), .A2(n_924), .B1(n_881), .B2(n_882), .Y(n_954) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_954), .B(n_843), .C(n_845), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_955), .A2(n_881), .B(n_885), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_956), .A2(n_916), .B1(n_900), .B2(n_906), .Y(n_957) );
endmodule