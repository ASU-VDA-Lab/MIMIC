module fake_netlist_5_1848_n_891 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_891);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_891;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_864;
wire n_859;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_867;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_171;
wire n_756;
wire n_878;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_862;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_570;
wire n_457;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_834;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_632;
wire n_489;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_170;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_884;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_647;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_180;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_163),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_57),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_138),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_62),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_82),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_131),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_77),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_134),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_75),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_52),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_120),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_29),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_10),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_43),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_98),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_108),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_42),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_16),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_156),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_91),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_71),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_119),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_88),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_85),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_63),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_83),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_66),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_155),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_58),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_6),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_61),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_127),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_99),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_78),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_44),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_68),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_29),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_11),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_72),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_165),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_3),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_28),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_26),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_87),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_32),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_153),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_38),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_145),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_45),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_139),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_146),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_118),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_161),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_5),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_166),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_89),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_80),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_79),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_111),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_122),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_55),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_14),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_157),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

AND2x4_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_218),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_0),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_225),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_189),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_0),
.Y(n_260)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_178),
.B(n_1),
.Y(n_262)
);

BUFx8_ASAP7_75t_SL g263 ( 
.A(n_167),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_196),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_30),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_189),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_211),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_186),
.B(n_1),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_205),
.B(n_2),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx6p67_ASAP7_75t_R g273 ( 
.A(n_215),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_219),
.B(n_2),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_205),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_193),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_201),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_168),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_170),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_224),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_193),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_173),
.Y(n_286)
);

BUFx8_ASAP7_75t_SL g287 ( 
.A(n_179),
.Y(n_287)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_193),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_186),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_210),
.B(n_3),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_169),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_217),
.B(n_4),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g297 ( 
.A(n_217),
.B(n_31),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_171),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g302 ( 
.A(n_174),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_172),
.B(n_33),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_180),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_242),
.Y(n_305)
);

CKINVDCx6p67_ASAP7_75t_R g306 ( 
.A(n_190),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_242),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_201),
.B(n_4),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_188),
.B(n_34),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_181),
.B(n_5),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_282),
.B(n_191),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_255),
.A2(n_198),
.B1(n_200),
.B2(n_208),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_175),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_268),
.B1(n_264),
.B2(n_260),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g318 ( 
.A1(n_262),
.A2(n_297),
.B1(n_265),
.B2(n_274),
.Y(n_318)
);

AO22x2_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_216),
.B1(n_241),
.B2(n_236),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_264),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_6),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_195),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_R g323 ( 
.A1(n_277),
.A2(n_251),
.B1(n_235),
.B2(n_226),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_268),
.A2(n_244),
.B1(n_248),
.B2(n_246),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_256),
.A2(n_249),
.B1(n_245),
.B2(n_243),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_301),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_176),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_273),
.A2(n_240),
.B1(n_238),
.B2(n_237),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_177),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_308),
.A2(n_206),
.B1(n_197),
.B2(n_204),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_265),
.A2(n_212),
.B1(n_214),
.B2(n_220),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_286),
.B(n_182),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_183),
.Y(n_334)
);

OA22x2_ASAP7_75t_L g335 ( 
.A1(n_258),
.A2(n_234),
.B1(n_232),
.B2(n_231),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_L g337 ( 
.A1(n_273),
.A2(n_230),
.B1(n_229),
.B2(n_223),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_301),
.Y(n_340)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_297),
.B(n_7),
.Y(n_341)
);

AO22x2_ASAP7_75t_L g342 ( 
.A1(n_265),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_294),
.A2(n_222),
.B1(n_213),
.B2(n_209),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_283),
.A2(n_207),
.B1(n_203),
.B2(n_202),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_254),
.A2(n_199),
.B1(n_194),
.B2(n_192),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_253),
.B(n_300),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_254),
.A2(n_185),
.B1(n_184),
.B2(n_201),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_267),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_272),
.A2(n_201),
.B1(n_9),
.B2(n_11),
.Y(n_352)
);

AO22x2_ASAP7_75t_L g353 ( 
.A1(n_253),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_283),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g356 ( 
.A1(n_272),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_356)
);

NAND3x1_ASAP7_75t_L g357 ( 
.A(n_271),
.B(n_15),
.C(n_17),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_291),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_253),
.B(n_201),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_291),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g362 ( 
.A1(n_306),
.A2(n_289),
.B1(n_292),
.B2(n_270),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g363 ( 
.A1(n_306),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_276),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_360),
.Y(n_365)
);

NAND2x1p5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_348),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_345),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_340),
.A2(n_359),
.B(n_318),
.Y(n_370)
);

OR2x6_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_302),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_302),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_343),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_311),
.B(n_303),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_305),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_321),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_333),
.B(n_303),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_355),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_320),
.B(n_305),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_324),
.B(n_263),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g384 ( 
.A(n_352),
.B(n_303),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_315),
.B(n_325),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_322),
.B(n_309),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_307),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_318),
.B(n_309),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_346),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_309),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_334),
.B(n_307),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_332),
.B(n_296),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_317),
.B(n_263),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_SL g402 ( 
.A(n_354),
.B(n_270),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_314),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_335),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_347),
.B(n_287),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_319),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_319),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_330),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_328),
.B(n_287),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_344),
.B(n_337),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_350),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_357),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_269),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_358),
.B(n_275),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_363),
.B(n_296),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_324),
.B(n_35),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_348),
.B(n_275),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_311),
.B(n_296),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_345),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_348),
.B(n_275),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_375),
.B(n_269),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_281),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_395),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_281),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_387),
.B(n_280),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_395),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_409),
.B(n_36),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_390),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_394),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

AND2x2_ASAP7_75t_SL g448 ( 
.A(n_384),
.B(n_280),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_376),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_392),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_393),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_370),
.A2(n_374),
.B(n_389),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_410),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_374),
.B(n_281),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_298),
.Y(n_459)
);

BUFx5_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_SL g461 ( 
.A(n_385),
.B(n_298),
.C(n_22),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_401),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_L g463 ( 
.A(n_370),
.B(n_298),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_396),
.B(n_276),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_408),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_428),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_389),
.B(n_37),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_365),
.B(n_39),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_276),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_390),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_366),
.B(n_420),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_366),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_372),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_429),
.A2(n_261),
.B(n_266),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_420),
.B(n_276),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_373),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_369),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_406),
.B(n_21),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_378),
.B(n_40),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_SL g484 ( 
.A(n_412),
.B(n_261),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_406),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_425),
.B(n_261),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_433),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_417),
.B(n_23),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_426),
.B(n_261),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_399),
.B(n_278),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_399),
.B(n_278),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_417),
.B(n_24),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_430),
.B(n_278),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_368),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_379),
.B(n_380),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_423),
.B(n_25),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_368),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_381),
.B(n_261),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_368),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_416),
.A2(n_295),
.B1(n_290),
.B2(n_285),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_422),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_437),
.B(n_441),
.Y(n_504)
);

BUFx12f_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

BUFx4f_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_503),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_503),
.Y(n_508)
);

CKINVDCx6p67_ASAP7_75t_R g509 ( 
.A(n_449),
.Y(n_509)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_468),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_448),
.B(n_419),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_466),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_437),
.B(n_414),
.Y(n_513)
);

BUFx2_ASAP7_75t_R g514 ( 
.A(n_452),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_448),
.B(n_488),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_475),
.B(n_371),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_440),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_473),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_442),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_465),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_474),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_485),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_440),
.Y(n_523)
);

NOR2x1_ASAP7_75t_R g524 ( 
.A(n_475),
.B(n_419),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_466),
.B(n_422),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_452),
.B(n_415),
.Y(n_526)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_455),
.B(n_427),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_452),
.B(n_371),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_447),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_447),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_443),
.B(n_421),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_452),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_441),
.B(n_371),
.Y(n_533)
);

BUFx8_ASAP7_75t_L g534 ( 
.A(n_474),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_456),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_477),
.B(n_498),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_448),
.B(n_367),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_450),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_481),
.B(n_431),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_464),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_492),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_481),
.B(n_413),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_468),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_482),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_494),
.B(n_411),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_442),
.B(n_418),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_468),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_434),
.B(n_413),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_439),
.B(n_402),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_451),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_442),
.B(n_413),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_434),
.B(n_400),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_439),
.B(n_278),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_469),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_442),
.B(n_41),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_461),
.B(n_383),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_469),
.B(n_46),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_496),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_469),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_483),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

NAND2x1p5_ASAP7_75t_L g564 ( 
.A(n_519),
.B(n_499),
.Y(n_564)
);

NAND2x1p5_ASAP7_75t_L g565 ( 
.A(n_519),
.B(n_499),
.Y(n_565)
);

NAND2x1p5_ASAP7_75t_L g566 ( 
.A(n_506),
.B(n_499),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_559),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_559),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_561),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_508),
.Y(n_570)
);

CKINVDCx11_ASAP7_75t_R g571 ( 
.A(n_509),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_518),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_505),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_522),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_492),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_543),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_534),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_526),
.Y(n_578)
);

BUFx2_ASAP7_75t_SL g579 ( 
.A(n_552),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_545),
.B(n_493),
.Y(n_580)
);

INVx3_ASAP7_75t_SL g581 ( 
.A(n_547),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_542),
.B(n_479),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_538),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_523),
.Y(n_585)
);

NAND2x1p5_ASAP7_75t_L g586 ( 
.A(n_506),
.B(n_499),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_520),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_552),
.Y(n_588)
);

BUFx4f_ASAP7_75t_L g589 ( 
.A(n_547),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_510),
.B(n_483),
.Y(n_590)
);

BUFx24_ASAP7_75t_L g591 ( 
.A(n_540),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_526),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_510),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_530),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_537),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_535),
.Y(n_596)
);

NAND2x1p5_ASAP7_75t_L g597 ( 
.A(n_556),
.B(n_483),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_529),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_534),
.Y(n_599)
);

BUFx12f_ASAP7_75t_L g600 ( 
.A(n_516),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_536),
.B(n_493),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_539),
.Y(n_602)
);

BUFx24_ASAP7_75t_L g603 ( 
.A(n_540),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_525),
.Y(n_604)
);

CKINVDCx6p67_ASAP7_75t_R g605 ( 
.A(n_516),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_538),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_542),
.B(n_479),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_504),
.B(n_464),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_551),
.Y(n_609)
);

BUFx4_ASAP7_75t_SL g610 ( 
.A(n_516),
.Y(n_610)
);

CKINVDCx6p67_ASAP7_75t_R g611 ( 
.A(n_528),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_521),
.Y(n_612)
);

CKINVDCx11_ASAP7_75t_R g613 ( 
.A(n_571),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_609),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_578),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_609),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_575),
.A2(n_546),
.B1(n_527),
.B2(n_515),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_585),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_571),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_601),
.A2(n_546),
.B1(n_515),
.B2(n_511),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_584),
.B(n_521),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_583),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_598),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_599),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_602),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_580),
.B(n_531),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_583),
.Y(n_627)
);

INVx3_ASAP7_75t_SL g628 ( 
.A(n_599),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_588),
.A2(n_511),
.B1(n_525),
.B2(n_544),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_597),
.A2(n_560),
.B1(n_555),
.B2(n_548),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_582),
.B(n_550),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_572),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_563),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_594),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_589),
.A2(n_556),
.B1(n_558),
.B2(n_533),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_597),
.A2(n_510),
.B1(n_533),
.B2(n_513),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_594),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_606),
.A2(n_558),
.B1(n_557),
.B2(n_528),
.Y(n_638)
);

CKINVDCx11_ASAP7_75t_R g639 ( 
.A(n_577),
.Y(n_639)
);

CKINVDCx6p67_ASAP7_75t_R g640 ( 
.A(n_591),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_595),
.Y(n_641)
);

CKINVDCx6p67_ASAP7_75t_R g642 ( 
.A(n_591),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_608),
.A2(n_541),
.B1(n_483),
.B2(n_462),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_589),
.A2(n_603),
.B1(n_576),
.B2(n_579),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_587),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_607),
.A2(n_451),
.B1(n_462),
.B2(n_454),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_603),
.Y(n_647)
);

INVx6_ASAP7_75t_L g648 ( 
.A(n_578),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_574),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_595),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_612),
.A2(n_553),
.B1(n_446),
.B2(n_445),
.Y(n_651)
);

INVx6_ASAP7_75t_L g652 ( 
.A(n_578),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_SL g653 ( 
.A1(n_577),
.A2(n_514),
.B1(n_478),
.B2(n_446),
.Y(n_653)
);

INVx6_ASAP7_75t_L g654 ( 
.A(n_578),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_562),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_590),
.A2(n_445),
.B1(n_512),
.B2(n_532),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_614),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_631),
.B(n_612),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_649),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_621),
.B(n_626),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_617),
.A2(n_581),
.B1(n_604),
.B2(n_600),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_SL g662 ( 
.A1(n_647),
.A2(n_600),
.B1(n_573),
.B2(n_604),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_616),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_613),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_620),
.A2(n_581),
.B1(n_512),
.B2(n_605),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_618),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_630),
.A2(n_573),
.B1(n_593),
.B2(n_587),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_620),
.A2(n_590),
.B1(n_605),
.B2(n_611),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_638),
.A2(n_611),
.B1(n_569),
.B2(n_590),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_640),
.A2(n_573),
.B1(n_596),
.B2(n_569),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_655),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_638),
.A2(n_407),
.B1(n_573),
.B2(n_592),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_627),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_651),
.B(n_592),
.Y(n_674)
);

CKINVDCx11_ASAP7_75t_R g675 ( 
.A(n_619),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_622),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_SL g677 ( 
.A1(n_636),
.A2(n_593),
.B1(n_569),
.B2(n_563),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_653),
.A2(n_569),
.B1(n_592),
.B2(n_453),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_653),
.A2(n_592),
.B1(n_453),
.B2(n_472),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_635),
.A2(n_593),
.B1(n_586),
.B2(n_566),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_651),
.A2(n_454),
.B1(n_472),
.B2(n_532),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_SL g682 ( 
.A1(n_644),
.A2(n_502),
.B(n_436),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_642),
.A2(n_570),
.B1(n_487),
.B2(n_490),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_644),
.A2(n_502),
.B(n_438),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_629),
.A2(n_487),
.B1(n_490),
.B2(n_495),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_632),
.A2(n_495),
.B1(n_497),
.B2(n_470),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_650),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_633),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_643),
.A2(n_470),
.B1(n_501),
.B2(n_491),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_643),
.A2(n_501),
.B1(n_491),
.B2(n_480),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_SL g691 ( 
.A1(n_624),
.A2(n_593),
.B1(n_563),
.B2(n_586),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_634),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_633),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_648),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_623),
.Y(n_695)
);

AOI222xp33_ASAP7_75t_L g696 ( 
.A1(n_628),
.A2(n_524),
.B1(n_457),
.B2(n_463),
.C1(n_459),
.C2(n_554),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_645),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_656),
.A2(n_480),
.B1(n_491),
.B2(n_463),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_637),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_615),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_615),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_641),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_625),
.B(n_524),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_615),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_648),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_648),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_652),
.Y(n_707)
);

INVx4_ASAP7_75t_L g708 ( 
.A(n_652),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_646),
.A2(n_480),
.B1(n_566),
.B2(n_484),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_661),
.A2(n_628),
.B1(n_639),
.B2(n_646),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_SL g711 ( 
.A1(n_672),
.A2(n_610),
.B(n_564),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_660),
.A2(n_654),
.B1(n_652),
.B2(n_568),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_SL g713 ( 
.A1(n_668),
.A2(n_654),
.B1(n_610),
.B2(n_568),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_665),
.A2(n_654),
.B1(n_568),
.B2(n_567),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_669),
.A2(n_484),
.B1(n_568),
.B2(n_567),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_658),
.B(n_567),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_674),
.A2(n_659),
.B1(n_684),
.B2(n_682),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_679),
.A2(n_567),
.B1(n_460),
.B2(n_564),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_678),
.A2(n_460),
.B1(n_565),
.B2(n_496),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_703),
.A2(n_565),
.B1(n_496),
.B2(n_476),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_696),
.A2(n_460),
.B1(n_496),
.B2(n_489),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_667),
.A2(n_460),
.B1(n_496),
.B2(n_486),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_683),
.A2(n_662),
.B1(n_686),
.B2(n_681),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_677),
.A2(n_460),
.B1(n_476),
.B2(n_435),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_SL g725 ( 
.A1(n_680),
.A2(n_285),
.B1(n_290),
.B2(n_295),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_691),
.A2(n_697),
.B1(n_685),
.B2(n_675),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_666),
.A2(n_285),
.B1(n_290),
.B2(n_295),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_SL g728 ( 
.A(n_664),
.B(n_500),
.C(n_26),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_670),
.A2(n_460),
.B1(n_435),
.B2(n_458),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_675),
.A2(n_460),
.B1(n_444),
.B2(n_435),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_695),
.A2(n_295),
.B1(n_285),
.B2(n_290),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_671),
.A2(n_460),
.B1(n_458),
.B2(n_444),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_671),
.A2(n_460),
.B1(n_458),
.B2(n_444),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_707),
.A2(n_471),
.B1(n_467),
.B2(n_288),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_709),
.B(n_288),
.C(n_266),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_664),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_689),
.A2(n_471),
.B1(n_467),
.B2(n_288),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_657),
.B(n_27),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_673),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_705),
.A2(n_471),
.B1(n_467),
.B2(n_288),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_705),
.A2(n_467),
.B1(n_471),
.B2(n_288),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_705),
.A2(n_266),
.B1(n_48),
.B2(n_49),
.Y(n_742)
);

OA21x2_ASAP7_75t_L g743 ( 
.A1(n_673),
.A2(n_47),
.B(n_50),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_657),
.A2(n_266),
.B1(n_53),
.B2(n_54),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_SL g745 ( 
.A1(n_688),
.A2(n_266),
.B1(n_56),
.B2(n_59),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_SL g746 ( 
.A1(n_688),
.A2(n_51),
.B1(n_60),
.B2(n_64),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_663),
.B(n_65),
.C(n_67),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_663),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_694),
.A2(n_74),
.B1(n_81),
.B2(n_84),
.Y(n_749)
);

OAI21xp33_ASAP7_75t_L g750 ( 
.A1(n_736),
.A2(n_728),
.B(n_710),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_717),
.B(n_692),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_717),
.B(n_692),
.C(n_699),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_716),
.B(n_699),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_739),
.B(n_702),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_738),
.B(n_702),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_726),
.B(n_676),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_743),
.B(n_676),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_713),
.B(n_687),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_743),
.B(n_687),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_712),
.B(n_700),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_711),
.A2(n_690),
.B1(n_708),
.B2(n_706),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_723),
.B(n_706),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_714),
.B(n_693),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_721),
.B(n_688),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_747),
.A2(n_708),
.B1(n_694),
.B2(n_693),
.Y(n_765)
);

OAI221xp5_ASAP7_75t_SL g766 ( 
.A1(n_749),
.A2(n_698),
.B1(n_701),
.B2(n_704),
.C(n_693),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_730),
.B(n_704),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_720),
.B(n_708),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_743),
.B(n_704),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_SL g770 ( 
.A(n_735),
.B(n_701),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_722),
.B(n_701),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_L g772 ( 
.A(n_748),
.B(n_86),
.C(n_90),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_725),
.B(n_92),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_724),
.B(n_93),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_715),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_746),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_776)
);

AND2x2_ASAP7_75t_SL g777 ( 
.A(n_719),
.B(n_104),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_718),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_745),
.B(n_110),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_729),
.B(n_744),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_742),
.B(n_113),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_754),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_769),
.B(n_727),
.Y(n_783)
);

NAND4xp75_ASAP7_75t_L g784 ( 
.A(n_751),
.B(n_741),
.C(n_731),
.D(n_116),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_769),
.B(n_734),
.Y(n_785)
);

NOR2x1_ASAP7_75t_L g786 ( 
.A(n_752),
.B(n_755),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_754),
.B(n_733),
.Y(n_787)
);

NOR2x1_ASAP7_75t_L g788 ( 
.A(n_752),
.B(n_732),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_SL g789 ( 
.A(n_766),
.B(n_114),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_757),
.B(n_737),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_753),
.B(n_115),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_757),
.B(n_740),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_750),
.A2(n_117),
.B1(n_121),
.B2(n_123),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_759),
.B(n_124),
.Y(n_794)
);

AOI211xp5_ASAP7_75t_L g795 ( 
.A1(n_750),
.A2(n_125),
.B(n_126),
.C(n_128),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_759),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_762),
.B(n_129),
.C(n_130),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_763),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_760),
.B(n_132),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_796),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_782),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_796),
.B(n_756),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_782),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_798),
.B(n_758),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_782),
.B(n_768),
.Y(n_805)
);

NAND4xp75_ASAP7_75t_L g806 ( 
.A(n_793),
.B(n_777),
.C(n_779),
.D(n_773),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_786),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_798),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_799),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_785),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_785),
.B(n_792),
.Y(n_811)
);

OA22x2_ASAP7_75t_L g812 ( 
.A1(n_807),
.A2(n_783),
.B1(n_794),
.B2(n_761),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_810),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_808),
.Y(n_814)
);

XOR2x2_ASAP7_75t_L g815 ( 
.A(n_806),
.B(n_795),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_807),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_801),
.Y(n_817)
);

OAI22x1_ASAP7_75t_L g818 ( 
.A1(n_816),
.A2(n_809),
.B1(n_811),
.B2(n_805),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_817),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_816),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_812),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_813),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_820),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_822),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_819),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_818),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_819),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_824),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_823),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_825),
.Y(n_830)
);

OAI221xp5_ASAP7_75t_L g831 ( 
.A1(n_829),
.A2(n_821),
.B1(n_826),
.B2(n_815),
.C(n_812),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_830),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_828),
.A2(n_821),
.B1(n_826),
.B2(n_806),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_828),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_834),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_833),
.B(n_827),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_832),
.Y(n_837)
);

NOR2x1_ASAP7_75t_L g838 ( 
.A(n_831),
.B(n_827),
.Y(n_838)
);

NOR2x1_ASAP7_75t_L g839 ( 
.A(n_833),
.B(n_797),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_832),
.B(n_811),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_833),
.A2(n_789),
.B1(n_809),
.B2(n_788),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_840),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_838),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_839),
.A2(n_836),
.B1(n_841),
.B2(n_837),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_835),
.B(n_814),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_840),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_837),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_837),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_840),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_840),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_847),
.B(n_848),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_843),
.A2(n_776),
.B1(n_784),
.B2(n_772),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_842),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_845),
.A2(n_791),
.B(n_804),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_845),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_846),
.Y(n_856)
);

AND5x1_ASAP7_75t_L g857 ( 
.A(n_844),
.B(n_770),
.C(n_805),
.D(n_794),
.E(n_777),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_851),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_855),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_853),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_856),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_857),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_852),
.A2(n_850),
.B1(n_849),
.B2(n_803),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_852),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_854),
.Y(n_865)
);

AO22x2_ASAP7_75t_L g866 ( 
.A1(n_858),
.A2(n_775),
.B1(n_773),
.B2(n_778),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_SL g867 ( 
.A1(n_858),
.A2(n_781),
.B1(n_765),
.B2(n_774),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_864),
.A2(n_783),
.B1(n_792),
.B2(n_802),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_861),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_859),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_860),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_865),
.Y(n_872)
);

AO22x2_ASAP7_75t_L g873 ( 
.A1(n_863),
.A2(n_802),
.B1(n_800),
.B2(n_780),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_869),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_870),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_872),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_871),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_873),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_874),
.A2(n_862),
.B1(n_866),
.B2(n_868),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_878),
.A2(n_876),
.B1(n_875),
.B2(n_877),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_875),
.A2(n_867),
.B1(n_780),
.B2(n_800),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_874),
.A2(n_790),
.B1(n_771),
.B2(n_767),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_880),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_879),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_881),
.Y(n_885)
);

AO22x2_ASAP7_75t_L g886 ( 
.A1(n_883),
.A2(n_882),
.B1(n_790),
.B2(n_764),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_884),
.A2(n_787),
.B1(n_140),
.B2(n_141),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_886),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_887),
.Y(n_889)
);

AO22x2_ASAP7_75t_L g890 ( 
.A1(n_888),
.A2(n_885),
.B1(n_143),
.B2(n_147),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_SL g891 ( 
.A1(n_890),
.A2(n_889),
.B1(n_787),
.B2(n_149),
.Y(n_891)
);


endmodule