module real_aes_12001_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1600;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_1606;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1584;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_0), .A2(n_248), .B1(n_360), .B2(n_361), .Y(n_359) );
INVxp33_ASAP7_75t_L g411 ( .A(n_0), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_1), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g1341 ( .A1(n_2), .A2(n_3), .B1(n_1329), .B2(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g495 ( .A(n_3), .Y(n_495) );
INVxp67_ASAP7_75t_SL g1205 ( .A(n_4), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_4), .A2(n_231), .B1(n_704), .B2(n_834), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_5), .A2(n_193), .B1(n_508), .B2(n_606), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_5), .A2(n_139), .B1(n_434), .B2(n_473), .C(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_6), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_6), .B(n_217), .Y(n_316) );
AND2x2_ASAP7_75t_L g420 ( .A(n_6), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g494 ( .A(n_6), .Y(n_494) );
INVx1_ASAP7_75t_L g1143 ( .A(n_7), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_7), .A2(n_206), .B1(n_736), .B2(n_898), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_8), .A2(n_18), .B1(n_533), .B2(n_534), .Y(n_532) );
INVx1_ASAP7_75t_L g571 ( .A(n_8), .Y(n_571) );
OA22x2_ASAP7_75t_L g647 ( .A1(n_9), .A2(n_648), .B1(n_722), .B2(n_723), .Y(n_647) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_9), .Y(n_723) );
OAI221xp5_ASAP7_75t_SL g852 ( .A1(n_10), .A2(n_61), .B1(n_853), .B2(n_855), .C(n_857), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_10), .A2(n_110), .B1(n_366), .B2(n_887), .C(n_891), .Y(n_886) );
INVx1_ASAP7_75t_L g876 ( .A(n_11), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g1165 ( .A1(n_12), .A2(n_55), .B1(n_472), .B2(n_1161), .Y(n_1165) );
INVx1_ASAP7_75t_L g1192 ( .A(n_12), .Y(n_1192) );
AOI22xp5_ASAP7_75t_L g1350 ( .A1(n_13), .A2(n_246), .B1(n_1336), .B2(n_1339), .Y(n_1350) );
CKINVDCx5p33_ASAP7_75t_R g1547 ( .A(n_14), .Y(n_1547) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_15), .A2(n_109), .B1(n_361), .B2(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g631 ( .A(n_15), .Y(n_631) );
OAI332xp33_ASAP7_75t_L g659 ( .A1(n_16), .A2(n_453), .A3(n_490), .B1(n_660), .B2(n_664), .B3(n_669), .C1(n_676), .C2(n_681), .Y(n_659) );
INVx1_ASAP7_75t_L g718 ( .A(n_16), .Y(n_718) );
INVx1_ASAP7_75t_L g917 ( .A(n_17), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_18), .A2(n_121), .B1(n_566), .B2(n_568), .C(n_570), .Y(n_565) );
CKINVDCx14_ASAP7_75t_R g1354 ( .A(n_19), .Y(n_1354) );
INVx1_ASAP7_75t_L g874 ( .A(n_20), .Y(n_874) );
INVxp67_ASAP7_75t_L g1204 ( .A(n_21), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g1232 ( .A1(n_21), .A2(n_172), .B1(n_378), .B2(n_530), .C(n_839), .Y(n_1232) );
INVxp33_ASAP7_75t_L g798 ( .A(n_22), .Y(n_798) );
AOI221xp5_ASAP7_75t_L g838 ( .A1(n_22), .A2(n_152), .B1(n_620), .B2(n_621), .C(n_839), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g954 ( .A1(n_23), .A2(n_244), .B1(n_955), .B2(n_957), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_23), .A2(n_244), .B1(n_1017), .B2(n_1019), .Y(n_1016) );
CKINVDCx5p33_ASAP7_75t_R g1532 ( .A(n_24), .Y(n_1532) );
INVx1_ASAP7_75t_L g1073 ( .A(n_25), .Y(n_1073) );
INVxp33_ASAP7_75t_L g1225 ( .A(n_26), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_26), .A2(n_105), .B1(n_932), .B2(n_1236), .Y(n_1235) );
INVx2_ASAP7_75t_L g325 ( .A(n_27), .Y(n_325) );
OR2x2_ASAP7_75t_L g339 ( .A(n_27), .B(n_323), .Y(n_339) );
INVx1_ASAP7_75t_L g845 ( .A(n_28), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g1551 ( .A(n_29), .Y(n_1551) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_30), .A2(n_50), .B1(n_534), .B2(n_739), .C(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g782 ( .A(n_30), .Y(n_782) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_31), .A2(n_74), .B1(n_440), .B2(n_802), .C(n_862), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_31), .A2(n_74), .B1(n_347), .B2(n_898), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g1096 ( .A(n_32), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_33), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g1589 ( .A1(n_34), .A2(n_146), .B1(n_919), .B2(n_923), .Y(n_1589) );
INVx1_ASAP7_75t_L g1607 ( .A(n_34), .Y(n_1607) );
OR2x2_ASAP7_75t_L g315 ( .A(n_35), .B(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g319 ( .A(n_35), .Y(n_319) );
BUFx2_ASAP7_75t_L g407 ( .A(n_35), .Y(n_407) );
INVx1_ASAP7_75t_L g419 ( .A(n_35), .Y(n_419) );
INVxp33_ASAP7_75t_L g1224 ( .A(n_36), .Y(n_1224) );
AOI21xp33_ASAP7_75t_L g1240 ( .A1(n_36), .A2(n_520), .B(n_1241), .Y(n_1240) );
CKINVDCx16_ASAP7_75t_R g1330 ( .A(n_37), .Y(n_1330) );
INVx1_ASAP7_75t_L g1539 ( .A(n_38), .Y(n_1539) );
AOI221xp5_ASAP7_75t_SL g1556 ( .A1(n_38), .A2(n_170), .B1(n_530), .B2(n_690), .C(n_1557), .Y(n_1556) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_39), .A2(n_161), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_39), .A2(n_148), .B1(n_548), .B2(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g1211 ( .A(n_40), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_41), .A2(n_121), .B1(n_528), .B2(n_529), .C(n_530), .Y(n_527) );
INVx1_ASAP7_75t_L g572 ( .A(n_41), .Y(n_572) );
INVx1_ASAP7_75t_L g1533 ( .A(n_42), .Y(n_1533) );
AOI221xp5_ASAP7_75t_L g1564 ( .A1(n_42), .A2(n_159), .B1(n_686), .B2(n_1565), .C(n_1566), .Y(n_1564) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_43), .Y(n_500) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_44), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_44), .A2(n_168), .B1(n_905), .B2(n_906), .Y(n_904) );
OAI22xp33_ASAP7_75t_R g1265 ( .A1(n_45), .A2(n_259), .B1(n_347), .B2(n_696), .Y(n_1265) );
OAI221xp5_ASAP7_75t_L g1283 ( .A1(n_45), .A2(n_259), .B1(n_440), .B2(n_802), .C(n_862), .Y(n_1283) );
OAI221xp5_ASAP7_75t_SL g341 ( .A1(n_46), .A2(n_242), .B1(n_342), .B2(n_347), .C(n_351), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_46), .A2(n_242), .B1(n_440), .B2(n_447), .C(n_450), .Y(n_439) );
INVx1_ASAP7_75t_L g817 ( .A(n_47), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_48), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_49), .A2(n_157), .B1(n_376), .B2(n_379), .C(n_383), .Y(n_375) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_49), .Y(n_470) );
INVx1_ASAP7_75t_L g786 ( .A(n_50), .Y(n_786) );
INVx1_ASAP7_75t_L g763 ( .A(n_51), .Y(n_763) );
INVx1_ASAP7_75t_L g1275 ( .A(n_52), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g1530 ( .A(n_53), .Y(n_1530) );
INVx1_ASAP7_75t_L g1542 ( .A(n_54), .Y(n_1542) );
AOI22xp33_ASAP7_75t_L g1559 ( .A1(n_54), .A2(n_63), .B1(n_1560), .B2(n_1561), .Y(n_1559) );
INVx1_ASAP7_75t_L g1172 ( .A(n_55), .Y(n_1172) );
OAI22xp5_ASAP7_75t_L g1610 ( .A1(n_56), .A2(n_214), .B1(n_1017), .B2(n_1019), .Y(n_1610) );
AOI22xp33_ASAP7_75t_L g1619 ( .A1(n_56), .A2(n_214), .B1(n_759), .B2(n_1620), .Y(n_1619) );
INVx1_ASAP7_75t_L g1583 ( .A(n_57), .Y(n_1583) );
AOI221xp5_ASAP7_75t_SL g517 ( .A1(n_58), .A2(n_78), .B1(n_366), .B2(n_518), .C(n_520), .Y(n_517) );
INVx1_ASAP7_75t_L g550 ( .A(n_58), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_59), .A2(n_210), .B1(n_587), .B2(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1126 ( .A(n_59), .Y(n_1126) );
INVx1_ASAP7_75t_L g514 ( .A(n_60), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_61), .A2(n_127), .B1(n_534), .B2(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_62), .A2(n_79), .B1(n_687), .B2(n_948), .Y(n_947) );
INVxp67_ASAP7_75t_L g1000 ( .A(n_62), .Y(n_1000) );
INVx1_ASAP7_75t_L g1537 ( .A(n_63), .Y(n_1537) );
INVx1_ASAP7_75t_L g512 ( .A(n_64), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g675 ( .A(n_65), .Y(n_675) );
INVx1_ASAP7_75t_L g374 ( .A(n_66), .Y(n_374) );
INVxp33_ASAP7_75t_L g1222 ( .A(n_67), .Y(n_1222) );
NAND2xp33_ASAP7_75t_SL g1238 ( .A(n_67), .B(n_1239), .Y(n_1238) );
INVxp33_ASAP7_75t_SL g868 ( .A(n_68), .Y(n_868) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_68), .A2(n_235), .B1(n_901), .B2(n_902), .C(n_903), .Y(n_900) );
AOI221xp5_ASAP7_75t_L g1259 ( .A1(n_69), .A2(n_141), .B1(n_948), .B2(n_1188), .C(n_1260), .Y(n_1259) );
INVxp33_ASAP7_75t_L g1280 ( .A(n_69), .Y(n_1280) );
AOI22xp5_ASAP7_75t_L g1351 ( .A1(n_70), .A2(n_96), .B1(n_1329), .B2(n_1342), .Y(n_1351) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_71), .A2(n_213), .B1(n_651), .B2(n_652), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_71), .Y(n_716) );
INVxp33_ASAP7_75t_SL g1032 ( .A(n_72), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_72), .A2(n_267), .B1(n_1058), .B2(n_1064), .C(n_1066), .Y(n_1063) );
OAI221xp5_ASAP7_75t_L g1593 ( .A1(n_73), .A2(n_994), .B1(n_1594), .B2(n_1597), .C(n_1601), .Y(n_1593) );
AOI22xp33_ASAP7_75t_SL g1617 ( .A1(n_73), .A2(n_279), .B1(n_528), .B2(n_1618), .Y(n_1617) );
AOI22xp5_ASAP7_75t_SL g1347 ( .A1(n_75), .A2(n_92), .B1(n_1323), .B2(n_1329), .Y(n_1347) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_76), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_77), .A2(n_230), .B1(n_780), .B2(n_1157), .Y(n_1166) );
INVx1_ASAP7_75t_L g1181 ( .A(n_77), .Y(n_1181) );
INVx1_ASAP7_75t_L g547 ( .A(n_78), .Y(n_547) );
INVxp67_ASAP7_75t_L g997 ( .A(n_79), .Y(n_997) );
INVx1_ASAP7_75t_L g1246 ( .A(n_80), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1524 ( .A1(n_81), .A2(n_1525), .B1(n_1569), .B2(n_1570), .Y(n_1524) );
CKINVDCx5p33_ASAP7_75t_R g1569 ( .A(n_81), .Y(n_1569) );
XOR2x2_ASAP7_75t_L g582 ( .A(n_82), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g1152 ( .A(n_83), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1174 ( .A1(n_83), .A2(n_108), .B1(n_523), .B2(n_1058), .C(n_1175), .Y(n_1174) );
CKINVDCx16_ASAP7_75t_R g1327 ( .A(n_84), .Y(n_1327) );
INVx1_ASAP7_75t_L g1596 ( .A(n_85), .Y(n_1596) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_85), .A2(n_226), .B1(n_1614), .B2(n_1615), .Y(n_1613) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_86), .A2(n_249), .B1(n_891), .B2(n_1273), .Y(n_1272) );
INVxp67_ASAP7_75t_SL g1292 ( .A(n_86), .Y(n_1292) );
OAI221xp5_ASAP7_75t_L g504 ( .A1(n_87), .A2(n_232), .B1(n_505), .B2(n_507), .C(n_510), .Y(n_504) );
INVx1_ASAP7_75t_L g561 ( .A(n_87), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_88), .Y(n_1151) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_89), .A2(n_154), .B1(n_314), .B2(n_654), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g714 ( .A(n_89), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g1216 ( .A1(n_90), .A2(n_185), .B1(n_658), .B2(n_801), .C(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1242 ( .A(n_90), .Y(n_1242) );
AOI221xp5_ASAP7_75t_L g1087 ( .A1(n_91), .A2(n_255), .B1(n_389), .B2(n_1059), .C(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1115 ( .A(n_91), .Y(n_1115) );
OA22x2_ASAP7_75t_L g1249 ( .A1(n_93), .A2(n_1250), .B1(n_1251), .B2(n_1296), .Y(n_1249) );
CKINVDCx16_ASAP7_75t_R g1296 ( .A(n_93), .Y(n_1296) );
INVx1_ASAP7_75t_L g400 ( .A(n_94), .Y(n_400) );
INVx1_ASAP7_75t_L g323 ( .A(n_95), .Y(n_323) );
INVx1_ASAP7_75t_L g368 ( .A(n_95), .Y(n_368) );
AO221x2_ASAP7_75t_L g1352 ( .A1(n_97), .A2(n_265), .B1(n_1329), .B2(n_1342), .C(n_1353), .Y(n_1352) );
CKINVDCx5p33_ASAP7_75t_R g1254 ( .A(n_98), .Y(n_1254) );
CKINVDCx5p33_ASAP7_75t_R g1548 ( .A(n_99), .Y(n_1548) );
INVx1_ASAP7_75t_L g935 ( .A(n_100), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_101), .A2(n_278), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g767 ( .A(n_101), .Y(n_767) );
INVx1_ASAP7_75t_L g511 ( .A(n_102), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_102), .A2(n_232), .B1(n_556), .B2(n_558), .C(n_560), .Y(n_555) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_103), .Y(n_809) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_103), .A2(n_222), .B1(n_378), .B2(n_528), .C(n_530), .Y(n_832) );
INVxp33_ASAP7_75t_SL g795 ( .A(n_104), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_104), .A2(n_120), .B1(n_529), .B2(n_841), .Y(n_840) );
INVxp33_ASAP7_75t_L g1220 ( .A(n_105), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1373 ( .A1(n_106), .A2(n_252), .B1(n_1336), .B2(n_1374), .Y(n_1373) );
CKINVDCx20_ASAP7_75t_R g1421 ( .A(n_107), .Y(n_1421) );
INVx1_ASAP7_75t_L g1147 ( .A(n_108), .Y(n_1147) );
OAI211xp5_ASAP7_75t_L g622 ( .A1(n_109), .A2(n_623), .B(n_625), .C(n_627), .Y(n_622) );
INVxp33_ASAP7_75t_SL g859 ( .A(n_110), .Y(n_859) );
INVx1_ASAP7_75t_L g537 ( .A(n_111), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g1534 ( .A1(n_112), .A2(n_142), .B1(n_657), .B2(n_658), .C(n_801), .Y(n_1534) );
OAI22xp5_ASAP7_75t_L g1563 ( .A1(n_112), .A2(n_142), .B1(n_696), .B2(n_697), .Y(n_1563) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_113), .Y(n_1090) );
INVxp33_ASAP7_75t_SL g925 ( .A(n_114), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_114), .A2(n_163), .B1(n_780), .B2(n_984), .C(n_986), .Y(n_983) );
INVx1_ASAP7_75t_L g813 ( .A(n_115), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_115), .A2(n_184), .B1(n_704), .B2(n_834), .Y(n_833) );
OAI22xp33_ASAP7_75t_SL g1106 ( .A1(n_116), .A2(n_224), .B1(n_588), .B2(n_742), .Y(n_1106) );
INVx1_ASAP7_75t_L g1130 ( .A(n_116), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_117), .A2(n_175), .B1(n_388), .B2(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g474 ( .A(n_117), .Y(n_474) );
INVx1_ASAP7_75t_L g287 ( .A(n_118), .Y(n_287) );
INVx1_ASAP7_75t_L g1212 ( .A(n_119), .Y(n_1212) );
INVxp33_ASAP7_75t_SL g799 ( .A(n_120), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_122), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_123), .A2(n_199), .B1(n_950), .B2(n_951), .Y(n_949) );
INVxp67_ASAP7_75t_SL g1011 ( .A(n_123), .Y(n_1011) );
INVx1_ASAP7_75t_L g1047 ( .A(n_124), .Y(n_1047) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_124), .A2(n_220), .B1(n_1058), .B2(n_1059), .C(n_1061), .Y(n_1057) );
AOI221xp5_ASAP7_75t_L g1094 ( .A1(n_125), .A2(n_166), .B1(n_608), .B2(n_957), .C(n_1095), .Y(n_1094) );
INVx1_ASAP7_75t_L g1134 ( .A(n_125), .Y(n_1134) );
INVx1_ASAP7_75t_L g750 ( .A(n_126), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_126), .A2(n_176), .B1(n_778), .B2(n_780), .Y(n_777) );
INVxp33_ASAP7_75t_SL g858 ( .A(n_127), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g1097 ( .A(n_128), .Y(n_1097) );
AOI221xp5_ASAP7_75t_L g1268 ( .A1(n_129), .A2(n_223), .B1(n_608), .B2(n_1269), .C(n_1271), .Y(n_1268) );
INVxp67_ASAP7_75t_SL g1287 ( .A(n_129), .Y(n_1287) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_130), .A2(n_156), .B1(n_1161), .B2(n_1163), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g1182 ( .A1(n_130), .A2(n_218), .B1(n_385), .B2(n_608), .C(n_1183), .Y(n_1182) );
AOI22xp5_ASAP7_75t_L g1346 ( .A1(n_131), .A2(n_240), .B1(n_1336), .B2(n_1339), .Y(n_1346) );
INVx1_ASAP7_75t_L g1074 ( .A(n_132), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_133), .A2(n_256), .B1(n_757), .B2(n_759), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_133), .A2(n_149), .B1(n_772), .B2(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g788 ( .A(n_134), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g656 ( .A1(n_135), .A2(n_237), .B1(n_440), .B2(n_657), .C(n_658), .Y(n_656) );
OAI222xp33_ASAP7_75t_L g695 ( .A1(n_135), .A2(n_154), .B1(n_237), .B2(n_536), .C1(n_696), .C2(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g1214 ( .A(n_136), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1375 ( .A1(n_137), .A2(n_138), .B1(n_1323), .B2(n_1376), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_137), .A2(n_1575), .B1(n_1577), .B2(n_1622), .Y(n_1574) );
XOR2xp5_ASAP7_75t_L g1578 ( .A(n_137), .B(n_1579), .Y(n_1578) );
AOI21xp33_ASAP7_75t_L g607 ( .A1(n_139), .A2(n_608), .B(n_610), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g1553 ( .A(n_140), .Y(n_1553) );
INVxp33_ASAP7_75t_L g1282 ( .A(n_141), .Y(n_1282) );
CKINVDCx14_ASAP7_75t_R g1355 ( .A(n_143), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_144), .A2(n_218), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_144), .A2(n_156), .B1(n_1187), .B2(n_1188), .Y(n_1186) );
AOI22xp5_ASAP7_75t_L g1335 ( .A1(n_145), .A2(n_243), .B1(n_1336), .B2(n_1339), .Y(n_1335) );
INVx1_ASAP7_75t_L g1604 ( .A(n_146), .Y(n_1604) );
INVx1_ASAP7_75t_L g1588 ( .A(n_147), .Y(n_1588) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_148), .A2(n_164), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_149), .A2(n_158), .B1(n_385), .B2(n_752), .C(n_754), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_150), .A2(n_229), .B1(n_429), .B2(n_1055), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_150), .A2(n_251), .B1(n_587), .B2(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1587 ( .A(n_151), .Y(n_1587) );
INVxp33_ASAP7_75t_L g796 ( .A(n_152), .Y(n_796) );
INVx1_ASAP7_75t_L g1584 ( .A(n_153), .Y(n_1584) );
CKINVDCx5p33_ASAP7_75t_R g1550 ( .A(n_155), .Y(n_1550) );
INVx1_ASAP7_75t_L g465 ( .A(n_157), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_158), .A2(n_256), .B1(n_548), .B2(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g1529 ( .A(n_159), .Y(n_1529) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_160), .A2(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g628 ( .A(n_160), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_161), .A2(n_164), .B1(n_414), .B2(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g762 ( .A(n_162), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_162), .A2(n_196), .B1(n_772), .B2(n_775), .Y(n_774) );
INVxp33_ASAP7_75t_SL g921 ( .A(n_163), .Y(n_921) );
AOI22xp33_ASAP7_75t_SL g952 ( .A1(n_165), .A2(n_177), .B1(n_951), .B2(n_953), .Y(n_952) );
OAI211xp5_ASAP7_75t_SL g973 ( .A1(n_165), .A2(n_974), .B(n_979), .C(n_988), .Y(n_973) );
INVx1_ASAP7_75t_L g1136 ( .A(n_166), .Y(n_1136) );
XNOR2xp5_ASAP7_75t_L g912 ( .A(n_167), .B(n_913), .Y(n_912) );
INVxp67_ASAP7_75t_SL g871 ( .A(n_168), .Y(n_871) );
OAI221xp5_ASAP7_75t_L g800 ( .A1(n_169), .A2(n_280), .B1(n_447), .B2(n_801), .C(n_802), .Y(n_800) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_169), .A2(n_280), .B1(n_342), .B2(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g1541 ( .A(n_170), .Y(n_1541) );
INVx1_ASAP7_75t_L g1598 ( .A(n_171), .Y(n_1598) );
AOI22xp33_ASAP7_75t_L g1612 ( .A1(n_171), .A2(n_203), .B1(n_388), .B2(n_1270), .Y(n_1612) );
INVxp33_ASAP7_75t_L g1208 ( .A(n_172), .Y(n_1208) );
INVx1_ASAP7_75t_L g1040 ( .A(n_173), .Y(n_1040) );
INVx1_ASAP7_75t_L g352 ( .A(n_174), .Y(n_352) );
INVx1_ASAP7_75t_L g459 ( .A(n_175), .Y(n_459) );
INVx1_ASAP7_75t_L g761 ( .A(n_176), .Y(n_761) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_177), .A2(n_994), .B1(n_996), .B2(n_1006), .C(n_1014), .Y(n_993) );
INVx1_ASAP7_75t_L g1169 ( .A(n_178), .Y(n_1169) );
INVx1_ASAP7_75t_L g1264 ( .A(n_179), .Y(n_1264) );
INVx1_ASAP7_75t_L g790 ( .A(n_180), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_181), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_182), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_182), .B(n_287), .Y(n_1310) );
AND3x2_ASAP7_75t_L g1326 ( .A(n_182), .B(n_287), .C(n_1313), .Y(n_1326) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_183), .Y(n_602) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_184), .Y(n_808) );
INVx1_ASAP7_75t_L g1243 ( .A(n_185), .Y(n_1243) );
AOI22xp5_ASAP7_75t_SL g1362 ( .A1(n_186), .A2(n_201), .B1(n_1323), .B2(n_1329), .Y(n_1362) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_187), .A2(n_228), .B1(n_591), .B2(n_597), .C(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g626 ( .A(n_187), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_188), .Y(n_670) );
INVx2_ASAP7_75t_L g300 ( .A(n_189), .Y(n_300) );
INVx1_ASAP7_75t_L g515 ( .A(n_190), .Y(n_515) );
XNOR2x2_ASAP7_75t_L g1028 ( .A(n_191), .B(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1257 ( .A(n_192), .Y(n_1257) );
INVx1_ASAP7_75t_L g641 ( .A(n_193), .Y(n_641) );
INVx1_ASAP7_75t_L g878 ( .A(n_194), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_195), .Y(n_677) );
INVx1_ASAP7_75t_L g733 ( .A(n_196), .Y(n_733) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_197), .Y(n_1149) );
AOI22xp5_ASAP7_75t_SL g1361 ( .A1(n_198), .A2(n_258), .B1(n_1336), .B2(n_1339), .Y(n_1361) );
INVxp67_ASAP7_75t_SL g1008 ( .A(n_199), .Y(n_1008) );
INVx1_ASAP7_75t_L g849 ( .A(n_200), .Y(n_849) );
INVx1_ASAP7_75t_L g1313 ( .A(n_202), .Y(n_1313) );
INVx1_ASAP7_75t_L g1599 ( .A(n_203), .Y(n_1599) );
INVx1_ASAP7_75t_L g1043 ( .A(n_204), .Y(n_1043) );
INVx1_ASAP7_75t_L g1034 ( .A(n_205), .Y(n_1034) );
INVx1_ASAP7_75t_L g1144 ( .A(n_206), .Y(n_1144) );
INVx1_ASAP7_75t_L g1267 ( .A(n_207), .Y(n_1267) );
AOI22x1_ASAP7_75t_L g1198 ( .A1(n_208), .A2(n_1199), .B1(n_1200), .B2(n_1247), .Y(n_1198) );
INVx1_ASAP7_75t_L g1247 ( .A(n_208), .Y(n_1247) );
AO221x2_ASAP7_75t_L g1418 ( .A1(n_208), .A2(n_281), .B1(n_1376), .B2(n_1419), .C(n_1420), .Y(n_1418) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_209), .Y(n_661) );
INVx1_ASAP7_75t_L g1128 ( .A(n_210), .Y(n_1128) );
INVx1_ASAP7_75t_L g1262 ( .A(n_211), .Y(n_1262) );
INVx1_ASAP7_75t_L g820 ( .A(n_212), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_213), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_215), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g1111 ( .A(n_216), .Y(n_1111) );
INVx1_ASAP7_75t_L g302 ( .A(n_217), .Y(n_302) );
INVx2_ASAP7_75t_L g421 ( .A(n_217), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g1110 ( .A(n_219), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_220), .A2(n_225), .B1(n_551), .B2(n_1049), .Y(n_1048) );
CKINVDCx14_ASAP7_75t_R g1423 ( .A(n_221), .Y(n_1423) );
INVxp67_ASAP7_75t_SL g812 ( .A(n_222), .Y(n_812) );
INVxp67_ASAP7_75t_SL g1291 ( .A(n_223), .Y(n_1291) );
INVx1_ASAP7_75t_L g1123 ( .A(n_224), .Y(n_1123) );
INVx1_ASAP7_75t_L g1062 ( .A(n_225), .Y(n_1062) );
INVx1_ASAP7_75t_L g1595 ( .A(n_226), .Y(n_1595) );
XOR2x1_ASAP7_75t_L g1139 ( .A(n_227), .B(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g646 ( .A(n_228), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g1078 ( .A1(n_229), .A2(n_261), .B1(n_591), .B2(n_740), .Y(n_1078) );
INVx1_ASAP7_75t_L g1191 ( .A(n_230), .Y(n_1191) );
INVxp33_ASAP7_75t_L g1207 ( .A(n_231), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_233), .A2(n_250), .B1(n_523), .B2(n_524), .Y(n_522) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_233), .A2(n_250), .B1(n_544), .B2(n_545), .C(n_546), .Y(n_543) );
INVx1_ASAP7_75t_L g818 ( .A(n_234), .Y(n_818) );
INVxp67_ASAP7_75t_SL g870 ( .A(n_235), .Y(n_870) );
INVx1_ASAP7_75t_L g879 ( .A(n_236), .Y(n_879) );
CKINVDCx16_ASAP7_75t_R g1320 ( .A(n_238), .Y(n_1320) );
INVx1_ASAP7_75t_L g930 ( .A(n_239), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_241), .Y(n_667) );
INVx1_ASAP7_75t_L g1314 ( .A(n_245), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_245), .B(n_1312), .Y(n_1319) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_247), .A2(n_364), .B(n_366), .Y(n_363) );
INVxp33_ASAP7_75t_L g427 ( .A(n_247), .Y(n_427) );
INVxp33_ASAP7_75t_L g432 ( .A(n_248), .Y(n_432) );
INVxp67_ASAP7_75t_SL g1286 ( .A(n_249), .Y(n_1286) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_251), .Y(n_1053) );
INVx1_ASAP7_75t_L g941 ( .A(n_253), .Y(n_941) );
INVx1_ASAP7_75t_L g1591 ( .A(n_254), .Y(n_1591) );
INVx1_ASAP7_75t_L g1121 ( .A(n_255), .Y(n_1121) );
INVx1_ASAP7_75t_L g1276 ( .A(n_257), .Y(n_1276) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_260), .A2(n_364), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g785 ( .A(n_260), .Y(n_785) );
INVxp67_ASAP7_75t_SL g1052 ( .A(n_261), .Y(n_1052) );
INVx1_ASAP7_75t_L g1215 ( .A(n_262), .Y(n_1215) );
INVx2_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_264), .Y(n_965) );
XNOR2x2_ASAP7_75t_L g1084 ( .A(n_266), .B(n_1085), .Y(n_1084) );
INVxp33_ASAP7_75t_SL g1036 ( .A(n_267), .Y(n_1036) );
INVx1_ASAP7_75t_L g396 ( .A(n_268), .Y(n_396) );
INVx1_ASAP7_75t_L g1038 ( .A(n_269), .Y(n_1038) );
CKINVDCx20_ASAP7_75t_R g1315 ( .A(n_270), .Y(n_1315) );
INVx1_ASAP7_75t_L g821 ( .A(n_271), .Y(n_821) );
BUFx3_ASAP7_75t_L g328 ( .A(n_272), .Y(n_328) );
INVx1_ASAP7_75t_L g357 ( .A(n_272), .Y(n_357) );
BUFx3_ASAP7_75t_L g330 ( .A(n_273), .Y(n_330) );
INVx1_ASAP7_75t_L g337 ( .A(n_273), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_274), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_275), .Y(n_1091) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_276), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g744 ( .A(n_277), .Y(n_744) );
INVx1_ASAP7_75t_L g766 ( .A(n_278), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g1602 ( .A1(n_279), .A2(n_974), .B1(n_1603), .B2(n_1606), .C(n_1608), .Y(n_1602) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_303), .B(n_1299), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
AND2x4_ASAP7_75t_L g1576 ( .A(n_285), .B(n_291), .Y(n_1576) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_SL g1573 ( .A(n_286), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1626 ( .A(n_286), .B(n_288), .Y(n_1626) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_288), .B(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g564 ( .A(n_294), .B(n_302), .Y(n_564) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g454 ( .A(n_295), .B(n_455), .Y(n_454) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
OR2x2_ASAP7_75t_L g314 ( .A(n_297), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g458 ( .A(n_297), .Y(n_458) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_297), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_297), .A2(n_602), .B1(n_641), .B2(n_642), .Y(n_640) );
INVx2_ASAP7_75t_SL g866 ( .A(n_297), .Y(n_866) );
INVx2_ASAP7_75t_SL g1010 ( .A(n_297), .Y(n_1010) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x4_ASAP7_75t_L g416 ( .A(n_299), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g425 ( .A(n_299), .Y(n_425) );
AND2x2_ASAP7_75t_L g431 ( .A(n_299), .B(n_300), .Y(n_431) );
INVx2_ASAP7_75t_L g436 ( .A(n_299), .Y(n_436) );
INVx1_ASAP7_75t_L g464 ( .A(n_299), .Y(n_464) );
INVx2_ASAP7_75t_L g417 ( .A(n_300), .Y(n_417) );
INVx1_ASAP7_75t_L g438 ( .A(n_300), .Y(n_438) );
INVx1_ASAP7_75t_L g445 ( .A(n_300), .Y(n_445) );
INVx1_ASAP7_75t_L g463 ( .A(n_300), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_300), .B(n_436), .Y(n_469) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_1023), .B1(n_1024), .B2(n_1298), .Y(n_303) );
INVx1_ASAP7_75t_L g1298 ( .A(n_304), .Y(n_1298) );
AO22x1_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_725), .B2(n_726), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
XNOR2x1_ASAP7_75t_L g307 ( .A(n_308), .B(n_496), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
XNOR2x1_ASAP7_75t_L g309 ( .A(n_310), .B(n_495), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_408), .Y(n_310) );
AOI21xp33_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_331), .B(n_332), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_312), .A2(n_405), .B1(n_731), .B2(n_763), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g1226 ( .A1(n_312), .A2(n_1227), .B1(n_1228), .B2(n_1246), .Y(n_1226) );
INVx5_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g846 ( .A(n_313), .Y(n_846) );
INVx1_ASAP7_75t_L g1168 ( .A(n_313), .Y(n_1168) );
INVx2_ASAP7_75t_L g1253 ( .A(n_313), .Y(n_1253) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
INVx2_ASAP7_75t_L g573 ( .A(n_314), .Y(n_573) );
INVx3_ASAP7_75t_L g446 ( .A(n_315), .Y(n_446) );
INVx1_ASAP7_75t_L g971 ( .A(n_316), .Y(n_971) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x6_ASAP7_75t_L g966 ( .A(n_318), .B(n_967), .Y(n_966) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x4_ASAP7_75t_L g959 ( .A(n_319), .B(n_367), .Y(n_959) );
INVx2_ASAP7_75t_L g536 ( .A(n_320), .Y(n_536) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_326), .Y(n_320) );
AND2x4_ASAP7_75t_L g343 ( .A(n_321), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g348 ( .A(n_321), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g393 ( .A(n_321), .Y(n_393) );
AND2x4_ASAP7_75t_L g513 ( .A(n_321), .B(n_344), .Y(n_513) );
BUFx2_ASAP7_75t_L g600 ( .A(n_321), .Y(n_600) );
AND2x2_ASAP7_75t_L g737 ( .A(n_321), .B(n_349), .Y(n_737) );
AND2x4_ASAP7_75t_L g844 ( .A(n_321), .B(n_349), .Y(n_844) );
NAND2x1p5_ASAP7_75t_L g940 ( .A(n_321), .B(n_491), .Y(n_940) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g367 ( .A(n_324), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g386 ( .A(n_325), .B(n_368), .Y(n_386) );
INVx6_ASAP7_75t_L g365 ( .A(n_326), .Y(n_365) );
BUFx2_ASAP7_75t_L g620 ( .A(n_326), .Y(n_620) );
INVx2_ASAP7_75t_L g928 ( .A(n_326), .Y(n_928) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g350 ( .A(n_327), .Y(n_350) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g336 ( .A(n_328), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g373 ( .A(n_328), .B(n_330), .Y(n_373) );
INVx1_ASAP7_75t_L g346 ( .A(n_329), .Y(n_346) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g362 ( .A(n_330), .B(n_357), .Y(n_362) );
AOI31xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_369), .A3(n_395), .B(n_404), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_340), .B(n_341), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_334), .A2(n_397), .B1(n_761), .B2(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g896 ( .A(n_334), .Y(n_896) );
AOI211xp5_ASAP7_75t_L g1171 ( .A1(n_334), .A2(n_1172), .B(n_1173), .C(n_1174), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_334), .A2(n_397), .B1(n_1211), .B2(n_1214), .Y(n_1244) );
HB1xp67_ASAP7_75t_L g1258 ( .A(n_334), .Y(n_1258) );
AOI211xp5_ASAP7_75t_L g1562 ( .A1(n_334), .A2(n_1547), .B(n_1563), .C(n_1564), .Y(n_1562) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
BUFx3_ASAP7_75t_L g523 ( .A(n_335), .Y(n_523) );
INVx2_ASAP7_75t_SL g956 ( .A(n_335), .Y(n_956) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_336), .Y(n_360) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
BUFx2_ASAP7_75t_L g529 ( .A(n_336), .Y(n_529) );
INVx2_ASAP7_75t_SL g609 ( .A(n_336), .Y(n_609) );
BUFx3_ASAP7_75t_L g618 ( .A(n_336), .Y(n_618) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_336), .Y(n_710) );
BUFx2_ASAP7_75t_L g901 ( .A(n_336), .Y(n_901) );
INVx1_ASAP7_75t_L g358 ( .A(n_337), .Y(n_358) );
AND2x4_ASAP7_75t_L g371 ( .A(n_338), .B(n_372), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g503 ( .A1(n_338), .A2(n_348), .B1(n_504), .B2(n_513), .C1(n_514), .C2(n_515), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g585 ( .A1(n_338), .A2(n_586), .B(n_589), .Y(n_585) );
AND2x2_ASAP7_75t_L g830 ( .A(n_338), .B(n_378), .Y(n_830) );
OAI21xp5_ASAP7_75t_L g1075 ( .A1(n_338), .A2(n_1076), .B(n_1078), .Y(n_1075) );
OAI21xp33_ASAP7_75t_L g1103 ( .A1(n_338), .A2(n_1104), .B(n_1106), .Y(n_1103) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g398 ( .A(n_339), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g402 ( .A(n_339), .B(n_403), .Y(n_402) );
A2O1A1Ixp33_ASAP7_75t_SL g683 ( .A1(n_339), .A2(n_684), .B(n_689), .C(n_694), .Y(n_683) );
OR2x2_ASAP7_75t_L g920 ( .A(n_339), .B(n_419), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_340), .A2(n_400), .B1(n_476), .B2(n_479), .Y(n_475) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx4_ASAP7_75t_L g1109 ( .A(n_343), .Y(n_1109) );
INVxp67_ASAP7_75t_L g597 ( .A(n_344), .Y(n_597) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g938 ( .A(n_345), .Y(n_938) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_348), .A2(n_513), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
INVx1_ASAP7_75t_L g598 ( .A(n_349), .Y(n_598) );
INVx2_ASAP7_75t_L g698 ( .A(n_349), .Y(n_698) );
BUFx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI211xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B(n_359), .C(n_363), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_352), .A2(n_411), .B1(n_412), .B2(n_422), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_353), .A2(n_1034), .B1(n_1040), .B2(n_1067), .C(n_1069), .Y(n_1066) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_SL g591 ( .A(n_354), .Y(n_591) );
INVx1_ASAP7_75t_L g1176 ( .A(n_354), .Y(n_1176) );
INVx1_ASAP7_75t_L g1261 ( .A(n_354), .Y(n_1261) );
BUFx4f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g604 ( .A(n_355), .Y(n_604) );
INVx1_ASAP7_75t_L g707 ( .A(n_355), .Y(n_707) );
BUFx2_ASAP7_75t_L g743 ( .A(n_355), .Y(n_743) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
OR2x2_ASAP7_75t_L g399 ( .A(n_356), .B(n_358), .Y(n_399) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g740 ( .A(n_360), .Y(n_740) );
INVx1_ASAP7_75t_L g1065 ( .A(n_360), .Y(n_1065) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_361), .Y(n_704) );
BUFx3_ASAP7_75t_L g957 ( .A(n_361), .Y(n_957) );
INVx1_ASAP7_75t_L g1105 ( .A(n_361), .Y(n_1105) );
INVx1_ASAP7_75t_L g1616 ( .A(n_361), .Y(n_1616) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
INVx2_ASAP7_75t_L g403 ( .A(n_362), .Y(n_403) );
INVx1_ASAP7_75t_L g525 ( .A(n_362), .Y(n_525) );
INVx1_ASAP7_75t_L g688 ( .A(n_362), .Y(n_688) );
BUFx3_ASAP7_75t_L g388 ( .A(n_364), .Y(n_388) );
HB1xp67_ASAP7_75t_L g1560 ( .A(n_364), .Y(n_1560) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g521 ( .A(n_365), .Y(n_521) );
INVx1_ASAP7_75t_L g533 ( .A(n_365), .Y(n_533) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_365), .Y(n_595) );
INVx1_ASAP7_75t_L g606 ( .A(n_365), .Y(n_606) );
INVx2_ASAP7_75t_SL g836 ( .A(n_365), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g621 ( .A(n_367), .Y(n_621) );
INVx2_ASAP7_75t_L g746 ( .A(n_367), .Y(n_746) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_367), .Y(n_1069) );
INVx2_ASAP7_75t_SL g1099 ( .A(n_367), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_374), .B1(n_375), .B2(n_387), .C(n_391), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_370), .A2(n_391), .B1(n_1551), .B2(n_1556), .C(n_1559), .Y(n_1555) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_SL g749 ( .A(n_371), .Y(n_749) );
INVx1_ASAP7_75t_L g908 ( .A(n_371), .Y(n_908) );
INVx1_ASAP7_75t_L g1180 ( .A(n_371), .Y(n_1180) );
INVx1_ASAP7_75t_L g1231 ( .A(n_371), .Y(n_1231) );
INVx2_ASAP7_75t_SL g519 ( .A(n_372), .Y(n_519) );
BUFx3_ASAP7_75t_L g528 ( .A(n_372), .Y(n_528) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_372), .Y(n_693) );
BUFx4f_ASAP7_75t_L g1270 ( .A(n_372), .Y(n_1270) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_373), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_374), .A2(n_396), .B1(n_483), .B2(n_486), .Y(n_482) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_378), .A2(n_394), .B1(n_511), .B2(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g588 ( .A(n_378), .Y(n_588) );
BUFx2_ASAP7_75t_L g894 ( .A(n_378), .Y(n_894) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_380), .B(n_963), .Y(n_1585) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_382), .Y(n_394) );
INVx2_ASAP7_75t_L g890 ( .A(n_382), .Y(n_890) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g1061 ( .A1(n_384), .A2(n_742), .B1(n_753), .B2(n_1043), .C(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g1271 ( .A(n_385), .Y(n_1271) );
INVx2_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g531 ( .A(n_386), .Y(n_531) );
INVx2_ASAP7_75t_L g612 ( .A(n_386), .Y(n_612) );
INVx1_ASAP7_75t_L g1093 ( .A(n_386), .Y(n_1093) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g590 ( .A(n_390), .Y(n_590) );
BUFx6f_ASAP7_75t_L g1058 ( .A(n_390), .Y(n_1058) );
INVx1_ASAP7_75t_L g1237 ( .A(n_390), .Y(n_1237) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_391), .A2(n_517), .B(n_522), .Y(n_516) );
INVx1_ASAP7_75t_L g694 ( .A(n_391), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_391), .A2(n_748), .B1(n_750), .B2(n_751), .C(n_756), .Y(n_747) );
AOI221xp5_ASAP7_75t_L g831 ( .A1(n_391), .A2(n_748), .B1(n_821), .B2(n_832), .C(n_833), .Y(n_831) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_391), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_391), .A2(n_1179), .B1(n_1181), .B2(n_1182), .C(n_1186), .Y(n_1178) );
AOI221xp5_ASAP7_75t_L g1229 ( .A1(n_391), .A2(n_1212), .B1(n_1230), .B2(n_1232), .C(n_1233), .Y(n_1229) );
AOI221xp5_ASAP7_75t_L g1266 ( .A1(n_391), .A2(n_1230), .B1(n_1267), .B2(n_1268), .C(n_1272), .Y(n_1266) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g697 ( .A(n_393), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g755 ( .A(n_394), .Y(n_755) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_394), .Y(n_839) );
INVx1_ASAP7_75t_L g1558 ( .A(n_394), .Y(n_1558) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_400), .B2(n_401), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_397), .A2(n_817), .B1(n_820), .B2(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_397), .A2(n_401), .B1(n_876), .B2(n_878), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_397), .A2(n_401), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_397), .A2(n_401), .B1(n_1275), .B2(n_1276), .Y(n_1274) );
AOI22xp33_ASAP7_75t_SL g1568 ( .A1(n_397), .A2(n_401), .B1(n_1548), .B2(n_1550), .Y(n_1568) );
INVx6_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g506 ( .A(n_399), .Y(n_506) );
INVx1_ASAP7_75t_L g1068 ( .A(n_399), .Y(n_1068) );
BUFx2_ASAP7_75t_L g1263 ( .A(n_399), .Y(n_1263) );
AOI211xp5_ASAP7_75t_L g732 ( .A1(n_401), .A2(n_733), .B(n_734), .C(n_738), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_401), .A2(n_818), .B1(n_838), .B2(n_840), .C(n_842), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_401), .B(n_1215), .Y(n_1245) );
INVx4_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g509 ( .A(n_403), .Y(n_509) );
INVx1_ASAP7_75t_L g841 ( .A(n_403), .Y(n_841) );
AOI31xp33_ASAP7_75t_L g1554 ( .A1(n_404), .A2(n_1555), .A3(n_1562), .B(n_1568), .Y(n_1554) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI31xp33_ASAP7_75t_SL g1086 ( .A1(n_405), .A2(n_1087), .A3(n_1094), .B(n_1100), .Y(n_1086) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g825 ( .A(n_406), .Y(n_825) );
BUFx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x6_ASAP7_75t_L g453 ( .A(n_407), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g540 ( .A(n_407), .Y(n_540) );
NOR3xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_439), .C(n_452), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_426), .Y(n_409) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g783 ( .A(n_413), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_413), .A2(n_858), .B1(n_859), .B2(n_860), .Y(n_857) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_413), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_413), .A2(n_422), .B1(n_1096), .B2(n_1134), .Y(n_1133) );
BUFx2_ASAP7_75t_L g1148 ( .A(n_413), .Y(n_1148) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_413), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_413), .A2(n_860), .B1(n_1262), .B2(n_1282), .Y(n_1281) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_418), .Y(n_413) );
BUFx3_ASAP7_75t_L g773 ( .A(n_414), .Y(n_773) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g481 ( .A(n_415), .Y(n_481) );
BUFx6f_ASAP7_75t_L g1046 ( .A(n_415), .Y(n_1046) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_416), .Y(n_473) );
INVx1_ASAP7_75t_L g1005 ( .A(n_416), .Y(n_1005) );
AND2x4_ASAP7_75t_L g424 ( .A(n_417), .B(n_425), .Y(n_424) );
AND2x6_ASAP7_75t_L g422 ( .A(n_418), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g428 ( .A(n_418), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g433 ( .A(n_418), .B(n_434), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_418), .A2(n_543), .B1(n_554), .B2(n_555), .Y(n_542) );
AND2x2_ASAP7_75t_L g624 ( .A(n_418), .B(n_434), .Y(n_624) );
AND2x2_ASAP7_75t_L g629 ( .A(n_418), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g632 ( .A(n_418), .B(n_481), .Y(n_632) );
AND2x2_ASAP7_75t_L g644 ( .A(n_418), .B(n_638), .Y(n_644) );
AND2x2_ASAP7_75t_L g787 ( .A(n_418), .B(n_434), .Y(n_787) );
AND2x2_ASAP7_75t_L g856 ( .A(n_418), .B(n_434), .Y(n_856) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_418), .B(n_434), .Y(n_1037) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
INVx2_ASAP7_75t_L g977 ( .A(n_420), .Y(n_977) );
AND2x4_ASAP7_75t_L g995 ( .A(n_420), .B(n_549), .Y(n_995) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_420), .B(n_435), .Y(n_1018) );
INVx1_ASAP7_75t_L g455 ( .A(n_421), .Y(n_455) );
INVx1_ASAP7_75t_L g493 ( .A(n_421), .Y(n_493) );
INVx1_ASAP7_75t_SL g652 ( .A(n_422), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_422), .A2(n_744), .B1(n_782), .B2(n_783), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_422), .A2(n_783), .B1(n_795), .B2(n_796), .Y(n_794) );
BUFx2_ASAP7_75t_L g860 ( .A(n_422), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_422), .A2(n_1032), .B1(n_1033), .B2(n_1034), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_422), .A2(n_1147), .B1(n_1148), .B2(n_1149), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_422), .A2(n_1220), .B1(n_1221), .B2(n_1222), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1528 ( .A1(n_422), .A2(n_1033), .B1(n_1529), .B2(n_1530), .Y(n_1528) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_423), .B(n_446), .Y(n_451) );
BUFx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_424), .Y(n_553) );
BUFx2_ASAP7_75t_L g581 ( .A(n_424), .Y(n_581) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_424), .Y(n_638) );
BUFx3_ASAP7_75t_L g978 ( .A(n_424), .Y(n_978) );
INVx1_ASAP7_75t_L g1159 ( .A(n_424), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_432), .B2(n_433), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_428), .A2(n_785), .B1(n_786), .B2(n_787), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_428), .A2(n_787), .B1(n_798), .B2(n_799), .Y(n_797) );
BUFx2_ASAP7_75t_L g854 ( .A(n_428), .Y(n_854) );
AOI21xp5_ASAP7_75t_L g1039 ( .A1(n_428), .A2(n_1040), .B(n_1041), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_428), .A2(n_433), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_428), .A2(n_787), .B1(n_1224), .B2(n_1225), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_428), .A2(n_856), .B1(n_1532), .B2(n_1533), .Y(n_1531) );
INVx2_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g630 ( .A(n_430), .Y(n_630) );
INVx2_ASAP7_75t_L g779 ( .A(n_430), .Y(n_779) );
INVx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_431), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g1135 ( .A1(n_433), .A2(n_573), .B1(n_1102), .B2(n_1136), .Y(n_1135) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g557 ( .A(n_435), .Y(n_557) );
INVx1_ASAP7_75t_L g567 ( .A(n_435), .Y(n_567) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_435), .Y(n_636) );
BUFx2_ASAP7_75t_L g772 ( .A(n_435), .Y(n_772) );
BUFx6f_ASAP7_75t_L g1162 ( .A(n_435), .Y(n_1162) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g449 ( .A(n_436), .Y(n_449) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_SL g801 ( .A(n_441), .Y(n_801) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2x1_ASAP7_75t_SL g442 ( .A(n_443), .B(n_446), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_445), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_446), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g575 ( .A(n_446), .B(n_576), .Y(n_575) );
AND2x4_ASAP7_75t_L g577 ( .A(n_446), .B(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g580 ( .A(n_446), .B(n_581), .Y(n_580) );
BUFx4f_ASAP7_75t_L g657 ( .A(n_447), .Y(n_657) );
BUFx4f_ASAP7_75t_L g1217 ( .A(n_447), .Y(n_1217) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x6_ASAP7_75t_L g992 ( .A(n_449), .B(n_970), .Y(n_992) );
BUFx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx3_ASAP7_75t_L g658 ( .A(n_451), .Y(n_658) );
BUFx2_ASAP7_75t_L g802 ( .A(n_451), .Y(n_802) );
OAI33xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_456), .A3(n_466), .B1(n_475), .B2(n_482), .B3(n_488), .Y(n_452) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_453), .Y(n_804) );
OAI33xp33_ASAP7_75t_L g863 ( .A1(n_453), .A2(n_864), .A3(n_869), .B1(n_873), .B2(n_877), .B3(n_880), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_453), .A2(n_488), .B1(n_1042), .B2(n_1051), .Y(n_1041) );
OAI33xp33_ASAP7_75t_L g1113 ( .A1(n_453), .A2(n_1114), .A3(n_1118), .B1(n_1122), .B2(n_1127), .B3(n_1131), .Y(n_1113) );
OAI33xp33_ASAP7_75t_L g1202 ( .A1(n_453), .A2(n_488), .A3(n_1203), .B1(n_1206), .B2(n_1210), .B3(n_1213), .Y(n_1202) );
OAI33xp33_ASAP7_75t_L g1284 ( .A1(n_453), .A2(n_1285), .A3(n_1288), .B1(n_1293), .B2(n_1294), .B3(n_1295), .Y(n_1284) );
OAI33xp33_ASAP7_75t_L g1535 ( .A1(n_453), .A2(n_488), .A3(n_1536), .B1(n_1540), .B2(n_1545), .B3(n_1549), .Y(n_1535) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_460), .B2(n_465), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g666 ( .A(n_458), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g1210 ( .A1(n_460), .A2(n_806), .B1(n_1211), .B2(n_1212), .Y(n_1210) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g487 ( .A(n_462), .Y(n_487) );
INVx2_ASAP7_75t_L g1015 ( .A(n_462), .Y(n_1015) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_463), .B(n_464), .Y(n_643) );
INVx1_ASAP7_75t_L g579 ( .A(n_464), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_470), .B1(n_471), .B2(n_474), .Y(n_466) );
BUFx2_ASAP7_75t_L g811 ( .A(n_467), .Y(n_811) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g1120 ( .A(n_468), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g1290 ( .A(n_468), .Y(n_1290) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g478 ( .A(n_469), .Y(n_478) );
BUFx2_ASAP7_75t_L g673 ( .A(n_469), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_471), .A2(n_476), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g875 ( .A(n_472), .Y(n_875) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_SL g545 ( .A(n_473), .Y(n_545) );
INVx2_ASAP7_75t_SL g569 ( .A(n_473), .Y(n_569) );
INVx4_ASAP7_75t_L g663 ( .A(n_473), .Y(n_663) );
INVx2_ASAP7_75t_SL g982 ( .A(n_473), .Y(n_982) );
INVx2_ASAP7_75t_SL g1164 ( .A(n_473), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_476), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
INVx2_ASAP7_75t_L g981 ( .A(n_476), .Y(n_981) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g544 ( .A(n_477), .Y(n_544) );
INVx2_ASAP7_75t_SL g999 ( .A(n_477), .Y(n_999) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g816 ( .A(n_478), .Y(n_816) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g559 ( .A(n_481), .Y(n_559) );
INVx2_ASAP7_75t_L g674 ( .A(n_481), .Y(n_674) );
INVx2_ASAP7_75t_L g776 ( .A(n_481), .Y(n_776) );
OAI22xp33_ASAP7_75t_L g1206 ( .A1(n_483), .A2(n_1207), .B1(n_1208), .B2(n_1209), .Y(n_1206) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_485), .A2(n_487), .B1(n_512), .B2(n_561), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_485), .A2(n_487), .B1(n_571), .B2(n_572), .Y(n_570) );
OAI22xp5_ASAP7_75t_SL g676 ( .A1(n_485), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g807 ( .A(n_485), .Y(n_807) );
OAI221xp5_ASAP7_75t_L g1597 ( .A1(n_485), .A2(n_642), .B1(n_1598), .B2(n_1599), .C(n_1600), .Y(n_1597) );
OAI221xp5_ASAP7_75t_L g1603 ( .A1(n_485), .A2(n_487), .B1(n_1588), .B2(n_1604), .C(n_1605), .Y(n_1603) );
OAI22xp33_ASAP7_75t_L g805 ( .A1(n_486), .A2(n_806), .B1(n_808), .B2(n_809), .Y(n_805) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI33xp33_ASAP7_75t_L g803 ( .A1(n_488), .A2(n_804), .A3(n_805), .B1(n_810), .B2(n_814), .B3(n_819), .Y(n_803) );
INVx1_ASAP7_75t_L g881 ( .A(n_488), .Y(n_881) );
CKINVDCx8_ASAP7_75t_R g488 ( .A(n_489), .Y(n_488) );
INVx5_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx6_ASAP7_75t_L g554 ( .A(n_490), .Y(n_554) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g987 ( .A(n_492), .Y(n_987) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
OAI22x1_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_647), .B2(n_724), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
XNOR2x1_ASAP7_75t_L g498 ( .A(n_499), .B(n_582), .Y(n_498) );
XNOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_541), .Y(n_501) );
AOI31xp33_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_516), .A3(n_526), .B(n_538), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g1566 ( .A1(n_505), .A2(n_1098), .B1(n_1530), .B2(n_1532), .C(n_1567), .Y(n_1566) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g587 ( .A(n_506), .Y(n_587) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_506), .Y(n_702) );
INVx2_ASAP7_75t_L g717 ( .A(n_506), .Y(n_717) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g1189 ( .A(n_509), .Y(n_1189) );
INVx2_ASAP7_75t_SL g696 ( .A(n_513), .Y(n_696) );
INVx2_ASAP7_75t_SL g735 ( .A(n_513), .Y(n_735) );
INVx1_ASAP7_75t_L g898 ( .A(n_513), .Y(n_898) );
AOI322xp5_ASAP7_75t_L g1234 ( .A1(n_513), .A2(n_737), .A3(n_1235), .B1(n_1238), .B2(n_1240), .C1(n_1242), .C2(n_1243), .Y(n_1234) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_514), .A2(n_515), .B1(n_575), .B2(n_577), .C(n_580), .Y(n_574) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g1239 ( .A(n_519), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_520), .Y(n_905) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g758 ( .A(n_521), .Y(n_758) );
INVxp67_ASAP7_75t_L g713 ( .A(n_523), .Y(n_713) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g534 ( .A(n_525), .Y(n_534) );
INVx1_ASAP7_75t_L g1273 ( .A(n_525), .Y(n_1273) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_532), .B1(n_535), .B2(n_537), .Y(n_526) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_531), .A2(n_661), .B1(n_667), .B2(n_706), .C(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g903 ( .A(n_531), .Y(n_903) );
BUFx2_ASAP7_75t_L g953 ( .A(n_533), .Y(n_953) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_537), .A2(n_563), .B1(n_565), .B2(n_573), .Y(n_562) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI211xp5_ASAP7_75t_L g583 ( .A1(n_539), .A2(n_584), .B(n_622), .C(n_633), .Y(n_583) );
NOR2xp67_ASAP7_75t_L g967 ( .A(n_539), .B(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g563 ( .A(n_540), .B(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g721 ( .A(n_540), .Y(n_721) );
OR2x6_ASAP7_75t_L g946 ( .A(n_540), .B(n_612), .Y(n_946) );
AND2x4_ASAP7_75t_L g1155 ( .A(n_540), .B(n_564), .Y(n_1155) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_562), .C(n_574), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g1540 ( .A1(n_544), .A2(n_1541), .B1(n_1542), .B2(n_1543), .Y(n_1540) );
OAI22xp5_ASAP7_75t_L g1594 ( .A1(n_545), .A2(n_999), .B1(n_1595), .B2(n_1596), .Y(n_1594) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_550), .B2(n_551), .Y(n_546) );
INVx1_ASAP7_75t_L g985 ( .A(n_548), .Y(n_985) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g1050 ( .A(n_549), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1157 ( .A(n_549), .Y(n_1157) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g770 ( .A(n_552), .Y(n_770) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AOI322xp5_ASAP7_75t_L g634 ( .A1(n_554), .A2(n_563), .A3(n_614), .B1(n_635), .B2(n_637), .C1(n_639), .C2(n_644), .Y(n_634) );
AOI33xp33_ASAP7_75t_L g768 ( .A1(n_554), .A2(n_563), .A3(n_769), .B1(n_771), .B2(n_774), .B3(n_777), .Y(n_768) );
INVx2_ASAP7_75t_L g1131 ( .A(n_554), .Y(n_1131) );
AOI33xp33_ASAP7_75t_L g1153 ( .A1(n_554), .A2(n_1154), .A3(n_1156), .B1(n_1160), .B2(n_1165), .B3(n_1166), .Y(n_1153) );
INVx1_ASAP7_75t_L g1295 ( .A(n_554), .Y(n_1295) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g1544 ( .A(n_559), .Y(n_1544) );
INVx1_ASAP7_75t_L g1013 ( .A(n_564), .Y(n_1013) );
BUFx2_ASAP7_75t_SL g1600 ( .A(n_564), .Y(n_1600) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_573), .A2(n_577), .B1(n_593), .B2(n_626), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_573), .A2(n_1036), .B1(n_1037), .B2(n_1038), .Y(n_1035) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_575), .A2(n_580), .B(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_575), .A2(n_577), .B1(n_580), .B2(n_766), .C(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g1083 ( .A(n_575), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g1142 ( .A1(n_575), .A2(n_1080), .B1(n_1143), .B2(n_1144), .C(n_1145), .Y(n_1142) );
AND2x2_ASAP7_75t_L g990 ( .A(n_576), .B(n_969), .Y(n_990) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_576), .B(n_969), .Y(n_1609) );
INVx1_ASAP7_75t_L g1081 ( .A(n_577), .Y(n_1081) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g1079 ( .A1(n_580), .A2(n_1073), .B1(n_1074), .B2(n_1080), .C(n_1082), .Y(n_1079) );
AOI221xp5_ASAP7_75t_L g1137 ( .A1(n_580), .A2(n_1080), .B1(n_1082), .B2(n_1110), .C(n_1111), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1145 ( .A(n_580), .Y(n_1145) );
NAND4xp25_ASAP7_75t_L g584 ( .A(n_585), .B(n_592), .C(n_601), .D(n_613), .Y(n_584) );
INVx1_ASAP7_75t_L g1565 ( .A(n_588), .Y(n_1565) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_590), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g759 ( .A(n_590), .Y(n_759) );
INVx1_ASAP7_75t_L g906 ( .A(n_590), .Y(n_906) );
OAI221xp5_ASAP7_75t_L g1095 ( .A1(n_591), .A2(n_1067), .B1(n_1096), .B2(n_1097), .C(n_1098), .Y(n_1095) );
A2O1A1Ixp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_596), .C(n_599), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_SL g1101 ( .A1(n_594), .A2(n_599), .B(n_754), .C(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx4_ASAP7_75t_L g685 ( .A(n_595), .Y(n_685) );
INVx2_ASAP7_75t_L g892 ( .A(n_595), .Y(n_892) );
A2O1A1Ixp33_ASAP7_75t_L g1071 ( .A1(n_599), .A2(n_620), .B(n_839), .C(n_1038), .Y(n_1071) );
BUFx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B(n_605), .C(n_607), .Y(n_601) );
BUFx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g616 ( .A(n_604), .Y(n_616) );
OR2x6_ASAP7_75t_L g923 ( .A(n_604), .B(n_920), .Y(n_923) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_606), .Y(n_950) );
INVx1_ASAP7_75t_L g1060 ( .A(n_606), .Y(n_1060) );
INVx2_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g932 ( .A(n_609), .Y(n_932) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_617), .C(n_619), .Y(n_613) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_SL g691 ( .A(n_618), .Y(n_691) );
BUFx3_ASAP7_75t_L g948 ( .A(n_618), .Y(n_948) );
INVx1_ASAP7_75t_L g719 ( .A(n_621), .Y(n_719) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g651 ( .A(n_624), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_631), .B2(n_632), .Y(n_627) );
INVx1_ASAP7_75t_L g681 ( .A(n_629), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_630), .B(n_969), .Y(n_968) );
INVx2_ASAP7_75t_L g654 ( .A(n_632), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_645), .Y(n_633) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_638), .Y(n_780) );
BUFx3_ASAP7_75t_L g668 ( .A(n_642), .Y(n_668) );
INVx2_ASAP7_75t_L g680 ( .A(n_642), .Y(n_680) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g724 ( .A(n_647), .Y(n_724) );
INVx1_ASAP7_75t_L g722 ( .A(n_648), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_655), .C(n_682), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_657), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_662), .A2(n_665), .B1(n_701), .B2(n_703), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_663), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_663), .A2(n_815), .B1(n_817), .B2(n_818), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_666), .A2(n_1090), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1127 ( .A1(n_666), .A2(n_1128), .B1(n_1129), .B2(n_1130), .Y(n_1127) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_668), .A2(n_865), .B1(n_867), .B2(n_868), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g877 ( .A1(n_668), .A2(n_865), .B1(n_878), .B2(n_879), .Y(n_877) );
BUFx3_ASAP7_75t_L g1007 ( .A(n_668), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_674), .B2(n_675), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_670), .A2(n_678), .B1(n_690), .B2(n_692), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g1042 ( .A1(n_671), .A2(n_1043), .B1(n_1044), .B2(n_1047), .C(n_1048), .Y(n_1042) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx2_ASAP7_75t_L g1546 ( .A(n_673), .Y(n_1546) );
OAI22xp5_ASAP7_75t_L g1203 ( .A1(n_674), .A2(n_811), .B1(n_1204), .B2(n_1205), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_675), .A2(n_677), .B1(n_685), .B2(n_686), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_679), .A2(n_806), .B1(n_820), .B2(n_821), .Y(n_819) );
OAI22xp33_ASAP7_75t_L g1285 ( .A1(n_679), .A2(n_1009), .B1(n_1286), .B2(n_1287), .Y(n_1285) );
OAI22xp33_ASAP7_75t_L g1294 ( .A1(n_679), .A2(n_982), .B1(n_1267), .B2(n_1276), .Y(n_1294) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g1129 ( .A(n_680), .Y(n_1129) );
INVx1_ASAP7_75t_L g1209 ( .A(n_680), .Y(n_1209) );
OAI31xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_695), .A3(n_699), .B(n_720), .Y(n_682) );
BUFx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OR2x6_ASAP7_75t_L g919 ( .A(n_688), .B(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_693), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_693), .B(n_963), .Y(n_962) );
OR2x6_ASAP7_75t_L g943 ( .A(n_698), .B(n_940), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_705), .B1(n_711), .B2(n_715), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g715 ( .A1(n_706), .A2(n_716), .B1(n_717), .B2(n_718), .C(n_719), .Y(n_715) );
BUFx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g753 ( .A(n_710), .Y(n_753) );
INVx2_ASAP7_75t_L g1621 ( .A(n_710), .Y(n_1621) );
OAI31xp33_ASAP7_75t_SL g1056 ( .A1(n_720), .A2(n_1057), .A3(n_1063), .B(n_1070), .Y(n_1056) );
CKINVDCx8_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
AOI31xp33_ASAP7_75t_L g1170 ( .A1(n_721), .A2(n_1171), .A3(n_1178), .B(n_1190), .Y(n_1170) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_847), .B1(n_1021), .B2(n_1022), .Y(n_726) );
INVx1_ASAP7_75t_L g1021 ( .A(n_727), .Y(n_1021) );
XOR2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_789), .Y(n_727) );
XNOR2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_788), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_764), .Y(n_729) );
NAND3xp33_ASAP7_75t_SL g731 ( .A(n_732), .B(n_747), .C(n_760), .Y(n_731) );
INVx2_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI21xp5_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_744), .B(n_745), .Y(n_741) );
INVx2_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g1089 ( .A(n_743), .Y(n_1089) );
INVx1_ASAP7_75t_L g1567 ( .A(n_743), .Y(n_1567) );
INVx1_ASAP7_75t_L g1177 ( .A(n_746), .Y(n_1177) );
BUFx2_ASAP7_75t_L g1241 ( .A(n_746), .Y(n_1241) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_753), .A2(n_1089), .B1(n_1090), .B2(n_1091), .C(n_1092), .Y(n_1088) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND4x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_768), .C(n_781), .D(n_784), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g872 ( .A(n_773), .Y(n_872) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx3_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
XNOR2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_822), .Y(n_791) );
NOR3xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_800), .C(n_803), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .Y(n_793) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_815), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_815), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_873) );
BUFx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_826), .B1(n_845), .B2(n_846), .Y(n_822) );
INVx1_ASAP7_75t_SL g911 ( .A(n_823), .Y(n_911) );
INVx5_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OAI31xp33_ASAP7_75t_L g1592 ( .A1(n_824), .A2(n_1593), .A3(n_1602), .B(n_1610), .Y(n_1592) );
BUFx8_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
OAI31xp33_ASAP7_75t_L g972 ( .A1(n_825), .A2(n_973), .A3(n_993), .B(n_1016), .Y(n_972) );
INVx2_ASAP7_75t_L g1227 ( .A(n_825), .Y(n_1227) );
AOI31xp33_ASAP7_75t_L g1255 ( .A1(n_825), .A2(n_1256), .A3(n_1266), .B(n_1274), .Y(n_1255) );
NAND3xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_831), .C(n_837), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_839), .Y(n_902) );
INVx1_ASAP7_75t_L g1077 ( .A(n_841), .Y(n_1077) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_844), .A2(n_1108), .B1(n_1110), .B2(n_1111), .Y(n_1107) );
AOI21xp5_ASAP7_75t_L g882 ( .A1(n_846), .A2(n_883), .B(n_884), .Y(n_882) );
INVx1_ASAP7_75t_L g1022 ( .A(n_847), .Y(n_1022) );
XOR2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_912), .Y(n_847) );
XNOR2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_882), .Y(n_850) );
NOR3xp33_ASAP7_75t_SL g851 ( .A(n_852), .B(n_861), .C(n_863), .Y(n_851) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
AOI21xp5_ASAP7_75t_L g1112 ( .A1(n_854), .A2(n_1097), .B(n_1113), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_854), .A2(n_856), .B1(n_1264), .B2(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx3_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AOI221xp5_ASAP7_75t_SL g885 ( .A1(n_874), .A2(n_886), .B1(n_893), .B2(n_895), .C(n_897), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g899 ( .A1(n_879), .A2(n_900), .B1(n_904), .B2(n_907), .C(n_909), .Y(n_899) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
AOI31xp33_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_899), .A3(n_910), .B(n_911), .Y(n_884) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx3_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g1185 ( .A(n_890), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
CKINVDCx5p33_ASAP7_75t_R g907 ( .A(n_908), .Y(n_907) );
AND3x1_ASAP7_75t_L g913 ( .A(n_914), .B(n_964), .C(n_972), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_915), .B(n_933), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_916), .B(n_924), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_918), .B1(n_921), .B2(n_922), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g979 ( .A1(n_917), .A2(n_930), .B1(n_980), .B2(n_982), .C(n_983), .Y(n_979) );
CKINVDCx6p67_ASAP7_75t_R g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g929 ( .A(n_920), .Y(n_929) );
CKINVDCx6p67_ASAP7_75t_R g922 ( .A(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_926), .B1(n_930), .B2(n_931), .Y(n_924) );
AOI221xp5_ASAP7_75t_L g1586 ( .A1(n_926), .A2(n_931), .B1(n_1587), .B2(n_1588), .C(n_1589), .Y(n_1586) );
AND2x2_ASAP7_75t_L g926 ( .A(n_927), .B(n_929), .Y(n_926) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_927), .Y(n_1187) );
INVx2_ASAP7_75t_SL g927 ( .A(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g1618 ( .A(n_928), .Y(n_1618) );
AND2x2_ASAP7_75t_L g931 ( .A(n_929), .B(n_932), .Y(n_931) );
NAND3xp33_ASAP7_75t_SL g933 ( .A(n_934), .B(n_944), .C(n_960), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_936), .B1(n_941), .B2(n_942), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_935), .A2(n_941), .B1(n_989), .B2(n_991), .Y(n_988) );
INVx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g1582 ( .A(n_937), .Y(n_1582) );
NAND2x1p5_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
INVx2_ASAP7_75t_SL g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g963 ( .A(n_940), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g1581 ( .A1(n_942), .A2(n_1582), .B1(n_1583), .B2(n_1584), .C(n_1585), .Y(n_1581) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
AOI33xp33_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_947), .A3(n_949), .B1(n_952), .B2(n_954), .B3(n_958), .Y(n_944) );
AOI33xp33_ASAP7_75t_L g1611 ( .A1(n_945), .A2(n_958), .A3(n_1612), .B1(n_1613), .B2(n_1617), .B3(n_1619), .Y(n_1611) );
CKINVDCx5p33_ASAP7_75t_R g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g1614 ( .A(n_956), .Y(n_1614) );
BUFx4f_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_966), .B(n_1591), .Y(n_1590) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_970), .B(n_1015), .Y(n_1014) );
OR2x6_ASAP7_75t_L g1601 ( .A(n_970), .B(n_1015), .Y(n_1601) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx8_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
AND2x4_ASAP7_75t_L g975 ( .A(n_976), .B(n_978), .Y(n_975) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_976), .B(n_1004), .Y(n_1020) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
BUFx6f_ASAP7_75t_L g1055 ( .A(n_978), .Y(n_1055) );
INVx2_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
OAI221xp5_ASAP7_75t_L g1051 ( .A1(n_982), .A2(n_999), .B1(n_1052), .B2(n_1053), .C(n_1054), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1288 ( .A1(n_982), .A2(n_1289), .B1(n_1291), .B2(n_1292), .Y(n_1288) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1605 ( .A(n_986), .Y(n_1605) );
INVx2_ASAP7_75t_SL g986 ( .A(n_987), .Y(n_986) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
AOI22xp5_ASAP7_75t_L g1608 ( .A1(n_991), .A2(n_1583), .B1(n_1584), .B2(n_1609), .Y(n_1608) );
CKINVDCx11_ASAP7_75t_R g991 ( .A(n_992), .Y(n_991) );
CKINVDCx6p67_ASAP7_75t_R g994 ( .A(n_995), .Y(n_994) );
OAI22xp5_ASAP7_75t_SL g996 ( .A1(n_997), .A2(n_998), .B1(n_1000), .B2(n_1001), .Y(n_996) );
OAI22xp33_ASAP7_75t_L g1293 ( .A1(n_998), .A2(n_1009), .B1(n_1257), .B2(n_1275), .Y(n_1293) );
BUFx2_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_999), .A2(n_1123), .B1(n_1124), .B2(n_1126), .Y(n_1122) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
OAI221xp5_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1009), .B2(n_1011), .C(n_1012), .Y(n_1006) );
OAI22xp33_ASAP7_75t_L g1536 ( .A1(n_1007), .A2(n_1537), .B1(n_1538), .B2(n_1539), .Y(n_1536) );
BUFx2_ASAP7_75t_L g1538 ( .A(n_1009), .Y(n_1538) );
INVx2_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1015), .Y(n_1117) );
INVx3_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx3_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
XNOR2xp5_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1195), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1138), .B1(n_1193), .B2(n_1194), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1193 ( .A(n_1027), .Y(n_1193) );
XOR2x2_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1084), .Y(n_1027) );
NAND4xp25_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1039), .C(n_1056), .D(n_1079), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1035), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1545 ( .A1(n_1044), .A2(n_1546), .B1(n_1547), .B2(n_1548), .Y(n_1545) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_1046), .A2(n_1091), .B1(n_1119), .B2(n_1121), .Y(n_1118) );
INVx3_ASAP7_75t_L g1125 ( .A(n_1046), .Y(n_1125) );
INVx2_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
HB1xp67_ASAP7_75t_L g1561 ( .A(n_1058), .Y(n_1561) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
OAI221xp5_ASAP7_75t_L g1175 ( .A1(n_1067), .A2(n_1149), .B1(n_1151), .B2(n_1176), .C(n_1177), .Y(n_1175) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
NAND3xp33_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1072), .C(n_1075), .Y(n_1070) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
NAND4xp25_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1112), .C(n_1132), .D(n_1137), .Y(n_1085) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
NAND3xp33_ASAP7_75t_SL g1100 ( .A(n_1101), .B(n_1103), .C(n_1107), .Y(n_1100) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1606 ( .A1(n_1119), .A2(n_1124), .B1(n_1587), .B2(n_1607), .Y(n_1606) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
OAI22xp33_ASAP7_75t_L g1549 ( .A1(n_1129), .A2(n_1538), .B1(n_1550), .B2(n_1551), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1135), .Y(n_1132) );
INVxp67_ASAP7_75t_L g1194 ( .A(n_1138), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1167), .Y(n_1140) );
AND4x1_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1146), .C(n_1150), .D(n_1153), .Y(n_1141) );
BUFx3_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
BUFx3_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
AOI21xp33_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1169), .B(n_1170), .Y(n_1167) );
AOI21xp5_ASAP7_75t_L g1552 ( .A1(n_1168), .A2(n_1553), .B(n_1554), .Y(n_1552) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_1177), .A2(n_1261), .B1(n_1262), .B2(n_1263), .C(n_1264), .Y(n_1260) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_1196), .A2(n_1248), .B1(n_1249), .B2(n_1297), .Y(n_1195) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1196), .Y(n_1297) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1226), .Y(n_1200) );
NOR3xp33_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1216), .C(n_1218), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1223), .Y(n_1218) );
NAND4xp25_ASAP7_75t_L g1228 ( .A(n_1229), .B(n_1234), .C(n_1244), .D(n_1245), .Y(n_1228) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx2_ASAP7_75t_SL g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1277), .Y(n_1251) );
AOI21xp5_ASAP7_75t_L g1252 ( .A1(n_1253), .A2(n_1254), .B(n_1255), .Y(n_1252) );
AOI211xp5_ASAP7_75t_L g1256 ( .A1(n_1257), .A2(n_1258), .B(n_1259), .C(n_1265), .Y(n_1256) );
BUFx2_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NOR3xp33_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1283), .C(n_1284), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1281), .Y(n_1278) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
OAI221xp5_ASAP7_75t_L g1299 ( .A1(n_1300), .A2(n_1523), .B1(n_1524), .B2(n_1571), .C(n_1574), .Y(n_1299) );
NOR2xp67_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1461), .Y(n_1300) );
OAI21xp33_ASAP7_75t_L g1301 ( .A1(n_1302), .A2(n_1416), .B(n_1425), .Y(n_1301) );
NOR5xp2_ASAP7_75t_SL g1302 ( .A(n_1303), .B(n_1356), .C(n_1384), .D(n_1396), .E(n_1404), .Y(n_1302) );
NOR2xp33_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1331), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1438 ( .A1(n_1304), .A2(n_1409), .B1(n_1439), .B2(n_1441), .Y(n_1438) );
OAI211xp5_ASAP7_75t_L g1468 ( .A1(n_1304), .A2(n_1399), .B(n_1469), .C(n_1471), .Y(n_1468) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1304), .B(n_1472), .Y(n_1488) );
HB1xp67_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx2_ASAP7_75t_SL g1379 ( .A(n_1305), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1305), .B(n_1345), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1305), .B(n_1360), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1305), .B(n_1459), .Y(n_1458) );
AND2x4_ASAP7_75t_L g1467 ( .A(n_1305), .B(n_1359), .Y(n_1467) );
NOR2xp33_ASAP7_75t_L g1476 ( .A(n_1305), .B(n_1459), .Y(n_1476) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1305), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_1305), .B(n_1450), .Y(n_1513) );
CKINVDCx5p33_ASAP7_75t_R g1305 ( .A(n_1306), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1306), .B(n_1359), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1306), .B(n_1360), .Y(n_1411) );
OR2x2_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1321), .Y(n_1306) );
OAI22xp5_ASAP7_75t_L g1307 ( .A1(n_1308), .A2(n_1315), .B1(n_1316), .B2(n_1320), .Y(n_1307) );
BUFx3_ASAP7_75t_L g1422 ( .A(n_1308), .Y(n_1422) );
BUFx6f_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1353 ( .A1(n_1309), .A2(n_1318), .B1(n_1354), .B2(n_1355), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1311), .Y(n_1309) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1310), .B(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1310), .Y(n_1338) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1311), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1314), .Y(n_1311) );
HB1xp67_ASAP7_75t_L g1624 ( .A(n_1312), .Y(n_1624) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1314), .Y(n_1325) );
HB1xp67_ASAP7_75t_L g1424 ( .A(n_1316), .Y(n_1424) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1319), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g1321 ( .A1(n_1322), .A2(n_1327), .B1(n_1328), .B2(n_1330), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
BUFx3_ASAP7_75t_L g1419 ( .A(n_1323), .Y(n_1419) );
AND2x4_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1326), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1324), .B(n_1326), .Y(n_1342) );
HB1xp67_ASAP7_75t_L g1625 ( .A(n_1324), .Y(n_1625) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
AND2x4_ASAP7_75t_L g1329 ( .A(n_1325), .B(n_1326), .Y(n_1329) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1328), .Y(n_1376) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1343), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1333), .B(n_1370), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1333), .B(n_1382), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1333), .B(n_1367), .Y(n_1496) );
INVxp67_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
BUFx3_ASAP7_75t_L g1366 ( .A(n_1334), .Y(n_1366) );
BUFx2_ASAP7_75t_L g1381 ( .A(n_1334), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1334), .B(n_1370), .Y(n_1409) );
AOI222xp33_ASAP7_75t_L g1443 ( .A1(n_1334), .A2(n_1380), .B1(n_1395), .B2(n_1411), .C1(n_1444), .C2(n_1445), .Y(n_1443) );
NOR3xp33_ASAP7_75t_L g1498 ( .A(n_1334), .B(n_1398), .C(n_1479), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1341), .Y(n_1334) );
AND2x4_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1338), .Y(n_1336) );
AND2x4_ASAP7_75t_L g1339 ( .A(n_1338), .B(n_1340), .Y(n_1339) );
BUFx2_ASAP7_75t_L g1374 ( .A(n_1339), .Y(n_1374) );
NOR2xp33_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1348), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1344), .B(n_1401), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1344), .B(n_1379), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_1344), .B(n_1467), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1516 ( .A(n_1344), .B(n_1517), .Y(n_1516) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
BUFx2_ASAP7_75t_L g1363 ( .A(n_1345), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1407 ( .A(n_1345), .B(n_1366), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1345), .B(n_1381), .Y(n_1431) );
INVx2_ASAP7_75t_L g1459 ( .A(n_1345), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1345), .B(n_1394), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1347), .Y(n_1345) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1348), .Y(n_1370) );
OR2x2_ASAP7_75t_L g1506 ( .A(n_1348), .B(n_1407), .Y(n_1506) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1352), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1349), .B(n_1368), .Y(n_1367) );
INVx2_ASAP7_75t_L g1383 ( .A(n_1349), .Y(n_1383) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_1349), .B(n_1366), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1349), .B(n_1352), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1349), .B(n_1366), .Y(n_1413) );
OAI321xp33_ASAP7_75t_L g1474 ( .A1(n_1349), .A2(n_1475), .A3(n_1477), .B1(n_1479), .B2(n_1481), .C(n_1482), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1351), .Y(n_1349) );
INVx2_ASAP7_75t_SL g1368 ( .A(n_1352), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1352), .B(n_1383), .Y(n_1382) );
OAI222xp33_ASAP7_75t_L g1426 ( .A1(n_1352), .A2(n_1359), .B1(n_1427), .B2(n_1429), .C1(n_1432), .C2(n_1433), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1352), .B(n_1366), .Y(n_1517) );
OAI22xp5_ASAP7_75t_L g1356 ( .A1(n_1357), .A2(n_1364), .B1(n_1371), .B2(n_1377), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1363), .Y(n_1357) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1358), .Y(n_1473) );
OAI311xp33_ASAP7_75t_L g1494 ( .A1(n_1358), .A2(n_1416), .A3(n_1495), .B1(n_1497), .C1(n_1500), .Y(n_1494) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
NOR2xp33_ASAP7_75t_L g1414 ( .A(n_1359), .B(n_1415), .Y(n_1414) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_1359), .B(n_1478), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1359), .B(n_1372), .Y(n_1480) );
INVx3_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1360), .B(n_1372), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1360), .B(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1360), .Y(n_1520) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1362), .Y(n_1360) );
NAND2xp5_ASAP7_75t_SL g1387 ( .A(n_1363), .B(n_1388), .Y(n_1387) );
INVx2_ASAP7_75t_L g1398 ( .A(n_1363), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1363), .B(n_1428), .Y(n_1444) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1363), .B(n_1446), .Y(n_1445) );
AOI221xp5_ASAP7_75t_L g1462 ( .A1(n_1363), .A2(n_1463), .B1(n_1468), .B2(n_1473), .C(n_1474), .Y(n_1462) );
NOR2xp33_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1369), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1365), .B(n_1459), .Y(n_1472) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1365), .Y(n_1481) );
OAI21xp5_ASAP7_75t_SL g1500 ( .A1(n_1365), .A2(n_1501), .B(n_1502), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1367), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1366), .B(n_1368), .Y(n_1386) );
OR2x2_ASAP7_75t_L g1399 ( .A(n_1366), .B(n_1400), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1366), .B(n_1442), .Y(n_1441) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_1366), .B(n_1383), .Y(n_1486) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1367), .Y(n_1406) );
NAND3xp33_ASAP7_75t_SL g1482 ( .A(n_1367), .B(n_1436), .C(n_1483), .Y(n_1482) );
AOI321xp33_ASAP7_75t_L g1489 ( .A1(n_1368), .A2(n_1379), .A3(n_1401), .B1(n_1490), .B2(n_1491), .C(n_1492), .Y(n_1489) );
NOR2x1_ASAP7_75t_L g1501 ( .A(n_1368), .B(n_1381), .Y(n_1501) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1369), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1370), .B(n_1393), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1370), .B(n_1431), .Y(n_1470) );
NOR2xp33_ASAP7_75t_L g1491 ( .A(n_1371), .B(n_1379), .Y(n_1491) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1371), .Y(n_1514) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1372), .Y(n_1391) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1372), .Y(n_1394) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1372), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1375), .Y(n_1372) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1378), .B(n_1380), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1378), .B(n_1440), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1378), .B(n_1470), .Y(n_1469) );
INVx2_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1379), .B(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1379), .Y(n_1403) );
NOR2xp33_ASAP7_75t_L g1505 ( .A(n_1379), .B(n_1506), .Y(n_1505) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1380), .B(n_1398), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1382), .Y(n_1380) );
NOR2xp33_ASAP7_75t_L g1446 ( .A(n_1381), .B(n_1383), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1382), .B(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1382), .Y(n_1464) );
A2O1A1Ixp33_ASAP7_75t_L g1384 ( .A1(n_1385), .A2(n_1387), .B(n_1389), .C(n_1392), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1388), .B(n_1398), .Y(n_1433) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
AOI211xp5_ASAP7_75t_L g1504 ( .A1(n_1390), .A2(n_1505), .B(n_1507), .C(n_1519), .Y(n_1504) );
NAND2xp5_ASAP7_75t_L g1518 ( .A(n_1390), .B(n_1512), .Y(n_1518) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1391), .Y(n_1436) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1391), .Y(n_1450) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1393), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1395), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1394), .B(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1394), .Y(n_1456) );
AOI32xp33_ASAP7_75t_L g1497 ( .A1(n_1395), .A2(n_1413), .A3(n_1490), .B1(n_1498), .B2(n_1499), .Y(n_1497) );
AOI21xp33_ASAP7_75t_L g1396 ( .A1(n_1397), .A2(n_1399), .B(n_1402), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1398), .B(n_1428), .Y(n_1432) );
OR2x2_ASAP7_75t_L g1495 ( .A(n_1398), .B(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1401), .B(n_1431), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1401), .B(n_1509), .Y(n_1508) );
A2O1A1Ixp33_ASAP7_75t_L g1404 ( .A1(n_1405), .A2(n_1408), .B(n_1410), .C(n_1412), .Y(n_1404) );
OR2x2_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1407), .Y(n_1405) );
NOR3xp33_ASAP7_75t_L g1492 ( .A(n_1406), .B(n_1456), .C(n_1493), .Y(n_1492) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1406), .B(n_1464), .Y(n_1499) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1407), .Y(n_1509) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
OR2x2_ASAP7_75t_L g1452 ( .A(n_1410), .B(n_1453), .Y(n_1452) );
CKINVDCx5p33_ASAP7_75t_R g1410 ( .A(n_1411), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1413), .B(n_1414), .Y(n_1412) );
INVx2_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx3_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1418), .B(n_1435), .Y(n_1434) );
INVx3_ASAP7_75t_L g1449 ( .A(n_1418), .Y(n_1449) );
AOI21xp5_ASAP7_75t_L g1484 ( .A1(n_1418), .A2(n_1485), .B(n_1494), .Y(n_1484) );
O2A1O1Ixp33_ASAP7_75t_L g1510 ( .A1(n_1418), .A2(n_1511), .B(n_1513), .C(n_1514), .Y(n_1510) );
CKINVDCx5p33_ASAP7_75t_R g1523 ( .A(n_1419), .Y(n_1523) );
OAI22xp33_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1422), .B1(n_1423), .B2(n_1424), .Y(n_1420) );
AOI221xp5_ASAP7_75t_L g1425 ( .A1(n_1426), .A2(n_1434), .B1(n_1437), .B2(n_1447), .C(n_1451), .Y(n_1425) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1521 ( .A(n_1428), .B(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
OAI222xp33_ASAP7_75t_L g1507 ( .A1(n_1433), .A2(n_1465), .B1(n_1508), .B2(n_1510), .C1(n_1515), .C2(n_1518), .Y(n_1507) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1436), .Y(n_1453) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1443), .Y(n_1437) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1450), .Y(n_1448) );
OAI211xp5_ASAP7_75t_L g1461 ( .A1(n_1449), .A2(n_1462), .B(n_1484), .C(n_1504), .Y(n_1461) );
O2A1O1Ixp33_ASAP7_75t_L g1519 ( .A1(n_1449), .A2(n_1506), .B(n_1520), .C(n_1521), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1450), .B(n_1467), .Y(n_1466) );
OAI21xp33_ASAP7_75t_L g1451 ( .A1(n_1452), .A2(n_1454), .B(n_1455), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1457), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1460), .Y(n_1457) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1458), .Y(n_1493) );
NOR2xp33_ASAP7_75t_L g1463 ( .A(n_1464), .B(n_1465), .Y(n_1463) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
OAI211xp5_ASAP7_75t_L g1485 ( .A1(n_1486), .A2(n_1487), .B(n_1488), .C(n_1489), .Y(n_1485) );
INVx2_ASAP7_75t_L g1522 ( .A(n_1496), .Y(n_1522) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1525), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1552), .Y(n_1525) );
NOR3xp33_ASAP7_75t_SL g1526 ( .A(n_1527), .B(n_1534), .C(n_1535), .Y(n_1526) );
NAND2xp5_ASAP7_75t_L g1527 ( .A(n_1528), .B(n_1531), .Y(n_1527) );
INVx2_ASAP7_75t_SL g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
CKINVDCx5p33_ASAP7_75t_R g1571 ( .A(n_1572), .Y(n_1571) );
A2O1A1Ixp33_ASAP7_75t_L g1622 ( .A1(n_1573), .A2(n_1623), .B(n_1625), .C(n_1626), .Y(n_1622) );
BUFx2_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
NAND4xp75_ASAP7_75t_SL g1579 ( .A(n_1580), .B(n_1590), .C(n_1592), .D(n_1611), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1586), .Y(n_1580) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVx2_ASAP7_75t_SL g1620 ( .A(n_1621), .Y(n_1620) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
endmodule