module fake_jpeg_1502_n_223 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_223);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx6f_ASAP7_75t_SL g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_13),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_84),
.Y(n_90)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_24),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_52),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_69),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_65),
.B1(n_75),
.B2(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_98),
.B1(n_59),
.B2(n_66),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_75),
.B1(n_65),
.B2(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_64),
.B1(n_83),
.B2(n_81),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_103),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_57),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_111),
.Y(n_124)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_119),
.B1(n_60),
.B2(n_70),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_54),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_61),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_66),
.B1(n_57),
.B2(n_76),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_88),
.B(n_73),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_71),
.B(n_74),
.Y(n_150)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_73),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_102),
.C(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_119),
.A2(n_78),
.B1(n_60),
.B2(n_67),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_135),
.B1(n_139),
.B2(n_141),
.Y(n_154)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_32),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_138),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_70),
.B1(n_56),
.B2(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_62),
.B1(n_58),
.B2(n_71),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_137),
.A2(n_118),
.B1(n_102),
.B2(n_105),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_43),
.B1(n_40),
.B2(n_39),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_152),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_162),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_74),
.B(n_71),
.C(n_51),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_151),
.A2(n_38),
.B(n_37),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_1),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_141),
.A2(n_71),
.B1(n_3),
.B2(n_4),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_157),
.B1(n_165),
.B2(n_139),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_48),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_162),
.C(n_149),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_R g158 ( 
.A(n_131),
.B(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_7),
.Y(n_169)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_120),
.B(n_47),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_164),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_171),
.C(n_185),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_129),
.B(n_133),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_151),
.B(n_154),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_174),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_25),
.C(n_45),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_175),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_152),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_46),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_177),
.B1(n_184),
.B2(n_175),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_184),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_35),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_178),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_196),
.B1(n_28),
.B2(n_26),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_147),
.B1(n_164),
.B2(n_153),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_181),
.B1(n_182),
.B2(n_173),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_148),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_195),
.B(n_181),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_166),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_203),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_171),
.C(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_202),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_188),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_193),
.B1(n_194),
.B2(n_187),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_34),
.C(n_33),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_10),
.C(n_12),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_10),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_186),
.B1(n_18),
.B2(n_19),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_209),
.A2(n_211),
.B1(n_14),
.B2(n_17),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_197),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_216),
.B(n_208),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_217),
.A2(n_215),
.B1(n_211),
.B2(n_216),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_218),
.A2(n_213),
.B(n_186),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_207),
.B(n_18),
.C(n_20),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_17),
.B(n_20),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_221),
.A2(n_21),
.B(n_22),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_22),
.Y(n_223)
);


endmodule