module fake_ariane_723_n_1907 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1907);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1907;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_39),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_177),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_72),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_74),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_149),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_32),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_11),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_88),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_87),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_20),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_26),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_94),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_53),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_115),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_1),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_95),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_98),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_43),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_80),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_13),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_45),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_67),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_61),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_61),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_23),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_162),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_176),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_86),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_56),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_110),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_59),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_129),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_68),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_137),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_12),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_0),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_153),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_76),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_42),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_126),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_151),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_91),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_141),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_100),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_107),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_144),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_40),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_23),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_125),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_179),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_9),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_50),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_128),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_24),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_32),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_24),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_27),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_27),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_145),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_3),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_155),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_14),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_33),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_22),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_34),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_92),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_182),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_28),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_136),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_170),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_64),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_49),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_169),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_143),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_39),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_12),
.Y(n_280)
);

BUFx8_ASAP7_75t_SL g281 ( 
.A(n_161),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_37),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_83),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_60),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_116),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_146),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_66),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_166),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_45),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_29),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_159),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_54),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_84),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_142),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_19),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_65),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_69),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_181),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_59),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_119),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_2),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_123),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_3),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_70),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_42),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_147),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_130),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_78),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_21),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_171),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_148),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_124),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_122),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_103),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_117),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_47),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_10),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_75),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_101),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_60),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_81),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_54),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_49),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_97),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_105),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_90),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_33),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_96),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_99),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_184),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_138),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_150),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_158),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_14),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_57),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_22),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_106),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_113),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_19),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_43),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_82),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_40),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_183),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_50),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_132),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_25),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_112),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_13),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_104),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_185),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_37),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_25),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_17),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_51),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_10),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_18),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_102),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_63),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_111),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_89),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_118),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_133),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_2),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_16),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_16),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_114),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_38),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_34),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_18),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_71),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_127),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_156),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_135),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_31),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_139),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_31),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_6),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_271),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_294),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_231),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_231),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_201),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_352),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_193),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_206),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_197),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_248),
.B(n_280),
.Y(n_390)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_186),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_209),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_300),
.B(n_0),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_210),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_213),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_235),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_261),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_252),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_189),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_205),
.B(n_1),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_189),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_186),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_266),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_279),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_205),
.B(n_4),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_282),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_216),
.B(n_5),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_283),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_216),
.B(n_6),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_189),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_290),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_315),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_304),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_196),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_306),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_335),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_324),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_304),
.B(n_7),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_357),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_196),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_346),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_370),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_348),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_380),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_262),
.Y(n_429)
);

NOR2xp67_ASAP7_75t_L g430 ( 
.A(n_219),
.B(n_310),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_268),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_376),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_196),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_310),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_355),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_221),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_187),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_237),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_187),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_272),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_188),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_262),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_188),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_199),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_262),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_262),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_190),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_190),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_286),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_268),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_366),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_192),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_262),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_191),
.B(n_7),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_351),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_351),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_192),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_195),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_351),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_195),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_202),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_281),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_233),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_351),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_202),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_199),
.B(n_8),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_351),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_194),
.B(n_8),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_233),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_328),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_200),
.B(n_11),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_379),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_218),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_268),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_269),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_239),
.Y(n_477)
);

INVxp33_ASAP7_75t_SL g478 ( 
.A(n_200),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_239),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_218),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_251),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_269),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_251),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_208),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_471),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_438),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_471),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_471),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_447),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_463),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_387),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_198),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_392),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_471),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_454),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_456),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_383),
.B(n_203),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_457),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_398),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_460),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_465),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_468),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_483),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_429),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_483),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_434),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_409),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_435),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_413),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_426),
.B(n_269),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_442),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_385),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_388),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_394),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_395),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_396),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_440),
.Y(n_521)
);

CKINVDCx11_ASAP7_75t_R g522 ( 
.A(n_450),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_400),
.B(n_223),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_397),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_452),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_389),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_400),
.B(n_223),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_404),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_405),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_417),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_407),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_473),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_425),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_418),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_384),
.B(n_208),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_420),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_381),
.Y(n_540)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_455),
.A2(n_211),
.B(n_207),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_421),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_427),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_432),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_437),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_422),
.Y(n_546)
);

OA21x2_ASAP7_75t_L g547 ( 
.A1(n_469),
.A2(n_215),
.B(n_214),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_437),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_389),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_428),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_403),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_475),
.B(n_288),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_401),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_439),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_439),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_441),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_441),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_464),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_402),
.B(n_226),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_419),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_444),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_470),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_444),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_513),
.B(n_431),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_517),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_513),
.B(n_414),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_517),
.B(n_445),
.Y(n_569)
);

INVx6_ASAP7_75t_L g570 ( 
.A(n_506),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_506),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_540),
.B(n_393),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_501),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_402),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_506),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_501),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_501),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_501),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_523),
.B(n_560),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_484),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_554),
.B(n_411),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_411),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_534),
.B(n_451),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_498),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_561),
.B(n_415),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_498),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_534),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_498),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_484),
.Y(n_589)
);

AND2x2_ASAP7_75t_SL g590 ( 
.A(n_541),
.B(n_393),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_541),
.A2(n_478),
.B1(n_391),
.B2(n_410),
.Y(n_591)
);

INVx4_ASAP7_75t_SL g592 ( 
.A(n_506),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_507),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_540),
.B(n_408),
.Y(n_594)
);

NOR2x1p5_ASAP7_75t_L g595 ( 
.A(n_545),
.B(n_549),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_527),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_555),
.B(n_448),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_553),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_562),
.B(n_415),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_539),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_498),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_498),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_539),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_493),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_507),
.B(n_424),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_490),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_546),
.Y(n_607)
);

AO22x2_ASAP7_75t_L g608 ( 
.A1(n_538),
.A2(n_482),
.B1(n_476),
.B2(n_259),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_546),
.B(n_433),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_541),
.A2(n_391),
.B1(n_478),
.B2(n_481),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_546),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_538),
.B(n_467),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_550),
.B(n_381),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_490),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_546),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_556),
.B(n_448),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_495),
.B(n_433),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_553),
.B(n_449),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_492),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_553),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_499),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_524),
.B(n_382),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_539),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_539),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_558),
.B(n_449),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_503),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_503),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_525),
.B(n_537),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_504),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_504),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_505),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_553),
.B(n_508),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_528),
.B(n_382),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_539),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_505),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_508),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_539),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_525),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_487),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_487),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_500),
.B(n_453),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_486),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_541),
.A2(n_477),
.B1(n_430),
.B2(n_472),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_525),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_537),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_487),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_552),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_537),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_522),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_486),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_487),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_518),
.B(n_453),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_563),
.B(n_386),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_487),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_486),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_565),
.B(n_458),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_518),
.B(n_458),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_515),
.B(n_459),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_491),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_509),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_509),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_494),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_511),
.Y(n_666)
);

INVxp33_ASAP7_75t_L g667 ( 
.A(n_485),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_487),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_515),
.B(n_480),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_516),
.B(n_459),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_516),
.B(n_461),
.Y(n_671)
);

NOR2x1p5_ASAP7_75t_L g672 ( 
.A(n_519),
.B(n_386),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_547),
.A2(n_519),
.B1(n_529),
.B2(n_520),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_520),
.B(n_204),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_511),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_529),
.B(n_461),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_530),
.B(n_462),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_530),
.B(n_462),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_532),
.B(n_204),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_532),
.B(n_466),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_533),
.B(n_466),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_533),
.B(n_474),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_491),
.Y(n_683)
);

BUFx8_ASAP7_75t_SL g684 ( 
.A(n_488),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_535),
.B(n_474),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_535),
.B(n_480),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_547),
.B(n_212),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_547),
.A2(n_254),
.B1(n_327),
.B2(n_363),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_542),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_548),
.B(n_373),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_547),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_496),
.Y(n_692)
);

OAI22x1_ASAP7_75t_L g693 ( 
.A1(n_485),
.A2(n_379),
.B1(n_284),
.B2(n_377),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_551),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_551),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_491),
.B(n_229),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_497),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_497),
.B(n_288),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_502),
.B(n_510),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_489),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_489),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_489),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_489),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_559),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_564),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_512),
.B(n_230),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_531),
.A2(n_222),
.B1(n_303),
.B2(n_224),
.Y(n_707)
);

AND3x4_ASAP7_75t_L g708 ( 
.A(n_521),
.B(n_314),
.C(n_220),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_580),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_576),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_576),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_579),
.A2(n_331),
.B1(n_222),
.B2(n_224),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_609),
.B(n_225),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_590),
.B(n_321),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_590),
.B(n_321),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_680),
.B(n_220),
.C(n_217),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_574),
.B(n_217),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_568),
.B(n_536),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_669),
.A2(n_303),
.B1(n_339),
.B2(n_330),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_581),
.B(n_323),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_582),
.B(n_544),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_577),
.Y(n_722)
);

AND2x2_ASAP7_75t_SL g723 ( 
.A(n_688),
.B(n_610),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_577),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_687),
.A2(n_314),
.B1(n_212),
.B2(n_244),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_580),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_589),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_640),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_640),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_585),
.B(n_323),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_599),
.B(n_326),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_589),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_593),
.B(n_330),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_567),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_687),
.A2(n_311),
.B1(n_278),
.B2(n_244),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_591),
.A2(n_227),
.B(n_228),
.C(n_377),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_598),
.B(n_334),
.Y(n_737)
);

NOR2x1p5_ASAP7_75t_L g738 ( 
.A(n_656),
.B(n_543),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_598),
.B(n_334),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_621),
.B(n_339),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_619),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_593),
.B(n_689),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_643),
.B(n_350),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_669),
.A2(n_353),
.B1(n_361),
.B2(n_375),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_646),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_619),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_617),
.B(n_526),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_621),
.B(n_353),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_655),
.B(n_361),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_625),
.B(n_364),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_604),
.B(n_227),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_655),
.B(n_364),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_660),
.B(n_369),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_694),
.A2(n_228),
.B(n_372),
.C(n_371),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_625),
.B(n_374),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_607),
.Y(n_756)
);

AO221x1_ASAP7_75t_L g757 ( 
.A1(n_693),
.A2(n_328),
.B1(n_313),
.B2(n_285),
.C(n_257),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_661),
.A2(n_374),
.B1(n_375),
.B2(n_378),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_661),
.B(n_236),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_678),
.A2(n_295),
.B1(n_292),
.B2(n_287),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_622),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_646),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_618),
.A2(n_677),
.B1(n_685),
.B2(n_670),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_SL g764 ( 
.A1(n_708),
.A2(n_372),
.B1(n_371),
.B2(n_367),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_622),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_647),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_647),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_625),
.B(n_232),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_650),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_678),
.B(n_240),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_682),
.B(n_249),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_682),
.B(n_250),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_608),
.A2(n_645),
.B1(n_679),
.B2(n_674),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_694),
.B(n_253),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_625),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_583),
.B(n_284),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_625),
.B(n_246),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_SL g778 ( 
.A(n_604),
.B(n_656),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_607),
.B(n_255),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_674),
.B(n_679),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_639),
.B(n_673),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_SL g782 ( 
.A1(n_708),
.A2(n_367),
.B1(n_359),
.B2(n_358),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_639),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_695),
.B(n_258),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_583),
.B(n_322),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_695),
.B(n_634),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_690),
.B(n_568),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_650),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_639),
.B(n_256),
.Y(n_789)
);

AND2x6_ASAP7_75t_SL g790 ( 
.A(n_572),
.B(n_322),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_630),
.B(n_260),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_628),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_639),
.B(n_263),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_573),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_630),
.B(n_264),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_608),
.A2(n_365),
.B1(n_362),
.B2(n_360),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_573),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_597),
.B(n_329),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_578),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_624),
.A2(n_299),
.B1(n_345),
.B2(n_343),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_608),
.A2(n_365),
.B1(n_362),
.B2(n_360),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_578),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_606),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_663),
.B(n_267),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_587),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_629),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_639),
.B(n_316),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_629),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_663),
.B(n_276),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_635),
.A2(n_332),
.B1(n_340),
.B2(n_301),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_614),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_664),
.B(n_291),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_664),
.B(n_293),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_649),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_633),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_649),
.B(n_329),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_666),
.B(n_296),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_666),
.B(n_675),
.Y(n_818)
);

INVx4_ASAP7_75t_L g819 ( 
.A(n_674),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_675),
.B(n_686),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_614),
.Y(n_821)
);

NAND3xp33_ASAP7_75t_L g822 ( 
.A(n_706),
.B(n_707),
.C(n_605),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_596),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_611),
.B(n_302),
.Y(n_824)
);

NOR2x1p5_ASAP7_75t_L g825 ( 
.A(n_652),
.B(n_336),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_691),
.A2(n_278),
.B(n_333),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_616),
.B(n_336),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_615),
.B(n_317),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_651),
.B(n_318),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_627),
.B(n_338),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_659),
.B(n_338),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_566),
.B(n_341),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_633),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_569),
.B(n_596),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_620),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_600),
.A2(n_311),
.B(n_333),
.C(n_234),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_600),
.B(n_328),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_575),
.A2(n_305),
.B(n_241),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_572),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_620),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_674),
.B(n_341),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_572),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_638),
.B(n_342),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_603),
.B(n_328),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_603),
.B(n_328),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_631),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_572),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_608),
.A2(n_356),
.B1(n_349),
.B2(n_347),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_631),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_674),
.B(n_344),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_674),
.A2(n_349),
.B1(n_347),
.B2(n_344),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_671),
.A2(n_15),
.B(n_20),
.C(n_21),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_684),
.Y(n_853)
);

OAI22xp33_ASAP7_75t_L g854 ( 
.A1(n_594),
.A2(n_320),
.B1(n_319),
.B2(n_312),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_674),
.A2(n_309),
.B1(n_308),
.B2(n_307),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_566),
.B(n_15),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_626),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_637),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_632),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_698),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_626),
.B(n_636),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_612),
.B(n_298),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_857),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_763),
.B(n_676),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_861),
.A2(n_681),
.B(n_571),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_776),
.B(n_623),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_822),
.A2(n_613),
.B(n_697),
.C(n_672),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_861),
.A2(n_571),
.B(n_636),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_SL g869 ( 
.A1(n_714),
.A2(n_702),
.B(n_588),
.C(n_584),
.Y(n_869)
);

INVx1_ASAP7_75t_SL g870 ( 
.A(n_834),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_709),
.A2(n_613),
.B1(n_612),
.B2(n_569),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_794),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_785),
.B(n_623),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_839),
.B(n_595),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_787),
.B(n_612),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_721),
.B(n_594),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_710),
.A2(n_703),
.B(n_648),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_775),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_853),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_743),
.B(n_612),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_711),
.A2(n_648),
.B(n_668),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_711),
.A2(n_668),
.B(n_703),
.Y(n_882)
);

OAI321xp33_ASAP7_75t_L g883 ( 
.A1(n_800),
.A2(n_594),
.A3(n_699),
.B1(n_705),
.B2(n_704),
.C(n_696),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_814),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_718),
.B(n_623),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_713),
.B(n_594),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_797),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_726),
.A2(n_672),
.B(n_584),
.C(n_586),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_722),
.A2(n_668),
.B(n_703),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_799),
.Y(n_890)
);

AOI221xp5_ASAP7_75t_L g891 ( 
.A1(n_832),
.A2(n_693),
.B1(n_692),
.B2(n_667),
.C(n_705),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_720),
.B(n_679),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_727),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_730),
.B(n_679),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_732),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_741),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_731),
.B(n_679),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_746),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_816),
.B(n_665),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_761),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_823),
.B(n_699),
.C(n_652),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_799),
.A2(n_602),
.B(n_586),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_781),
.A2(n_588),
.B(n_602),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_747),
.A2(n_665),
.B1(n_570),
.B2(n_704),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_765),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_857),
.Y(n_906)
);

NOR2x1p5_ASAP7_75t_SL g907 ( 
.A(n_802),
.B(n_644),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_792),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_734),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_749),
.B(n_665),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_742),
.B(n_698),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_842),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_806),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_752),
.B(n_570),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_857),
.Y(n_915)
);

INVx11_ASAP7_75t_L g916 ( 
.A(n_778),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_724),
.A2(n_657),
.B(n_642),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_751),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_819),
.B(n_601),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_802),
.A2(n_642),
.B(n_657),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_723),
.A2(n_658),
.B1(n_644),
.B2(n_683),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_819),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_836),
.A2(n_657),
.B(n_653),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_753),
.B(n_653),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_808),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_714),
.A2(n_701),
.B(n_700),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_815),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_728),
.Y(n_928)
);

CKINVDCx10_ASAP7_75t_R g929 ( 
.A(n_825),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_723),
.B(n_683),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_833),
.B(n_662),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_715),
.A2(n_701),
.B(n_700),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_728),
.A2(n_662),
.B(n_658),
.Y(n_933)
);

NOR3xp33_ASAP7_75t_L g934 ( 
.A(n_764),
.B(n_782),
.C(n_798),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_715),
.A2(n_745),
.B(n_729),
.Y(n_935)
);

BUFx12f_ASAP7_75t_L g936 ( 
.A(n_790),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_858),
.B(n_601),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_738),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_810),
.A2(n_570),
.B1(n_601),
.B2(n_238),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_745),
.A2(n_601),
.B(n_641),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_735),
.A2(n_641),
.B1(n_654),
.B2(n_297),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_848),
.A2(n_592),
.B1(n_242),
.B2(n_273),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_762),
.A2(n_641),
.B(n_654),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_827),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_766),
.A2(n_654),
.B(n_274),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_852),
.A2(n_270),
.B(n_289),
.C(n_277),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_791),
.B(n_592),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_766),
.A2(n_654),
.B(n_275),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_775),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_767),
.A2(n_788),
.B(n_769),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_826),
.A2(n_781),
.B(n_841),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_759),
.B(n_30),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_859),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_767),
.A2(n_265),
.B(n_247),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_769),
.A2(n_245),
.B(n_243),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_795),
.B(n_592),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_819),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_788),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_770),
.B(n_771),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_772),
.B(n_30),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_756),
.B(n_35),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_756),
.B(n_35),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_803),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_847),
.B(n_36),
.Y(n_964)
);

NAND2xp33_ASAP7_75t_L g965 ( 
.A(n_775),
.B(n_36),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_716),
.B(n_41),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_811),
.A2(n_79),
.B(n_160),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_821),
.A2(n_77),
.B(n_157),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_775),
.B(n_41),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_805),
.B(n_44),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_725),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_773),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_736),
.A2(n_760),
.B(n_712),
.C(n_831),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_856),
.B(n_733),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_736),
.A2(n_52),
.B(n_53),
.C(n_55),
.Y(n_975)
);

AOI21x1_ASAP7_75t_L g976 ( 
.A1(n_837),
.A2(n_93),
.B(n_131),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_754),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_719),
.A2(n_58),
.B1(n_62),
.B2(n_108),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_796),
.A2(n_109),
.B1(n_173),
.B2(n_801),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_774),
.B(n_817),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_783),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_835),
.A2(n_840),
.B(n_849),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_840),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_SL g984 ( 
.A(n_805),
.B(n_854),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_783),
.B(n_849),
.Y(n_985)
);

AOI21x1_ASAP7_75t_L g986 ( 
.A1(n_837),
.A2(n_845),
.B(n_844),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_783),
.B(n_860),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_844),
.A2(n_845),
.B(n_793),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_830),
.A2(n_846),
.B(n_758),
.C(n_841),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_784),
.B(n_813),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_779),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_717),
.A2(n_744),
.B1(n_739),
.B2(n_740),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_804),
.B(n_809),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_779),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_717),
.A2(n_737),
.B1(n_739),
.B2(n_740),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_851),
.B(n_855),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_812),
.B(n_843),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_829),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_862),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_824),
.A2(n_828),
.B(n_750),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_780),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_750),
.A2(n_755),
.B(n_793),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_755),
.A2(n_768),
.B(n_777),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_768),
.A2(n_777),
.B(n_807),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_789),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_748),
.A2(n_850),
.B(n_838),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_850),
.B(n_757),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_789),
.B(n_807),
.Y(n_1008)
);

INVx11_ASAP7_75t_L g1009 ( 
.A(n_853),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_820),
.B(n_579),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_794),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_820),
.A2(n_786),
.B(n_818),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_820),
.B(n_579),
.Y(n_1013)
);

AO21x1_ASAP7_75t_L g1014 ( 
.A1(n_826),
.A2(n_781),
.B(n_715),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_820),
.A2(n_786),
.B(n_818),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_776),
.B(n_568),
.Y(n_1016)
);

OAI321xp33_ASAP7_75t_L g1017 ( 
.A1(n_800),
.A2(n_523),
.A3(n_848),
.B1(n_390),
.B2(n_610),
.C(n_712),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_820),
.A2(n_786),
.B(n_818),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_878),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_878),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_1001),
.B(n_922),
.Y(n_1023)
);

AO31x2_ASAP7_75t_L g1024 ( 
.A1(n_1014),
.A2(n_951),
.A3(n_935),
.B(n_930),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_903),
.A2(n_982),
.B(n_950),
.Y(n_1025)
);

OAI22x1_ASAP7_75t_L g1026 ( 
.A1(n_876),
.A2(n_944),
.B1(n_992),
.B2(n_864),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1016),
.B(n_876),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_866),
.B(n_873),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_952),
.A2(n_973),
.B(n_966),
.C(n_989),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_980),
.B(n_990),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_993),
.B(n_997),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_878),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_918),
.B(n_984),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_940),
.A2(n_986),
.B(n_932),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_998),
.B(n_959),
.Y(n_1035)
);

AO21x1_ASAP7_75t_L g1036 ( 
.A1(n_1000),
.A2(n_996),
.B(n_1006),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_892),
.A2(n_897),
.B(n_894),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_872),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_958),
.B(n_893),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_926),
.A2(n_923),
.B(n_902),
.Y(n_1040)
);

AOI21x1_ASAP7_75t_L g1041 ( 
.A1(n_985),
.A2(n_988),
.B(n_956),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_910),
.B(n_875),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_952),
.A2(n_973),
.B(n_966),
.C(n_989),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_870),
.B(n_885),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_934),
.A2(n_918),
.B1(n_871),
.B2(n_910),
.Y(n_1045)
);

OAI22x1_ASAP7_75t_L g1046 ( 
.A1(n_995),
.A2(n_991),
.B1(n_904),
.B2(n_970),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_867),
.A2(n_888),
.B(n_882),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_1017),
.B(n_909),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_SL g1049 ( 
.A1(n_880),
.A2(n_886),
.B(n_1002),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_895),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_888),
.A2(n_889),
.B(n_881),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_909),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_999),
.B(n_896),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_898),
.B(n_900),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_937),
.A2(n_877),
.B(n_917),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_933),
.A2(n_1004),
.B(n_943),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_905),
.B(n_908),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_947),
.A2(n_1007),
.B(n_919),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_920),
.A2(n_869),
.B(n_868),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_879),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_967),
.A2(n_968),
.B(n_919),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_878),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_934),
.A2(n_974),
.B(n_960),
.C(n_996),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_SL g1064 ( 
.A1(n_972),
.A2(n_970),
.B(n_977),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_SL g1065 ( 
.A1(n_922),
.A2(n_957),
.B(n_1001),
.Y(n_1065)
);

AOI222xp33_ASAP7_75t_L g1066 ( 
.A1(n_972),
.A2(n_891),
.B1(n_883),
.B2(n_971),
.C1(n_936),
.C2(n_942),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_899),
.B(n_884),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_874),
.B(n_938),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_976),
.A2(n_1003),
.B(n_921),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_916),
.B(n_884),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_945),
.A2(n_948),
.B(n_924),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_931),
.A2(n_865),
.B(n_946),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_L g1073 ( 
.A(n_901),
.B(n_874),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_994),
.B(n_1001),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_921),
.A2(n_983),
.B(n_963),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_912),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_SL g1077 ( 
.A1(n_961),
.A2(n_962),
.B(n_946),
.C(n_969),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_961),
.A2(n_962),
.B(n_914),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_913),
.Y(n_1079)
);

AO32x2_ASAP7_75t_L g1080 ( 
.A1(n_941),
.A2(n_975),
.A3(n_907),
.B1(n_969),
.B2(n_965),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_949),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_925),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_927),
.A2(n_979),
.B1(n_975),
.B2(n_942),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_964),
.B(n_953),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_987),
.A2(n_928),
.B(n_911),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_987),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_957),
.B(n_981),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_863),
.A2(n_906),
.B(n_915),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_887),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_863),
.A2(n_906),
.B(n_915),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_890),
.B(n_1011),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_1009),
.Y(n_1092)
);

INVx5_ASAP7_75t_L g1093 ( 
.A(n_949),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_955),
.A2(n_1008),
.B(n_978),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1008),
.B(n_949),
.Y(n_1095)
);

OAI22x1_ASAP7_75t_L g1096 ( 
.A1(n_1005),
.A2(n_939),
.B1(n_929),
.B2(n_981),
.Y(n_1096)
);

AOI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_981),
.A2(n_864),
.B(n_952),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_954),
.B(n_1016),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_903),
.A2(n_935),
.B(n_982),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_944),
.B(n_814),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_864),
.A2(n_952),
.B(n_723),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_864),
.A2(n_952),
.B(n_973),
.C(n_876),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_935),
.A2(n_1015),
.B(n_1012),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_893),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_903),
.A2(n_935),
.B(n_982),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_903),
.A2(n_951),
.B(n_1000),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1014),
.A2(n_951),
.A3(n_935),
.B(n_930),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_903),
.A2(n_935),
.B(n_982),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_909),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_991),
.B(n_874),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_878),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_879),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_878),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_903),
.A2(n_935),
.B(n_982),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_864),
.A2(n_1013),
.B1(n_1010),
.B2(n_972),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1014),
.A2(n_951),
.A3(n_935),
.B(n_930),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1126)
);

NOR2xp67_ASAP7_75t_L g1127 ( 
.A(n_918),
.B(n_692),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_991),
.B(n_874),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_991),
.B(n_874),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_991),
.B(n_874),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_893),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1014),
.A2(n_951),
.A3(n_935),
.B(n_930),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_879),
.B(n_839),
.Y(n_1137)
);

AOI221x1_ASAP7_75t_L g1138 ( 
.A1(n_973),
.A2(n_864),
.B1(n_989),
.B2(n_975),
.C(n_1007),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_879),
.B(n_839),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_903),
.A2(n_935),
.B(n_982),
.Y(n_1142)
);

INVx4_ASAP7_75t_SL g1143 ( 
.A(n_878),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_909),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1009),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_903),
.A2(n_935),
.B(n_982),
.Y(n_1147)
);

AOI21x1_ASAP7_75t_L g1148 ( 
.A1(n_903),
.A2(n_951),
.B(n_1000),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_935),
.A2(n_1015),
.B(n_1012),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1012),
.A2(n_1018),
.B(n_1015),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_893),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1014),
.A2(n_951),
.A3(n_935),
.B(n_930),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_918),
.B(n_692),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_L g1155 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_893),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_870),
.B(n_834),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_903),
.A2(n_935),
.B(n_982),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1016),
.B(n_870),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_878),
.Y(n_1160)
);

INVx3_ASAP7_75t_SL g1161 ( 
.A(n_1092),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1157),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1050),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1022),
.A2(n_1111),
.B(n_1109),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_1020),
.B(n_1093),
.Y(n_1165)
);

AOI21xp33_ASAP7_75t_SL g1166 ( 
.A1(n_1124),
.A2(n_1026),
.B(n_1045),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1120),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1146),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1028),
.B(n_1102),
.Y(n_1169)
);

CKINVDCx20_ASAP7_75t_R g1170 ( 
.A(n_1060),
.Y(n_1170)
);

INVx3_ASAP7_75t_SL g1171 ( 
.A(n_1068),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1020),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1020),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1044),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1079),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1038),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1082),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1124),
.B(n_1102),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1107),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1066),
.A2(n_1101),
.B1(n_1048),
.B2(n_1033),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1159),
.B(n_1052),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1106),
.A2(n_1150),
.B(n_1119),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1104),
.B(n_1105),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1093),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1134),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1114),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1076),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1152),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1019),
.B(n_1126),
.Y(n_1189)
);

O2A1O1Ixp5_ASAP7_75t_SL g1190 ( 
.A1(n_1101),
.A2(n_1097),
.B(n_1150),
.C(n_1106),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1116),
.A2(n_1140),
.B(n_1122),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1104),
.B(n_1105),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1056),
.A2(n_1025),
.B(n_1034),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1141),
.A2(n_1145),
.B(n_1151),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1117),
.B(n_1129),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1029),
.A2(n_1043),
.B(n_1155),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1093),
.B(n_1115),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1156),
.Y(n_1198)
);

AO32x2_ASAP7_75t_L g1199 ( 
.A1(n_1083),
.A2(n_1138),
.A3(n_1112),
.B1(n_1024),
.B2(n_1135),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1054),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1064),
.A2(n_1066),
.B1(n_1027),
.B2(n_1117),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1057),
.Y(n_1202)
);

NOR2x1p5_ASAP7_75t_SL g1203 ( 
.A(n_1110),
.B(n_1148),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1039),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1094),
.A2(n_1063),
.B(n_1030),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1128),
.B(n_1130),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_L g1207 ( 
.A(n_1131),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1042),
.B(n_1031),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1031),
.B(n_1132),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1039),
.Y(n_1210)
);

INVx8_ASAP7_75t_L g1211 ( 
.A(n_1137),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1064),
.A2(n_1133),
.B1(n_1136),
.B2(n_1149),
.Y(n_1212)
);

OR2x2_ASAP7_75t_SL g1213 ( 
.A(n_1035),
.B(n_1053),
.Y(n_1213)
);

INVx4_ASAP7_75t_L g1214 ( 
.A(n_1143),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1089),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_1065),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1084),
.A2(n_1098),
.B1(n_1144),
.B2(n_1078),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1070),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1061),
.A2(n_1037),
.B(n_1051),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1067),
.B(n_1154),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1095),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1072),
.A2(n_1069),
.B(n_1047),
.C(n_1095),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1074),
.B(n_1091),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1100),
.B(n_1073),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1137),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1077),
.A2(n_1049),
.B(n_1072),
.C(n_1047),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1139),
.B(n_1127),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1032),
.Y(n_1228)
);

BUFx10_ASAP7_75t_L g1229 ( 
.A(n_1032),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1143),
.B(n_1139),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1046),
.B(n_1074),
.Y(n_1231)
);

BUFx8_ASAP7_75t_L g1232 ( 
.A(n_1032),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1021),
.B(n_1081),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1062),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1075),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1086),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1062),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1062),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1160),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1096),
.A2(n_1036),
.B1(n_1121),
.B2(n_1118),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1021),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1081),
.B(n_1121),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1143),
.B(n_1118),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1160),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1160),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1023),
.Y(n_1246)
);

BUFx4_ASAP7_75t_SL g1247 ( 
.A(n_1080),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_L g1248 ( 
.A(n_1023),
.B(n_1087),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1085),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1080),
.B(n_1024),
.Y(n_1250)
);

BUFx8_ASAP7_75t_L g1251 ( 
.A(n_1080),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1040),
.A2(n_1058),
.B(n_1090),
.Y(n_1252)
);

INVx8_ASAP7_75t_L g1253 ( 
.A(n_1088),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1071),
.A2(n_1041),
.B1(n_1125),
.B2(n_1135),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1099),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1125),
.B(n_1153),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1108),
.A2(n_1113),
.B1(n_1123),
.B2(n_1142),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1147),
.B(n_1158),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1124),
.A2(n_1101),
.B1(n_1048),
.B2(n_864),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1019),
.B(n_1126),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1115),
.B(n_1128),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1020),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1159),
.B(n_870),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1020),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1101),
.A2(n_864),
.B(n_1103),
.C(n_876),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1159),
.B(n_870),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_L g1267 ( 
.A(n_1020),
.B(n_1093),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1120),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1106),
.A2(n_1150),
.B(n_1109),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1124),
.A2(n_1101),
.B1(n_1048),
.B2(n_864),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1124),
.B(n_1102),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1115),
.B(n_1128),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1020),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1050),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1157),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1050),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1050),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1050),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1101),
.A2(n_864),
.B(n_1103),
.C(n_876),
.Y(n_1279)
);

INVx5_ASAP7_75t_L g1280 ( 
.A(n_1137),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1120),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1159),
.B(n_870),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1020),
.Y(n_1283)
);

OA21x2_ASAP7_75t_L g1284 ( 
.A1(n_1106),
.A2(n_1150),
.B(n_1109),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1020),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1028),
.B(n_944),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1157),
.B(n_870),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1092),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1159),
.B(n_870),
.Y(n_1289)
);

AND2x6_ASAP7_75t_L g1290 ( 
.A(n_1074),
.B(n_1086),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1124),
.B(n_1102),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1066),
.A2(n_723),
.B1(n_708),
.B2(n_1101),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1050),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1092),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1022),
.A2(n_1111),
.B(n_1109),
.Y(n_1295)
);

CKINVDCx8_ASAP7_75t_R g1296 ( 
.A(n_1115),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1159),
.B(n_870),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1092),
.Y(n_1298)
);

OR2x6_ASAP7_75t_L g1299 ( 
.A(n_1137),
.B(n_1139),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1022),
.A2(n_1111),
.B(n_1109),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1022),
.A2(n_1111),
.B(n_1109),
.Y(n_1301)
);

INVx8_ASAP7_75t_L g1302 ( 
.A(n_1211),
.Y(n_1302)
);

INVx4_ASAP7_75t_L g1303 ( 
.A(n_1214),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1292),
.A2(n_1180),
.B1(n_1201),
.B2(n_1251),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1235),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1201),
.A2(n_1251),
.B1(n_1212),
.B2(n_1259),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1259),
.A2(n_1270),
.B(n_1254),
.Y(n_1307)
);

INVx5_ASAP7_75t_L g1308 ( 
.A(n_1214),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1163),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1175),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1177),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1179),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1181),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_SL g1314 ( 
.A1(n_1205),
.A2(n_1196),
.B(n_1178),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1270),
.A2(n_1205),
.B1(n_1174),
.B2(n_1271),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1169),
.B(n_1195),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1232),
.Y(n_1317)
);

INVx3_ASAP7_75t_SL g1318 ( 
.A(n_1294),
.Y(n_1318)
);

AO21x1_ASAP7_75t_L g1319 ( 
.A1(n_1166),
.A2(n_1226),
.B(n_1178),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1230),
.B(n_1243),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1185),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1211),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1188),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1247),
.A2(n_1291),
.B1(n_1271),
.B2(n_1217),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1198),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1265),
.A2(n_1279),
.B1(n_1291),
.B2(n_1166),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1230),
.B(n_1243),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1274),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1276),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1170),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1298),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1277),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1278),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1232),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1209),
.B(n_1183),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1293),
.Y(n_1336)
);

BUFx2_ASAP7_75t_R g1337 ( 
.A(n_1296),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1215),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1295),
.A2(n_1301),
.B(n_1300),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1286),
.A2(n_1224),
.B1(n_1208),
.B2(n_1209),
.Y(n_1340)
);

BUFx8_ASAP7_75t_L g1341 ( 
.A(n_1268),
.Y(n_1341)
);

BUFx10_ASAP7_75t_L g1342 ( 
.A(n_1218),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1174),
.A2(n_1162),
.B1(n_1231),
.B2(n_1263),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1200),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1256),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1202),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1221),
.B(n_1250),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1199),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1254),
.A2(n_1219),
.B(n_1222),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1204),
.B(n_1210),
.Y(n_1350)
);

BUFx5_ASAP7_75t_L g1351 ( 
.A(n_1249),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1176),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1281),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1161),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1253),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1211),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1217),
.A2(n_1192),
.B1(n_1183),
.B2(n_1162),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1192),
.B(n_1189),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1199),
.B(n_1190),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1260),
.B(n_1240),
.Y(n_1360)
);

INVx3_ASAP7_75t_SL g1361 ( 
.A(n_1171),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1182),
.B(n_1269),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1220),
.A2(n_1289),
.B1(n_1282),
.B2(n_1297),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1239),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1213),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1223),
.Y(n_1366)
);

CKINVDCx11_ASAP7_75t_R g1367 ( 
.A(n_1288),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1261),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1284),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1186),
.Y(n_1370)
);

NOR2x1_ASAP7_75t_R g1371 ( 
.A(n_1168),
.B(n_1187),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1266),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1223),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1287),
.A2(n_1275),
.B1(n_1290),
.B2(n_1236),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1241),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1252),
.A2(n_1257),
.B(n_1193),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1239),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_1167),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1280),
.A2(n_1290),
.B1(n_1207),
.B2(n_1225),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1284),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1238),
.B(n_1228),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1233),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1234),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1233),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1261),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1272),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1242),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1245),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1242),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1253),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1299),
.A2(n_1206),
.B1(n_1227),
.B2(n_1197),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1253),
.Y(n_1392)
);

BUFx2_ASAP7_75t_R g1393 ( 
.A(n_1244),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1246),
.A2(n_1248),
.B1(n_1285),
.B2(n_1262),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1262),
.A2(n_1285),
.B1(n_1283),
.B2(n_1273),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1229),
.Y(n_1396)
);

OAI21xp33_ASAP7_75t_L g1397 ( 
.A1(n_1203),
.A2(n_1255),
.B(n_1258),
.Y(n_1397)
);

AO21x1_ASAP7_75t_L g1398 ( 
.A1(n_1255),
.A2(n_1238),
.B(n_1239),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1264),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1237),
.B(n_1184),
.Y(n_1400)
);

BUFx12f_ASAP7_75t_L g1401 ( 
.A(n_1264),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1229),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1237),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1172),
.A2(n_1173),
.B(n_1184),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1165),
.A2(n_1267),
.B(n_1173),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1172),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1273),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1273),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1165),
.B(n_1267),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1283),
.B(n_1169),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1259),
.A2(n_1270),
.B(n_1254),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1164),
.A2(n_1194),
.B(n_1191),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1294),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1251),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1163),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1163),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1268),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1292),
.A2(n_723),
.B1(n_1066),
.B2(n_708),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1253),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1268),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1163),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1181),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1216),
.A2(n_1103),
.B(n_1043),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1262),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1163),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1259),
.B(n_1270),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1251),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1163),
.Y(n_1428)
);

BUFx10_ASAP7_75t_L g1429 ( 
.A(n_1294),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1163),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1251),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1305),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1355),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1326),
.A2(n_1426),
.B(n_1423),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1355),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1370),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1347),
.B(n_1348),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1347),
.B(n_1348),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1307),
.B(n_1411),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1307),
.B(n_1411),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1330),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1382),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1384),
.Y(n_1443)
);

AO21x1_ASAP7_75t_SL g1444 ( 
.A1(n_1306),
.A2(n_1315),
.B(n_1397),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1411),
.B(n_1359),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1387),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1390),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1389),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1359),
.B(n_1362),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1372),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1335),
.B(n_1358),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1314),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1401),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1418),
.A2(n_1324),
.B1(n_1304),
.B2(n_1340),
.Y(n_1454)
);

AOI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1339),
.A2(n_1412),
.B(n_1319),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1362),
.B(n_1350),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1351),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1350),
.B(n_1313),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1360),
.A2(n_1431),
.B1(n_1414),
.B2(n_1427),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1390),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1314),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1422),
.B(n_1309),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1310),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1311),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1312),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1321),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1369),
.A2(n_1380),
.B(n_1319),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1323),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1325),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1328),
.B(n_1329),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1351),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1332),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_SL g1473 ( 
.A(n_1337),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1333),
.B(n_1336),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1415),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1383),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1316),
.B(n_1357),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1416),
.B(n_1421),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1392),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1392),
.A2(n_1419),
.B(n_1404),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1425),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1351),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1428),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1430),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1338),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1375),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1351),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1344),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1388),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1351),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1346),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1349),
.B(n_1345),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1366),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1373),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1406),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1365),
.B(n_1431),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1398),
.A2(n_1360),
.B(n_1352),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1403),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1427),
.B(n_1381),
.Y(n_1499)
);

NAND2xp33_ASAP7_75t_R g1500 ( 
.A(n_1413),
.B(n_1405),
.Y(n_1500)
);

NOR2xp67_ASAP7_75t_L g1501 ( 
.A(n_1308),
.B(n_1408),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1376),
.Y(n_1502)
);

OR2x6_ASAP7_75t_L g1503 ( 
.A(n_1302),
.B(n_1409),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1376),
.Y(n_1504)
);

AO21x2_ASAP7_75t_L g1505 ( 
.A1(n_1376),
.A2(n_1410),
.B(n_1400),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1381),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1405),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1354),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1407),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1303),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1417),
.A2(n_1420),
.B(n_1394),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1320),
.B(n_1327),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1363),
.B(n_1343),
.Y(n_1513)
);

AO21x2_ASAP7_75t_L g1514 ( 
.A1(n_1320),
.A2(n_1327),
.B(n_1374),
.Y(n_1514)
);

AO21x2_ASAP7_75t_L g1515 ( 
.A1(n_1320),
.A2(n_1327),
.B(n_1391),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1408),
.B(n_1368),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1409),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1330),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1505),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1456),
.B(n_1342),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1512),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1437),
.B(n_1361),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1456),
.B(n_1342),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1437),
.B(n_1438),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1438),
.B(n_1449),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1434),
.A2(n_1378),
.B1(n_1396),
.B2(n_1402),
.C(n_1354),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1449),
.B(n_1342),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1512),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1467),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1445),
.B(n_1440),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1440),
.B(n_1353),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1454),
.A2(n_1378),
.B1(n_1361),
.B2(n_1396),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1442),
.B(n_1424),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1512),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1432),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1505),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1498),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1439),
.B(n_1317),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1505),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1457),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1506),
.B(n_1317),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1436),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1492),
.B(n_1334),
.Y(n_1543)
);

OAI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1477),
.A2(n_1302),
.B1(n_1386),
.B2(n_1385),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1452),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1492),
.B(n_1334),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1480),
.B(n_1356),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1512),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1452),
.B(n_1377),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1442),
.B(n_1364),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1461),
.B(n_1364),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1480),
.B(n_1457),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1461),
.B(n_1303),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1443),
.B(n_1341),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1458),
.B(n_1399),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1458),
.B(n_1399),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1502),
.B(n_1318),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1502),
.B(n_1504),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1511),
.A2(n_1379),
.B1(n_1356),
.B2(n_1322),
.C(n_1395),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1435),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1443),
.B(n_1341),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1435),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1504),
.B(n_1318),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1495),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1455),
.B(n_1429),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1508),
.B(n_1371),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1446),
.B(n_1341),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1446),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1568),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1542),
.B(n_1450),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1542),
.B(n_1462),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1532),
.A2(n_1559),
.B1(n_1500),
.B2(n_1526),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1537),
.B(n_1462),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_L g1574 ( 
.A(n_1557),
.B(n_1563),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1526),
.B(n_1495),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1565),
.B(n_1435),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1532),
.A2(n_1459),
.B1(n_1441),
.B2(n_1518),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1527),
.B(n_1499),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1537),
.B(n_1476),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1527),
.B(n_1471),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1564),
.B(n_1489),
.Y(n_1581)
);

NOR3xp33_ASAP7_75t_L g1582 ( 
.A(n_1565),
.B(n_1563),
.C(n_1557),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1564),
.B(n_1451),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1568),
.B(n_1470),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1565),
.B(n_1560),
.Y(n_1585)
);

AOI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1530),
.A2(n_1491),
.B1(n_1488),
.B2(n_1494),
.C(n_1493),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1527),
.B(n_1474),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1559),
.A2(n_1529),
.B(n_1538),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1530),
.B(n_1474),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1522),
.A2(n_1473),
.B1(n_1496),
.B2(n_1503),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1522),
.A2(n_1503),
.B1(n_1402),
.B2(n_1510),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1530),
.A2(n_1488),
.B1(n_1491),
.B2(n_1494),
.C(n_1493),
.Y(n_1592)
);

NOR3xp33_ASAP7_75t_L g1593 ( 
.A(n_1554),
.B(n_1509),
.C(n_1447),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1525),
.B(n_1471),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1560),
.B(n_1562),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_L g1596 ( 
.A(n_1554),
.B(n_1509),
.C(n_1433),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1555),
.B(n_1478),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1538),
.A2(n_1444),
.B1(n_1513),
.B2(n_1514),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1529),
.A2(n_1483),
.B1(n_1472),
.B2(n_1463),
.C(n_1475),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_L g1600 ( 
.A(n_1545),
.B(n_1448),
.C(n_1486),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1555),
.B(n_1448),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1525),
.B(n_1482),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1560),
.B(n_1435),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1556),
.B(n_1463),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1520),
.B(n_1482),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1556),
.B(n_1464),
.Y(n_1606)
);

NOR3xp33_ASAP7_75t_L g1607 ( 
.A(n_1561),
.B(n_1460),
.C(n_1433),
.Y(n_1607)
);

NAND3xp33_ASAP7_75t_L g1608 ( 
.A(n_1545),
.B(n_1486),
.C(n_1507),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_L g1609 ( 
.A(n_1538),
.B(n_1507),
.C(n_1485),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1523),
.B(n_1487),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1550),
.B(n_1533),
.C(n_1549),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1522),
.A2(n_1503),
.B1(n_1510),
.B2(n_1453),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1519),
.A2(n_1536),
.B1(n_1539),
.B2(n_1466),
.C(n_1468),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1521),
.B(n_1517),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1523),
.B(n_1487),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1556),
.B(n_1465),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1531),
.A2(n_1497),
.B1(n_1514),
.B2(n_1515),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1524),
.B(n_1465),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1562),
.B(n_1479),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1523),
.B(n_1466),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1543),
.B(n_1490),
.Y(n_1621)
);

AND4x1_ASAP7_75t_L g1622 ( 
.A(n_1566),
.B(n_1367),
.C(n_1516),
.D(n_1331),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1567),
.B(n_1367),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1569),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1583),
.B(n_1561),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1574),
.B(n_1552),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1594),
.B(n_1552),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1614),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1608),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1584),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1604),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1594),
.B(n_1552),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1618),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1602),
.B(n_1552),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1552),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1582),
.B(n_1540),
.Y(n_1638)
);

NAND4xp25_ASAP7_75t_L g1639 ( 
.A(n_1572),
.B(n_1567),
.C(n_1553),
.D(n_1551),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1598),
.A2(n_1444),
.B1(n_1531),
.B2(n_1514),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1578),
.B(n_1521),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1606),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1578),
.B(n_1528),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1586),
.B(n_1558),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1616),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1609),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1621),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1592),
.B(n_1558),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1601),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1589),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1571),
.B(n_1550),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1599),
.B(n_1558),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1595),
.B(n_1534),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1570),
.B(n_1541),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1611),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1620),
.Y(n_1656)
);

AND2x2_ASAP7_75t_SL g1657 ( 
.A(n_1593),
.B(n_1531),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1597),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1613),
.B(n_1535),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1588),
.A2(n_1544),
.B(n_1533),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1575),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1596),
.B(n_1535),
.Y(n_1662)
);

NAND2x1_ASAP7_75t_L g1663 ( 
.A(n_1580),
.B(n_1547),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1579),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1614),
.Y(n_1665)
);

INVx4_ASAP7_75t_L g1666 ( 
.A(n_1614),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1585),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1585),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1663),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1625),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1646),
.B(n_1503),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1646),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1657),
.A2(n_1661),
.B1(n_1652),
.B2(n_1644),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1657),
.Y(n_1674)
);

AOI211xp5_ASAP7_75t_L g1675 ( 
.A1(n_1639),
.A2(n_1577),
.B(n_1575),
.C(n_1590),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1625),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1657),
.B(n_1580),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1629),
.B(n_1573),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1629),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1656),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1656),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1657),
.B(n_1605),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1627),
.B(n_1548),
.Y(n_1683)
);

NAND2x1_ASAP7_75t_SL g1684 ( 
.A(n_1631),
.B(n_1543),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1652),
.B(n_1581),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1655),
.B(n_1587),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1642),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1642),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1631),
.B(n_1468),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1638),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1631),
.B(n_1469),
.Y(n_1691)
);

OA211x2_ASAP7_75t_L g1692 ( 
.A1(n_1663),
.A2(n_1624),
.B(n_1576),
.C(n_1623),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1666),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1646),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1655),
.B(n_1469),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1645),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1644),
.B(n_1472),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1645),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1653),
.B(n_1607),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1647),
.B(n_1605),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1633),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1647),
.B(n_1610),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1638),
.B(n_1610),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1633),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1638),
.B(n_1627),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1627),
.B(n_1630),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1649),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1648),
.B(n_1475),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1648),
.B(n_1481),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1649),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1630),
.B(n_1615),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1630),
.B(n_1615),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1686),
.B(n_1664),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1701),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1678),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1677),
.B(n_1661),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1679),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1674),
.B(n_1666),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1686),
.B(n_1664),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1679),
.B(n_1659),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1677),
.B(n_1666),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1672),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1701),
.Y(n_1723)
);

AND2x4_ASAP7_75t_SL g1724 ( 
.A(n_1706),
.B(n_1653),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1695),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1695),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1689),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1689),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1691),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1678),
.B(n_1659),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1685),
.B(n_1651),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1701),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1691),
.Y(n_1733)
);

OAI21xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1673),
.A2(n_1639),
.B(n_1666),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1670),
.Y(n_1735)
);

INVx1_ASAP7_75t_SL g1736 ( 
.A(n_1674),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1674),
.B(n_1666),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1670),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1673),
.A2(n_1643),
.B(n_1641),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1704),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1685),
.B(n_1651),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1704),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1669),
.B(n_1653),
.Y(n_1743)
);

OR2x2_ASAP7_75t_SL g1744 ( 
.A(n_1672),
.B(n_1667),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1697),
.B(n_1651),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1676),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1697),
.B(n_1654),
.Y(n_1747)
);

NOR2xp67_ASAP7_75t_L g1748 ( 
.A(n_1669),
.B(n_1667),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1676),
.Y(n_1749)
);

NAND2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1669),
.B(n_1622),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1682),
.B(n_1667),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1672),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1682),
.B(n_1668),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1675),
.A2(n_1640),
.B1(n_1617),
.B2(n_1660),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1694),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1694),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1690),
.B(n_1653),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1700),
.B(n_1668),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1724),
.B(n_1690),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1720),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1717),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1754),
.A2(n_1694),
.B1(n_1640),
.B2(n_1660),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1717),
.B(n_1730),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1736),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1744),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1715),
.B(n_1731),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1750),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1750),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1741),
.B(n_1708),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1735),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1724),
.B(n_1757),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1757),
.B(n_1705),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1734),
.A2(n_1675),
.B1(n_1671),
.B2(n_1708),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1725),
.B(n_1709),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1757),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1716),
.B(n_1705),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1738),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1716),
.A2(n_1671),
.B1(n_1709),
.B2(n_1692),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1726),
.B(n_1700),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1713),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1719),
.B(n_1747),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1746),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1745),
.B(n_1680),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1727),
.B(n_1728),
.Y(n_1784)
);

AND2x2_ASAP7_75t_SL g1785 ( 
.A(n_1718),
.B(n_1706),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1729),
.B(n_1702),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1733),
.B(n_1702),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1718),
.Y(n_1788)
);

NOR2x1_ASAP7_75t_L g1789 ( 
.A(n_1748),
.B(n_1693),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1749),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1714),
.Y(n_1791)
);

NAND4xp75_ASAP7_75t_L g1792 ( 
.A(n_1739),
.B(n_1692),
.C(n_1699),
.D(n_1703),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1758),
.B(n_1680),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1714),
.Y(n_1794)
);

INVx1_ASAP7_75t_SL g1795 ( 
.A(n_1718),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1758),
.B(n_1681),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1785),
.B(n_1751),
.Y(n_1797)
);

OAI31xp33_ASAP7_75t_L g1798 ( 
.A1(n_1762),
.A2(n_1722),
.A3(n_1755),
.B(n_1752),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1792),
.A2(n_1773),
.B1(n_1762),
.B2(n_1778),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1765),
.A2(n_1671),
.B1(n_1722),
.B2(n_1756),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1761),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1759),
.A2(n_1743),
.B1(n_1703),
.B2(n_1737),
.Y(n_1802)
);

NOR2x1_ASAP7_75t_L g1803 ( 
.A(n_1767),
.B(n_1737),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1763),
.A2(n_1742),
.B1(n_1740),
.B2(n_1723),
.C(n_1732),
.Y(n_1804)
);

AOI221x1_ASAP7_75t_L g1805 ( 
.A1(n_1763),
.A2(n_1737),
.B1(n_1742),
.B2(n_1740),
.C(n_1723),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1764),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1770),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1768),
.A2(n_1662),
.B(n_1751),
.Y(n_1808)
);

OAI21xp33_ASAP7_75t_SL g1809 ( 
.A1(n_1785),
.A2(n_1721),
.B(n_1684),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1777),
.Y(n_1810)
);

NAND3x2_ASAP7_75t_L g1811 ( 
.A(n_1771),
.B(n_1743),
.C(n_1721),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1788),
.Y(n_1812)
);

OAI321xp33_ASAP7_75t_L g1813 ( 
.A1(n_1765),
.A2(n_1671),
.A3(n_1753),
.B1(n_1732),
.B2(n_1544),
.C(n_1536),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1782),
.Y(n_1814)
);

CKINVDCx14_ASAP7_75t_R g1815 ( 
.A(n_1771),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1790),
.Y(n_1816)
);

AO22x1_ASAP7_75t_L g1817 ( 
.A1(n_1759),
.A2(n_1743),
.B1(n_1753),
.B2(n_1683),
.Y(n_1817)
);

O2A1O1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1760),
.A2(n_1662),
.B(n_1671),
.C(n_1668),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1781),
.Y(n_1819)
);

OAI221xp5_ASAP7_75t_L g1820 ( 
.A1(n_1766),
.A2(n_1684),
.B1(n_1704),
.B2(n_1710),
.C(n_1707),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1784),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1772),
.B(n_1711),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1772),
.B(n_1711),
.Y(n_1823)
);

AO22x1_ASAP7_75t_L g1824 ( 
.A1(n_1759),
.A2(n_1683),
.B1(n_1693),
.B2(n_1712),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1806),
.B(n_1780),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1806),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1799),
.A2(n_1774),
.B1(n_1793),
.B2(n_1794),
.C(n_1791),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1815),
.B(n_1775),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1797),
.Y(n_1829)
);

INVxp67_ASAP7_75t_SL g1830 ( 
.A(n_1801),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1819),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1815),
.B(n_1775),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1812),
.B(n_1776),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1800),
.A2(n_1776),
.B1(n_1794),
.B2(n_1791),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1821),
.B(n_1779),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1803),
.B(n_1795),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1808),
.B(n_1769),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1808),
.B(n_1786),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1822),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1823),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1807),
.B(n_1796),
.Y(n_1841)
);

NOR3xp33_ASAP7_75t_L g1842 ( 
.A(n_1804),
.B(n_1813),
.C(n_1809),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1810),
.Y(n_1843)
);

CKINVDCx16_ASAP7_75t_R g1844 ( 
.A(n_1802),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1817),
.B(n_1787),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1826),
.A2(n_1805),
.B(n_1798),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1837),
.A2(n_1820),
.B1(n_1796),
.B2(n_1783),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1826),
.B(n_1814),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_SL g1849 ( 
.A(n_1832),
.B(n_1413),
.Y(n_1849)
);

OAI211xp5_ASAP7_75t_L g1850 ( 
.A1(n_1842),
.A2(n_1811),
.B(n_1816),
.C(n_1789),
.Y(n_1850)
);

AOI21x1_ASAP7_75t_L g1851 ( 
.A1(n_1836),
.A2(n_1824),
.B(n_1784),
.Y(n_1851)
);

OAI222xp33_ASAP7_75t_L g1852 ( 
.A1(n_1838),
.A2(n_1818),
.B1(n_1783),
.B2(n_1519),
.C1(n_1539),
.C2(n_1687),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1844),
.B(n_1331),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1842),
.A2(n_1818),
.B(n_1687),
.Y(n_1854)
);

OAI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1834),
.A2(n_1681),
.B1(n_1710),
.B2(n_1707),
.C(n_1698),
.Y(n_1855)
);

OAI21xp33_ASAP7_75t_SL g1856 ( 
.A1(n_1830),
.A2(n_1712),
.B(n_1693),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1839),
.B(n_1688),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1825),
.B(n_1688),
.Y(n_1858)
);

NAND4xp25_ASAP7_75t_L g1859 ( 
.A(n_1846),
.B(n_1832),
.C(n_1828),
.D(n_1833),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1853),
.B(n_1839),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1848),
.B(n_1840),
.Y(n_1861)
);

OAI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1851),
.A2(n_1830),
.B(n_1836),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1849),
.B(n_1829),
.Y(n_1863)
);

NOR2x1p5_ASAP7_75t_SL g1864 ( 
.A(n_1858),
.B(n_1829),
.Y(n_1864)
);

NAND4xp25_ASAP7_75t_L g1865 ( 
.A(n_1850),
.B(n_1831),
.C(n_1827),
.D(n_1845),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1856),
.B(n_1841),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1854),
.B(n_1843),
.C(n_1835),
.Y(n_1867)
);

NOR3xp33_ASAP7_75t_L g1868 ( 
.A(n_1852),
.B(n_1453),
.C(n_1696),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1857),
.B(n_1626),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1852),
.A2(n_1698),
.B(n_1696),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1863),
.B(n_1855),
.Y(n_1871)
);

O2A1O1Ixp33_ASAP7_75t_SL g1872 ( 
.A1(n_1862),
.A2(n_1847),
.B(n_1693),
.C(n_1429),
.Y(n_1872)
);

NOR2x1_ASAP7_75t_L g1873 ( 
.A(n_1865),
.B(n_1429),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1860),
.B(n_1628),
.Y(n_1874)
);

AND3x1_ASAP7_75t_L g1875 ( 
.A(n_1866),
.B(n_1626),
.C(n_1641),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_L g1876 ( 
.A(n_1867),
.B(n_1635),
.C(n_1683),
.Y(n_1876)
);

NOR3xp33_ASAP7_75t_L g1877 ( 
.A(n_1859),
.B(n_1546),
.C(n_1543),
.Y(n_1877)
);

OAI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1861),
.A2(n_1623),
.B(n_1603),
.C(n_1619),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1875),
.A2(n_1860),
.B1(n_1868),
.B2(n_1869),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1873),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1874),
.B(n_1864),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1876),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1871),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1877),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1872),
.Y(n_1885)
);

OAI21xp33_ASAP7_75t_L g1886 ( 
.A1(n_1879),
.A2(n_1878),
.B(n_1870),
.Y(n_1886)
);

NOR3xp33_ASAP7_75t_L g1887 ( 
.A(n_1883),
.B(n_1393),
.C(n_1546),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1881),
.Y(n_1888)
);

OAI21xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1882),
.A2(n_1634),
.B(n_1628),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1880),
.A2(n_1683),
.B(n_1635),
.Y(n_1890)
);

NOR2x1p5_ASAP7_75t_L g1891 ( 
.A(n_1885),
.B(n_1401),
.Y(n_1891)
);

NOR2x1_ASAP7_75t_L g1892 ( 
.A(n_1888),
.B(n_1891),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1890),
.B(n_1884),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1889),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1886),
.Y(n_1895)
);

AO22x2_ASAP7_75t_L g1896 ( 
.A1(n_1894),
.A2(n_1887),
.B1(n_1654),
.B2(n_1632),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1895),
.Y(n_1897)
);

NAND3xp33_ASAP7_75t_L g1898 ( 
.A(n_1897),
.B(n_1892),
.C(n_1893),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1898),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1898),
.B(n_1896),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1899),
.B1(n_1632),
.B2(n_1650),
.Y(n_1901)
);

OA21x2_ASAP7_75t_L g1902 ( 
.A1(n_1899),
.A2(n_1650),
.B(n_1658),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1665),
.B1(n_1633),
.B2(n_1483),
.Y(n_1903)
);

OAI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1901),
.B(n_1654),
.Y(n_1904)
);

AOI322xp5_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1665),
.A3(n_1546),
.B1(n_1628),
.B2(n_1634),
.C1(n_1636),
.C2(n_1637),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1905),
.A2(n_1665),
.B1(n_1485),
.B2(n_1484),
.Y(n_1906)
);

AOI211xp5_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1591),
.B(n_1612),
.C(n_1501),
.Y(n_1907)
);


endmodule