module fake_jpeg_1975_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx2_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_17),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_43),
.B(n_44),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g44 ( 
.A(n_23),
.B(n_1),
.CON(n_44),
.SN(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_12),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_1),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_69),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_11),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_75),
.Y(n_94)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_4),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_37),
.Y(n_82)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_78),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_75),
.B1(n_68),
.B2(n_46),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_86),
.A2(n_109),
.B1(n_85),
.B2(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_102),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_72),
.A2(n_27),
.B1(n_36),
.B2(n_28),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_115),
.B1(n_81),
.B2(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_38),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_104),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_25),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_45),
.A2(n_27),
.B1(n_36),
.B2(n_28),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_41),
.A2(n_26),
.B1(n_37),
.B2(n_34),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_26),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_95),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_47),
.A2(n_34),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_118),
.A2(n_35),
.B1(n_6),
.B2(n_9),
.Y(n_130)
);

NAND2x1p5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_51),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_125),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_135),
.Y(n_157)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_122),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_58),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_129),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_113),
.B(n_93),
.C(n_108),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_133),
.B(n_147),
.C(n_98),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_4),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_81),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_140),
.B1(n_100),
.B2(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_133)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_83),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_10),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_138),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_90),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_10),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_143),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_112),
.B(n_114),
.C(n_119),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_112),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_85),
.B1(n_117),
.B2(n_97),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_162),
.B1(n_169),
.B2(n_135),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_120),
.C(n_125),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_157),
.C(n_158),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_95),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_129),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_156),
.B1(n_164),
.B2(n_128),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_99),
.B1(n_100),
.B2(n_132),
.Y(n_156)
);

AO21x2_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_126),
.B(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_172),
.B1(n_169),
.B2(n_153),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_168),
.B(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_171),
.B(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_162),
.A2(n_141),
.B1(n_148),
.B2(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_128),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_133),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_131),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_136),
.C(n_143),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_169),
.B1(n_150),
.B2(n_164),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_198),
.B1(n_199),
.B2(n_193),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_181),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_197),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_169),
.B1(n_153),
.B2(n_158),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_179),
.B(n_177),
.C(n_183),
.D(n_152),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_203),
.B(n_204),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_174),
.B(n_163),
.C(n_131),
.D(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_205),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_175),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_155),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_209),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_149),
.B1(n_153),
.B2(n_130),
.Y(n_209)
);

XNOR2x2_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_191),
.Y(n_210)
);

AOI31xp67_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_203),
.A3(n_209),
.B(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_194),
.C(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_220),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_221),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_197),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_206),
.B(n_201),
.C(n_189),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_223),
.B(n_195),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_211),
.A2(n_195),
.B(n_122),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_215),
.B1(n_210),
.B2(n_212),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_215),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_213),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_229),
.B(n_230),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_225),
.A2(n_213),
.B(n_159),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_228),
.A2(n_227),
.B(n_224),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_231),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_159),
.C(n_138),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_232),
.B(n_134),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);


endmodule