module fake_jpeg_27105_n_67 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_24),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_12),
.B1(n_22),
.B2(n_21),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_26),
.B1(n_29),
.B2(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_9),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.C(n_1),
.Y(n_34)
);

OR2x4_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_4),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_31),
.C(n_30),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_43),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_48),
.B1(n_10),
.B2(n_11),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_7),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_14),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_16),
.C(n_20),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_11),
.C(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_35),
.B1(n_15),
.B2(n_13),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_54),
.B1(n_58),
.B2(n_57),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_53),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_57),
.Y(n_60)
);

XNOR2x1_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_51),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_56),
.C(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_59),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_55),
.C(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_52),
.Y(n_67)
);


endmodule