module fake_jpeg_3722_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_5),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_3),
.B(n_4),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_3),
.B(n_5),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx9p33_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_18),
.B1(n_17),
.B2(n_24),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_0),
.Y(n_17)
);

OAI21xp33_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_23),
.B(n_11),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_9),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_22),
.B(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_9),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_10),
.C(n_19),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_13),
.A2(n_15),
.B1(n_14),
.B2(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_7),
.B(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

AO21x1_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_34),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_29),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_10),
.C(n_23),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_30),
.B(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_17),
.C(n_10),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_35),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_31),
.B(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_41),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_44),
.C(n_43),
.Y(n_48)
);

AOI321xp33_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_40),
.A3(n_45),
.B1(n_47),
.B2(n_39),
.C(n_37),
.Y(n_49)
);


endmodule