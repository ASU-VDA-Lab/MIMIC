module fake_netlist_5_387_n_79 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_79);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_79;

wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_45;
wire n_46;
wire n_38;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_23;
wire n_29;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

INVxp67_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

OAI21x1_ASAP7_75t_L g29 ( 
.A1(n_15),
.A2(n_0),
.B(n_7),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_2),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_1),
.A2(n_19),
.B1(n_10),
.B2(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_38),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_9),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_12),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_21),
.B1(n_37),
.B2(n_36),
.Y(n_48)
);

OAI21x1_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_29),
.B(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

OAI22x1_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

O2A1O1Ixp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_42),
.B(n_39),
.C(n_47),
.Y(n_54)
);

OA21x2_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_39),
.B(n_31),
.Y(n_55)
);

OAI21x1_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_40),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_25),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_25),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_55),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_63),
.B(n_65),
.C(n_61),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_61),
.C(n_26),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_68),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_67),
.B(n_55),
.C(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OA21x2_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_56),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_76),
.Y(n_79)
);


endmodule