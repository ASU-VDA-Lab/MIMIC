module fake_jpeg_24654_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_38),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_37),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_2),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_26),
.B1(n_42),
.B2(n_29),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_20),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_28),
.B(n_18),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_29),
.C(n_32),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_18),
.B1(n_33),
.B2(n_19),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_27),
.B1(n_24),
.B2(n_31),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_2),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_35),
.B(n_40),
.C(n_43),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_72),
.B1(n_48),
.B2(n_61),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_25),
.B1(n_36),
.B2(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_77),
.B1(n_56),
.B2(n_47),
.Y(n_104)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_78),
.Y(n_105)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_17),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_15),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_80),
.B1(n_21),
.B2(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_32),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_92),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_90),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_21),
.B1(n_31),
.B2(n_27),
.Y(n_94)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_46),
.B(n_17),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_102),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_66),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_66),
.B1(n_91),
.B2(n_5),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_70),
.B(n_79),
.C(n_73),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_24),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_110),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_88),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_36),
.C(n_61),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_135),
.C(n_101),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_77),
.B(n_69),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_131),
.B(n_104),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_132),
.B1(n_102),
.B2(n_100),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_95),
.B1(n_94),
.B2(n_98),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_97),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_67),
.B(n_63),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_9),
.C(n_14),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_113),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_146),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_105),
.B1(n_106),
.B2(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_105),
.B(n_112),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_124),
.C(n_131),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_122),
.C(n_123),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_101),
.B1(n_9),
.B2(n_15),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_153),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_113),
.B(n_4),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_118),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_10),
.C(n_11),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_145),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_166),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_143),
.C(n_139),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_122),
.C(n_134),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_125),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_168),
.C(n_162),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_142),
.B(n_137),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_164),
.B(n_158),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_120),
.B1(n_144),
.B2(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_164),
.B1(n_161),
.B2(n_128),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_138),
.C(n_150),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_176),
.C(n_159),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_148),
.C(n_128),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_179),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_182),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_175),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_155),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_183),
.Y(n_189)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_167),
.C(n_173),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_119),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_188),
.Y(n_193)
);

FAx1_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_171),
.CI(n_170),
.CON(n_187),
.SN(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_11),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_178),
.B1(n_119),
.B2(n_113),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_188),
.C(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_4),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_187),
.C(n_189),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_193),
.B(n_6),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_5),
.C(n_7),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_199),
.B(n_7),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_7),
.Y(n_202)
);


endmodule