module fake_jpeg_18491_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

CKINVDCx6p67_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_40),
.Y(n_41)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_10),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_17),
.B1(n_30),
.B2(n_18),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_52),
.B(n_25),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_24),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_30),
.B1(n_17),
.B2(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_70),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_63),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_25),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_36),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_16),
.B(n_23),
.C(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_48),
.B1(n_39),
.B2(n_29),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_76),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_15),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_44),
.B1(n_15),
.B2(n_16),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_80),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_72),
.A2(n_43),
.B1(n_48),
.B2(n_23),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_48),
.B1(n_27),
.B2(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_90),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_68),
.B1(n_62),
.B2(n_64),
.Y(n_90)
);

NOR2xp67_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_13),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_26),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_104),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_90),
.B(n_86),
.C(n_89),
.D(n_87),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_29),
.B(n_69),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_91),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_61),
.B1(n_73),
.B2(n_69),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_57),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_11),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_11),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_69),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_82),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_131),
.B1(n_107),
.B2(n_105),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_128),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_73),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_122),
.C(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_126),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_97),
.C(n_79),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_82),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_57),
.C(n_20),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_134),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_127),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_140),
.B(n_124),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_101),
.C(n_98),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_118),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_111),
.B1(n_108),
.B2(n_109),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_118),
.B1(n_121),
.B2(n_130),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_145),
.B1(n_151),
.B2(n_152),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_139),
.C(n_133),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_125),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_143),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_102),
.B1(n_123),
.B2(n_125),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_109),
.B1(n_75),
.B2(n_59),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_138),
.B(n_142),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_159),
.B(n_0),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_157),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_158),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_75),
.C(n_9),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_0),
.B(n_1),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_162),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_7),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_158),
.C(n_152),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_168),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_6),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_9),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_167),
.B(n_171),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_173),
.B(n_12),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_14),
.Y(n_175)
);


endmodule