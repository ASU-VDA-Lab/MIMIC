module fake_jpeg_19987_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_19),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_69),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_28),
.B1(n_18),
.B2(n_33),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_61),
.B1(n_22),
.B2(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_31),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_25),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_63),
.B1(n_43),
.B2(n_18),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_34),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_25),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_72),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_74),
.A2(n_76),
.B1(n_89),
.B2(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_108),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_82),
.Y(n_125)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_109),
.Y(n_114)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_84),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_88),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_18),
.B(n_48),
.C(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_93),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_98),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_95),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_36),
.B(n_24),
.C(n_35),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_96),
.A2(n_80),
.B(n_108),
.C(n_110),
.Y(n_142)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_97),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_29),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_99),
.B(n_101),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_65),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_53),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_42),
.B1(n_39),
.B2(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_29),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_45),
.C(n_39),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_17),
.Y(n_146)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_45),
.Y(n_108)
);

AND2x4_ASAP7_75t_SL g109 ( 
.A(n_60),
.B(n_48),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_52),
.A2(n_33),
.B1(n_41),
.B2(n_36),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_27),
.B1(n_35),
.B2(n_57),
.Y(n_135)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_59),
.B1(n_50),
.B2(n_56),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_113),
.A2(n_135),
.B1(n_143),
.B2(n_97),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_55),
.B(n_58),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_115),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_58),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_16),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_56),
.A3(n_50),
.B1(n_51),
.B2(n_27),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_21),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_145),
.Y(n_165)
);

OR2x2_ASAP7_75t_SL g136 ( 
.A(n_96),
.B(n_17),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_11),
.C(n_15),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_87),
.A2(n_51),
.A3(n_57),
.B1(n_33),
.B2(n_47),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_16),
.B(n_9),
.C(n_10),
.D(n_14),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_78),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_76),
.A2(n_47),
.B1(n_51),
.B2(n_32),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_0),
.B(n_1),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_78),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_74),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_149),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_112),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_106),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_113),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_89),
.B1(n_83),
.B2(n_81),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_162),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_86),
.B1(n_111),
.B2(n_79),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_168),
.B(n_172),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_72),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_174),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_84),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_157),
.B(n_163),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_79),
.B1(n_82),
.B2(n_91),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_150),
.B1(n_165),
.B2(n_151),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_115),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_91),
.B1(n_32),
.B2(n_26),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_85),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_116),
.A2(n_32),
.B1(n_26),
.B2(n_90),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_166),
.B1(n_167),
.B2(n_125),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_32),
.B1(n_26),
.B2(n_90),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_26),
.B1(n_16),
.B2(n_3),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_8),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_11),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_121),
.B(n_1),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_173),
.B(n_177),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_7),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_119),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_114),
.B(n_118),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_7),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_128),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_180),
.A2(n_188),
.B(n_200),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_179),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_194),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_172),
.C(n_154),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_201),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

AOI32xp33_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_114),
.A3(n_120),
.B1(n_142),
.B2(n_118),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_143),
.C(n_120),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_168),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_135),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_138),
.Y(n_195)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_203),
.B1(n_176),
.B2(n_152),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_169),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_150),
.A2(n_132),
.B1(n_141),
.B2(n_140),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_132),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_205),
.B(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_127),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_153),
.A2(n_140),
.B1(n_127),
.B2(n_130),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_209),
.A2(n_160),
.B1(n_175),
.B2(n_165),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_227),
.B1(n_208),
.B2(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_212),
.B(n_213),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_204),
.B(n_197),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_220),
.B(n_184),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_224),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_151),
.B(n_157),
.Y(n_220)
);

AOI22x1_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_194),
.B1(n_193),
.B2(n_158),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_231),
.B1(n_232),
.B2(n_202),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_173),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_168),
.B1(n_166),
.B2(n_164),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_162),
.B1(n_127),
.B2(n_130),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

INVxp33_ASAP7_75t_SL g230 ( 
.A(n_208),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_192),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_207),
.B1(n_201),
.B2(n_181),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_261)
);

AO22x1_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_209),
.B1(n_188),
.B2(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_244),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_237),
.B1(n_238),
.B2(n_235),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_184),
.B(n_202),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_247),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_190),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_248),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_134),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_190),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_205),
.C(n_189),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_134),
.C(n_14),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_214),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_264),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_256),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_248),
.B(n_212),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_232),
.C(n_210),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_270),
.C(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_221),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_266),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_245),
.A2(n_216),
.B1(n_233),
.B2(n_206),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_265),
.B(n_250),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_227),
.B1(n_218),
.B2(n_185),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_206),
.B1(n_182),
.B2(n_192),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_159),
.B1(n_124),
.B2(n_134),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_2),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_260),
.B1(n_277),
.B2(n_281),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_241),
.B(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_235),
.CI(n_246),
.CON(n_276),
.SN(n_276)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_280),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_268),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_278),
.Y(n_286)
);

NAND4xp25_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_249),
.C(n_236),
.D(n_12),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_9),
.B(n_3),
.Y(n_282)
);

AO221x1_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_259),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_262),
.C(n_255),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_264),
.B1(n_261),
.B2(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_290),
.B(n_274),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_267),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_296),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_270),
.C(n_273),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_295),
.C(n_297),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_273),
.C(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_253),
.C(n_255),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_292),
.B(n_276),
.Y(n_301)
);

NOR2x1_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_286),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_290),
.B1(n_279),
.B2(n_254),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_3),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_276),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_4),
.B(n_5),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_307),
.C(n_302),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_300),
.C(n_303),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_R g311 ( 
.A(n_310),
.B(n_308),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_5),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_5),
.Y(n_313)
);


endmodule