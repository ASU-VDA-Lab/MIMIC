module real_aes_11409_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_0), .A2(n_194), .B1(n_349), .B2(n_352), .Y(n_348) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_0), .A2(n_5), .B1(n_417), .B2(n_435), .Y(n_434) );
AOI21xp33_ASAP7_75t_L g575 ( .A1(n_1), .A2(n_522), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g602 ( .A(n_1), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g804 ( .A1(n_2), .A2(n_63), .B1(n_441), .B2(n_797), .Y(n_804) );
INVxp67_ASAP7_75t_SL g821 ( .A(n_2), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g1143 ( .A1(n_3), .A2(n_4), .B1(n_1138), .B2(n_1144), .Y(n_1143) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_5), .A2(n_161), .B1(n_342), .B2(n_344), .C(n_346), .Y(n_341) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_6), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_6), .B(n_185), .Y(n_285) );
AND2x2_ASAP7_75t_L g404 ( .A(n_6), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g447 ( .A(n_6), .Y(n_447) );
INVxp67_ASAP7_75t_L g639 ( .A(n_7), .Y(n_639) );
OAI222xp33_ASAP7_75t_L g657 ( .A1(n_7), .A2(n_38), .B1(n_237), .B2(n_658), .C1(n_659), .C2(n_661), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g1148 ( .A1(n_8), .A2(n_214), .B1(n_1122), .B2(n_1130), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_9), .A2(n_39), .B1(n_1393), .B2(n_1395), .Y(n_1392) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_9), .A2(n_39), .B1(n_507), .B2(n_702), .Y(n_1398) );
AOI221xp5_ASAP7_75t_L g1079 ( .A1(n_10), .A2(n_164), .B1(n_322), .B2(n_1080), .C(n_1081), .Y(n_1079) );
INVx1_ASAP7_75t_L g1098 ( .A(n_10), .Y(n_1098) );
INVx1_ASAP7_75t_L g1339 ( .A(n_11), .Y(n_1339) );
AO22x2_ASAP7_75t_L g451 ( .A1(n_12), .A2(n_452), .B1(n_540), .B2(n_541), .Y(n_451) );
CKINVDCx14_ASAP7_75t_R g540 ( .A(n_12), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_13), .A2(n_71), .B1(n_702), .B2(n_703), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_13), .A2(n_24), .B1(n_729), .B2(n_743), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_14), .A2(n_33), .B1(n_317), .B2(n_322), .Y(n_316) );
INVxp33_ASAP7_75t_SL g415 ( .A(n_14), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_15), .A2(n_224), .B1(n_673), .B2(n_702), .Y(n_1088) );
INVx1_ASAP7_75t_L g1106 ( .A(n_15), .Y(n_1106) );
AOI221xp5_ASAP7_75t_L g838 ( .A1(n_16), .A2(n_236), .B1(n_680), .B2(n_681), .C(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g862 ( .A(n_16), .Y(n_862) );
OAI221xp5_ASAP7_75t_L g548 ( .A1(n_17), .A2(n_549), .B1(n_550), .B2(n_556), .C(n_561), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_17), .A2(n_162), .B1(n_584), .B2(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_18), .A2(n_135), .B1(n_584), .B2(n_751), .C(n_752), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_18), .A2(n_207), .B1(n_770), .B2(n_771), .Y(n_769) );
INVx2_ASAP7_75t_L g294 ( .A(n_19), .Y(n_294) );
OR2x2_ASAP7_75t_L g328 ( .A(n_19), .B(n_292), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g915 ( .A1(n_20), .A2(n_175), .B1(n_800), .B2(n_916), .C(n_918), .Y(n_915) );
INVx1_ASAP7_75t_L g926 ( .A(n_20), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_21), .A2(n_54), .B1(n_503), .B2(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g741 ( .A(n_21), .Y(n_741) );
OAI221xp5_ASAP7_75t_L g1032 ( .A1(n_22), .A2(n_95), .B1(n_867), .B2(n_1033), .C(n_1035), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_22), .A2(n_95), .B1(n_653), .B2(n_844), .Y(n_1060) );
INVx1_ASAP7_75t_L g642 ( .A(n_23), .Y(n_642) );
OAI222xp33_ASAP7_75t_L g764 ( .A1(n_24), .A2(n_135), .B1(n_139), .B2(n_286), .C1(n_765), .C2(n_768), .Y(n_764) );
OR2x2_ASAP7_75t_L g284 ( .A(n_25), .B(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g288 ( .A(n_25), .Y(n_288) );
BUFx2_ASAP7_75t_L g377 ( .A(n_25), .Y(n_377) );
INVx1_ASAP7_75t_L g403 ( .A(n_25), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g1176 ( .A(n_26), .Y(n_1176) );
INVx1_ASAP7_75t_L g455 ( .A(n_27), .Y(n_455) );
AOI21xp33_ASAP7_75t_L g528 ( .A1(n_27), .A2(n_319), .B(n_346), .Y(n_528) );
INVx1_ASAP7_75t_L g900 ( .A(n_28), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_29), .Y(n_480) );
INVx1_ASAP7_75t_L g1346 ( .A(n_30), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_30), .A2(n_82), .B1(n_584), .B2(n_597), .Y(n_1389) );
INVx1_ASAP7_75t_L g956 ( .A(n_31), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_32), .A2(n_123), .B1(n_319), .B2(n_323), .Y(n_574) );
INVx1_ASAP7_75t_L g604 ( .A(n_32), .Y(n_604) );
INVxp33_ASAP7_75t_SL g396 ( .A(n_33), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_34), .A2(n_170), .B1(n_441), .B2(n_797), .Y(n_796) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_34), .A2(n_229), .B1(n_823), .B2(n_824), .C(n_826), .Y(n_822) );
INVx1_ASAP7_75t_L g626 ( .A(n_35), .Y(n_626) );
INVx1_ASAP7_75t_L g1352 ( .A(n_36), .Y(n_1352) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_36), .A2(n_132), .B1(n_1367), .B2(n_1369), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_37), .A2(n_45), .B1(n_592), .B2(n_747), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_37), .A2(n_45), .B1(n_354), .B2(n_847), .Y(n_1399) );
INVxp67_ASAP7_75t_L g637 ( .A(n_38), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g529 ( .A1(n_40), .A2(n_202), .B1(n_530), .B2(n_531), .C(n_533), .Y(n_529) );
INVx1_ASAP7_75t_L g538 ( .A(n_40), .Y(n_538) );
INVx1_ASAP7_75t_L g907 ( .A(n_41), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_42), .A2(n_44), .B1(n_916), .B2(n_1422), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1463 ( .A1(n_42), .A2(n_56), .B1(n_770), .B2(n_771), .Y(n_1463) );
INVx1_ASAP7_75t_L g720 ( .A(n_43), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g755 ( .A1(n_43), .A2(n_72), .B1(n_756), .B2(n_760), .C(n_761), .Y(n_755) );
INVxp67_ASAP7_75t_SL g1460 ( .A(n_44), .Y(n_1460) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_46), .A2(n_80), .B1(n_799), .B2(n_801), .Y(n_803) );
INVxp33_ASAP7_75t_SL g832 ( .A(n_46), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_47), .A2(n_162), .B1(n_366), .B2(n_372), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_47), .A2(n_243), .B1(n_587), .B2(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g1434 ( .A(n_48), .Y(n_1434) );
CKINVDCx5p33_ASAP7_75t_R g1083 ( .A(n_49), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_50), .A2(n_180), .B1(n_958), .B2(n_959), .Y(n_957) );
INVxp67_ASAP7_75t_SL g1003 ( .A(n_50), .Y(n_1003) );
INVx1_ASAP7_75t_L g1053 ( .A(n_51), .Y(n_1053) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_52), .Y(n_1009) );
AOI22xp5_ASAP7_75t_L g1149 ( .A1(n_53), .A2(n_73), .B1(n_1138), .B2(n_1144), .Y(n_1149) );
INVx1_ASAP7_75t_L g740 ( .A(n_54), .Y(n_740) );
AOI22xp5_ASAP7_75t_SL g1133 ( .A1(n_55), .A2(n_67), .B1(n_1134), .B2(n_1138), .Y(n_1133) );
AOI221xp5_ASAP7_75t_L g1424 ( .A1(n_56), .A2(n_176), .B1(n_752), .B2(n_1393), .C(n_1395), .Y(n_1424) );
INVxp33_ASAP7_75t_SL g1040 ( .A(n_57), .Y(n_1040) );
AOI221xp5_ASAP7_75t_L g1065 ( .A1(n_57), .A2(n_86), .B1(n_847), .B2(n_930), .C(n_932), .Y(n_1065) );
AOI221xp5_ASAP7_75t_L g902 ( .A1(n_58), .A2(n_113), .B1(n_747), .B2(n_903), .C(n_904), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_58), .A2(n_78), .B1(n_934), .B2(n_935), .Y(n_933) );
CKINVDCx16_ASAP7_75t_R g1174 ( .A(n_59), .Y(n_1174) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_60), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_60), .A2(n_131), .B1(n_849), .B2(n_1403), .Y(n_1402) );
INVxp33_ASAP7_75t_SL g364 ( .A(n_61), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_61), .A2(n_100), .B1(n_431), .B2(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_62), .A2(n_218), .B1(n_322), .B2(n_565), .Y(n_840) );
INVx1_ASAP7_75t_L g863 ( .A(n_62), .Y(n_863) );
INVxp33_ASAP7_75t_L g831 ( .A(n_63), .Y(n_831) );
INVx1_ASAP7_75t_L g906 ( .A(n_64), .Y(n_906) );
AOI221xp5_ASAP7_75t_L g928 ( .A1(n_64), .A2(n_113), .B1(n_929), .B2(n_930), .C(n_932), .Y(n_928) );
INVxp33_ASAP7_75t_L g1026 ( .A(n_65), .Y(n_1026) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_65), .A2(n_247), .B1(n_322), .B2(n_929), .C(n_1062), .Y(n_1061) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_66), .A2(n_129), .B1(n_678), .B2(n_680), .C(n_681), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_66), .A2(n_143), .B1(n_685), .B2(n_686), .C(n_688), .Y(n_684) );
INVxp33_ASAP7_75t_SL g1334 ( .A(n_68), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g1387 ( .A1(n_68), .A2(n_160), .B1(n_747), .B2(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g292 ( .A(n_69), .Y(n_292) );
INVx1_ASAP7_75t_L g315 ( .A(n_69), .Y(n_315) );
INVxp33_ASAP7_75t_L g370 ( .A(n_70), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_70), .A2(n_190), .B1(n_417), .B2(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g754 ( .A(n_71), .Y(n_754) );
INVx1_ASAP7_75t_L g716 ( .A(n_72), .Y(n_716) );
INVx1_ASAP7_75t_L g919 ( .A(n_74), .Y(n_919) );
OAI221xp5_ASAP7_75t_L g923 ( .A1(n_74), .A2(n_175), .B1(n_659), .B2(n_924), .C(n_925), .Y(n_923) );
AO221x2_ASAP7_75t_L g1150 ( .A1(n_75), .A2(n_234), .B1(n_1138), .B2(n_1144), .C(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g557 ( .A(n_76), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_76), .A2(n_138), .B1(n_583), .B2(n_584), .Y(n_582) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_77), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_77), .A2(n_201), .B1(n_811), .B2(n_812), .Y(n_810) );
INVxp67_ASAP7_75t_SL g905 ( .A(n_78), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_79), .A2(n_114), .B1(n_322), .B2(n_967), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_79), .A2(n_114), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_80), .Y(n_809) );
INVx1_ASAP7_75t_L g913 ( .A(n_81), .Y(n_913) );
AOI221xp5_ASAP7_75t_L g937 ( .A1(n_81), .A2(n_126), .B1(n_502), .B2(n_938), .C(n_939), .Y(n_937) );
INVxp33_ASAP7_75t_SL g1329 ( .A(n_82), .Y(n_1329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_83), .A2(n_227), .B1(n_331), .B2(n_336), .Y(n_330) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_83), .Y(n_384) );
INVx1_ASAP7_75t_L g1436 ( .A(n_84), .Y(n_1436) );
AOI221xp5_ASAP7_75t_L g1442 ( .A1(n_84), .A2(n_240), .B1(n_344), .B2(n_1443), .C(n_1444), .Y(n_1442) );
XNOR2xp5_ASAP7_75t_L g611 ( .A(n_85), .B(n_612), .Y(n_611) );
INVxp67_ASAP7_75t_SL g1043 ( .A(n_86), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_87), .A2(n_545), .B1(n_607), .B2(n_608), .Y(n_544) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_87), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_88), .Y(n_852) );
INVxp67_ASAP7_75t_L g622 ( .A(n_89), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_89), .A2(n_148), .B1(n_507), .B2(n_665), .C(n_666), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_90), .A2(n_221), .B1(n_1122), .B2(n_1188), .Y(n_1187) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_91), .A2(n_142), .B1(n_680), .B2(n_700), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g737 ( .A1(n_91), .A2(n_473), .B(n_489), .Y(n_737) );
OAI21xp33_ASAP7_75t_L g896 ( .A1(n_92), .A2(n_897), .B(n_921), .Y(n_896) );
INVx1_ASAP7_75t_L g944 ( .A(n_92), .Y(n_944) );
CKINVDCx20_ASAP7_75t_R g1197 ( .A(n_93), .Y(n_1197) );
INVx1_ASAP7_75t_L g920 ( .A(n_94), .Y(n_920) );
AOI221xp5_ASAP7_75t_L g846 ( .A1(n_96), .A2(n_204), .B1(n_560), .B2(n_839), .C(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g879 ( .A(n_96), .Y(n_879) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_97), .A2(n_220), .B1(n_718), .B2(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g989 ( .A(n_97), .Y(n_989) );
INVxp33_ASAP7_75t_SL g1379 ( .A(n_98), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1401 ( .A1(n_98), .A2(n_211), .B1(n_507), .B2(n_702), .Y(n_1401) );
INVx1_ASAP7_75t_L g255 ( .A(n_99), .Y(n_255) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_100), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_101), .Y(n_1090) );
CKINVDCx5p33_ASAP7_75t_R g854 ( .A(n_102), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_103), .Y(n_477) );
OA22x2_ASAP7_75t_L g833 ( .A1(n_104), .A2(n_834), .B1(n_890), .B2(n_891), .Y(n_833) );
INVx1_ASAP7_75t_L g891 ( .A(n_104), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_105), .Y(n_300) );
INVx1_ASAP7_75t_L g964 ( .A(n_106), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_106), .A2(n_992), .B1(n_994), .B2(n_1000), .C(n_1004), .Y(n_991) );
XOR2x2_ASAP7_75t_L g946 ( .A(n_107), .B(n_947), .Y(n_946) );
OAI221xp5_ASAP7_75t_SL g910 ( .A1(n_108), .A2(n_217), .B1(n_739), .B2(n_911), .C(n_912), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_108), .A2(n_217), .B1(n_343), .B2(n_354), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_109), .A2(n_203), .B1(n_1122), .B2(n_1130), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_110), .A2(n_177), .B1(n_981), .B2(n_982), .C(n_984), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_110), .A2(n_155), .B1(n_770), .B2(n_771), .Y(n_1014) );
INVx1_ASAP7_75t_L g1054 ( .A(n_111), .Y(n_1054) );
OAI222xp33_ASAP7_75t_L g614 ( .A1(n_112), .A2(n_147), .B1(n_241), .B2(n_283), .C1(n_615), .C2(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g651 ( .A(n_112), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_115), .A2(n_116), .B1(n_1134), .B2(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g977 ( .A(n_117), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_117), .A2(n_177), .B1(n_765), .B2(n_768), .Y(n_1015) );
INVx1_ASAP7_75t_L g1440 ( .A(n_118), .Y(n_1440) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_119), .Y(n_484) );
CKINVDCx14_ASAP7_75t_R g1153 ( .A(n_120), .Y(n_1153) );
AOI22xp5_ASAP7_75t_L g1142 ( .A1(n_121), .A2(n_141), .B1(n_1122), .B2(n_1130), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_122), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_123), .A2(n_232), .B1(n_497), .B2(n_606), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_124), .Y(n_569) );
XNOR2xp5_ASAP7_75t_L g690 ( .A(n_125), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g914 ( .A(n_126), .Y(n_914) );
INVx1_ASAP7_75t_L g1048 ( .A(n_127), .Y(n_1048) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_128), .A2(n_244), .B1(n_665), .B2(n_932), .C(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1105 ( .A(n_128), .Y(n_1105) );
OAI332xp33_ASAP7_75t_L g620 ( .A1(n_129), .A2(n_472), .A3(n_494), .B1(n_621), .B2(n_627), .B3(n_632), .C1(n_638), .C2(n_645), .Y(n_620) );
INVx1_ASAP7_75t_L g459 ( .A(n_130), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_130), .A2(n_179), .B1(n_323), .B2(n_527), .Y(n_526) );
INVxp33_ASAP7_75t_L g1373 ( .A(n_131), .Y(n_1373) );
INVx1_ASAP7_75t_L g1348 ( .A(n_132), .Y(n_1348) );
CKINVDCx5p33_ASAP7_75t_R g1076 ( .A(n_133), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1425 ( .A1(n_134), .A2(n_193), .B1(n_756), .B2(n_760), .Y(n_1425) );
OAI221xp5_ASAP7_75t_L g1452 ( .A1(n_134), .A2(n_193), .B1(n_1453), .B2(n_1455), .C(n_1456), .Y(n_1452) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_136), .Y(n_806) );
XNOR2xp5_ASAP7_75t_L g1071 ( .A(n_137), .B(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g553 ( .A(n_138), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_139), .A2(n_207), .B1(n_747), .B2(n_748), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_140), .A2(n_152), .B1(n_706), .B2(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g730 ( .A(n_140), .Y(n_730) );
XOR2x2_ASAP7_75t_L g778 ( .A(n_141), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g736 ( .A(n_142), .Y(n_736) );
INVx1_ASAP7_75t_L g676 ( .A(n_143), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_144), .A2(n_172), .B1(n_492), .B2(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g513 ( .A(n_144), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_145), .A2(n_197), .B1(n_283), .B2(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_145), .A2(n_172), .B1(n_319), .B2(n_323), .Y(n_518) );
AOI21xp33_ASAP7_75t_L g559 ( .A1(n_146), .A2(n_343), .B(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_146), .A2(n_231), .B1(n_587), .B2(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g671 ( .A(n_147), .Y(n_671) );
INVx1_ASAP7_75t_L g628 ( .A(n_148), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_149), .Y(n_478) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_150), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_150), .B(n_255), .Y(n_1129) );
AND3x2_ASAP7_75t_L g1137 ( .A(n_150), .B(n_255), .C(n_1126), .Y(n_1137) );
OA332x1_ASAP7_75t_L g453 ( .A1(n_151), .A2(n_454), .A3(n_463), .B1(n_472), .B2(n_475), .B3(n_479), .C1(n_486), .C2(n_487), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_151), .A2(n_520), .B(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g732 ( .A(n_152), .Y(n_732) );
INVxp33_ASAP7_75t_L g1038 ( .A(n_153), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_153), .A2(n_181), .B1(n_934), .B2(n_935), .Y(n_1066) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_154), .A2(n_222), .B1(n_304), .B2(n_309), .C(n_312), .Y(n_303) );
INVxp33_ASAP7_75t_SL g406 ( .A(n_154), .Y(n_406) );
INVx1_ASAP7_75t_L g979 ( .A(n_155), .Y(n_979) );
INVx1_ASAP7_75t_L g1068 ( .A(n_156), .Y(n_1068) );
OAI22xp33_ASAP7_75t_SL g1077 ( .A1(n_157), .A2(n_171), .B1(n_653), .B2(n_1078), .Y(n_1077) );
OAI221xp5_ASAP7_75t_L g1099 ( .A1(n_157), .A2(n_171), .B1(n_867), .B2(n_1033), .C(n_1035), .Y(n_1099) );
INVx2_ASAP7_75t_L g268 ( .A(n_158), .Y(n_268) );
AOI22xp5_ASAP7_75t_SL g1192 ( .A1(n_159), .A2(n_225), .B1(n_1122), .B2(n_1130), .Y(n_1192) );
INVxp33_ASAP7_75t_SL g1343 ( .A(n_160), .Y(n_1343) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_161), .A2(n_194), .B1(n_428), .B2(n_431), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_163), .A2(n_226), .B1(n_680), .B2(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g875 ( .A(n_163), .Y(n_875) );
INVx1_ASAP7_75t_L g1096 ( .A(n_164), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_165), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_166), .Y(n_792) );
INVx1_ASAP7_75t_L g899 ( .A(n_167), .Y(n_899) );
INVxp33_ASAP7_75t_SL g793 ( .A(n_168), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g813 ( .A1(n_168), .A2(n_212), .B1(n_814), .B2(n_816), .C(n_817), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_169), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_170), .A2(n_191), .B1(n_354), .B2(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g1126 ( .A(n_173), .Y(n_1126) );
AOI22xp5_ASAP7_75t_SL g1193 ( .A1(n_174), .A2(n_200), .B1(n_1134), .B2(n_1138), .Y(n_1193) );
INVxp67_ASAP7_75t_SL g1462 ( .A(n_176), .Y(n_1462) );
INVx1_ASAP7_75t_L g1433 ( .A(n_178), .Y(n_1433) );
INVx1_ASAP7_75t_L g464 ( .A(n_179), .Y(n_464) );
INVxp67_ASAP7_75t_SL g1001 ( .A(n_180), .Y(n_1001) );
INVxp67_ASAP7_75t_SL g1044 ( .A(n_181), .Y(n_1044) );
AO221x2_ASAP7_75t_L g1194 ( .A1(n_182), .A2(n_248), .B1(n_1190), .B2(n_1195), .C(n_1196), .Y(n_1194) );
OAI211xp5_ASAP7_75t_L g1419 ( .A1(n_183), .A2(n_973), .B(n_1420), .C(n_1426), .Y(n_1419) );
AOI221xp5_ASAP7_75t_L g1446 ( .A1(n_183), .A2(n_189), .B1(n_824), .B2(n_1447), .C(n_1448), .Y(n_1446) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_184), .Y(n_278) );
INVx1_ASAP7_75t_L g270 ( .A(n_185), .Y(n_270) );
INVx2_ASAP7_75t_L g405 ( .A(n_185), .Y(n_405) );
INVx1_ASAP7_75t_L g1427 ( .A(n_186), .Y(n_1427) );
OR2x2_ASAP7_75t_L g546 ( .A(n_187), .B(n_282), .Y(n_546) );
CKINVDCx14_ASAP7_75t_R g1199 ( .A(n_188), .Y(n_1199) );
OAI221xp5_ASAP7_75t_L g1429 ( .A1(n_189), .A2(n_992), .B1(n_1004), .B2(n_1430), .C(n_1435), .Y(n_1429) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_190), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_191), .A2(n_229), .B1(n_799), .B2(n_801), .Y(n_798) );
INVx1_ASAP7_75t_L g1051 ( .A(n_192), .Y(n_1051) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_195), .Y(n_1085) );
INVx1_ASAP7_75t_L g1030 ( .A(n_196), .Y(n_1030) );
INVx1_ASAP7_75t_L g534 ( .A(n_197), .Y(n_534) );
INVx1_ASAP7_75t_L g954 ( .A(n_198), .Y(n_954) );
CKINVDCx16_ASAP7_75t_R g1171 ( .A(n_199), .Y(n_1171) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_201), .Y(n_786) );
INVx1_ASAP7_75t_L g539 ( .A(n_202), .Y(n_539) );
INVx1_ASAP7_75t_L g1021 ( .A(n_203), .Y(n_1021) );
INVx1_ASAP7_75t_L g876 ( .A(n_204), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_205), .Y(n_841) );
INVx1_ASAP7_75t_L g790 ( .A(n_206), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_208), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_209), .A2(n_216), .B1(n_843), .B2(n_844), .Y(n_842) );
OAI221xp5_ASAP7_75t_L g864 ( .A1(n_209), .A2(n_216), .B1(n_865), .B2(n_867), .C(n_868), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_210), .A2(n_1414), .B1(n_1415), .B2(n_1416), .Y(n_1413) );
CKINVDCx5p33_ASAP7_75t_R g1414 ( .A(n_210), .Y(n_1414) );
INVxp67_ASAP7_75t_SL g1362 ( .A(n_211), .Y(n_1362) );
INVxp33_ASAP7_75t_SL g788 ( .A(n_212), .Y(n_788) );
INVx1_ASAP7_75t_L g1127 ( .A(n_213), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_213), .B(n_1125), .Y(n_1132) );
XOR2x2_ASAP7_75t_L g1325 ( .A(n_214), .B(n_1326), .Y(n_1325) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_214), .A2(n_1410), .B1(n_1412), .B2(n_1464), .Y(n_1409) );
INVx1_ASAP7_75t_L g654 ( .A(n_215), .Y(n_654) );
INVx1_ASAP7_75t_L g859 ( .A(n_218), .Y(n_859) );
INVx1_ASAP7_75t_L g631 ( .A(n_219), .Y(n_631) );
INVx1_ASAP7_75t_L g986 ( .A(n_220), .Y(n_986) );
INVxp33_ASAP7_75t_L g410 ( .A(n_222), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g1082 ( .A(n_223), .Y(n_1082) );
INVx1_ASAP7_75t_L g1102 ( .A(n_224), .Y(n_1102) );
INVx1_ASAP7_75t_L g881 ( .A(n_226), .Y(n_881) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_227), .Y(n_389) );
INVx2_ASAP7_75t_L g267 ( .A(n_228), .Y(n_267) );
INVx1_ASAP7_75t_L g965 ( .A(n_230), .Y(n_965) );
OAI211xp5_ASAP7_75t_SL g972 ( .A1(n_230), .A2(n_973), .B(n_974), .C(n_985), .Y(n_972) );
INVx1_ASAP7_75t_L g555 ( .A(n_231), .Y(n_555) );
INVx1_ASAP7_75t_L g572 ( .A(n_232), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_233), .Y(n_467) );
INVx1_ASAP7_75t_L g1428 ( .A(n_235), .Y(n_1428) );
INVx1_ASAP7_75t_L g860 ( .A(n_236), .Y(n_860) );
INVxp67_ASAP7_75t_L g633 ( .A(n_237), .Y(n_633) );
INVx1_ASAP7_75t_L g1028 ( .A(n_238), .Y(n_1028) );
INVx1_ASAP7_75t_L g1092 ( .A(n_239), .Y(n_1092) );
AOI21xp33_ASAP7_75t_L g1437 ( .A1(n_240), .A2(n_473), .B(n_1393), .Y(n_1437) );
INVx1_ASAP7_75t_L g655 ( .A(n_241), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g1168 ( .A(n_242), .Y(n_1168) );
OAI211xp5_ASAP7_75t_SL g562 ( .A1(n_243), .A2(n_563), .B(n_566), .C(n_571), .Y(n_562) );
INVx1_ASAP7_75t_L g1103 ( .A(n_244), .Y(n_1103) );
BUFx3_ASAP7_75t_L g297 ( .A(n_245), .Y(n_297) );
INVx1_ASAP7_75t_L g325 ( .A(n_245), .Y(n_325) );
BUFx3_ASAP7_75t_L g299 ( .A(n_246), .Y(n_299) );
INVx1_ASAP7_75t_L g321 ( .A(n_246), .Y(n_321) );
INVxp33_ASAP7_75t_L g1031 ( .A(n_247), .Y(n_1031) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_271), .B(n_1114), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_258), .Y(n_252) );
AND2x4_ASAP7_75t_L g1408 ( .A(n_253), .B(n_259), .Y(n_1408) );
NOR2xp33_ASAP7_75t_SL g253 ( .A(n_254), .B(n_256), .Y(n_253) );
INVx1_ASAP7_75t_SL g1411 ( .A(n_254), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_254), .B(n_256), .Y(n_1467) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_256), .B(n_1411), .Y(n_1410) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_264), .Y(n_259) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g1384 ( .A(n_261), .B(n_288), .Y(n_1384) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g426 ( .A(n_262), .B(n_270), .Y(n_426) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g473 ( .A(n_263), .B(n_474), .Y(n_473) );
INVx8_ASAP7_75t_L g1380 ( .A(n_264), .Y(n_1380) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
OR2x2_ASAP7_75t_L g283 ( .A(n_265), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_SL g466 ( .A(n_265), .Y(n_466) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_265), .Y(n_476) );
INVx1_ASAP7_75t_L g641 ( .A(n_265), .Y(n_641) );
BUFx2_ASAP7_75t_L g874 ( .A(n_265), .Y(n_874) );
OAI22xp33_ASAP7_75t_L g904 ( .A1(n_265), .A2(n_469), .B1(n_905), .B2(n_906), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g918 ( .A1(n_265), .A2(n_469), .B1(n_919), .B2(n_920), .Y(n_918) );
INVx2_ASAP7_75t_SL g998 ( .A(n_265), .Y(n_998) );
OR2x6_ASAP7_75t_L g1382 ( .A(n_265), .B(n_1372), .Y(n_1382) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g388 ( .A(n_267), .Y(n_388) );
INVx1_ASAP7_75t_L g393 ( .A(n_267), .Y(n_393) );
AND2x4_ASAP7_75t_L g401 ( .A(n_267), .B(n_394), .Y(n_401) );
AND2x2_ASAP7_75t_L g414 ( .A(n_267), .B(n_268), .Y(n_414) );
INVx2_ASAP7_75t_L g419 ( .A(n_267), .Y(n_419) );
INVx1_ASAP7_75t_L g382 ( .A(n_268), .Y(n_382) );
INVx2_ASAP7_75t_L g394 ( .A(n_268), .Y(n_394) );
INVx1_ASAP7_75t_L g421 ( .A(n_268), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_268), .B(n_419), .Y(n_458) );
INVx1_ASAP7_75t_L g471 ( .A(n_268), .Y(n_471) );
AND2x4_ASAP7_75t_L g1368 ( .A(n_269), .B(n_382), .Y(n_1368) );
INVx2_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_270), .B(n_387), .Y(n_1369) );
XNOR2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_774), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_609), .B2(n_610), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
XOR2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_448), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
XNOR2x1_ASAP7_75t_SL g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_378), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_300), .B(n_301), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_281), .A2(n_806), .B(n_807), .Y(n_805) );
INVx5_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_SL g855 ( .A(n_282), .Y(n_855) );
INVx2_ASAP7_75t_L g1069 ( .A(n_282), .Y(n_1069) );
AND2x4_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx2_ASAP7_75t_L g908 ( .A(n_283), .Y(n_908) );
INVx3_ASAP7_75t_L g383 ( .A(n_284), .Y(n_383) );
INVx1_ASAP7_75t_L g744 ( .A(n_285), .Y(n_744) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x6_ASAP7_75t_L g1010 ( .A(n_287), .B(n_1011), .Y(n_1010) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AND2x4_ASAP7_75t_L g709 ( .A(n_288), .B(n_314), .Y(n_709) );
AND2x4_ASAP7_75t_L g962 ( .A(n_288), .B(n_314), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_289), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g650 ( .A(n_289), .Y(n_650) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_295), .Y(n_289) );
AND2x4_ASAP7_75t_L g332 ( .A(n_290), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g337 ( .A(n_290), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g362 ( .A(n_290), .Y(n_362) );
BUFx2_ASAP7_75t_L g510 ( .A(n_290), .Y(n_510) );
AND2x2_ASAP7_75t_L g532 ( .A(n_290), .B(n_338), .Y(n_532) );
AND2x4_ASAP7_75t_L g568 ( .A(n_290), .B(n_333), .Y(n_568) );
AND2x4_ASAP7_75t_L g570 ( .A(n_290), .B(n_338), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g715 ( .A(n_290), .B(n_444), .Y(n_715) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g314 ( .A(n_293), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g347 ( .A(n_294), .B(n_315), .Y(n_347) );
INVx1_ASAP7_75t_L g1332 ( .A(n_294), .Y(n_1332) );
INVx1_ASAP7_75t_L g1337 ( .A(n_294), .Y(n_1337) );
HB1xp67_ASAP7_75t_L g1342 ( .A(n_294), .Y(n_1342) );
INVx6_ASAP7_75t_L g311 ( .A(n_295), .Y(n_311) );
INVx2_ASAP7_75t_L g521 ( .A(n_295), .Y(n_521) );
AND2x4_ASAP7_75t_L g1340 ( .A(n_295), .B(n_1341), .Y(n_1340) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g339 ( .A(n_296), .Y(n_339) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g308 ( .A(n_297), .B(n_299), .Y(n_308) );
AND2x4_ASAP7_75t_L g320 ( .A(n_297), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g324 ( .A(n_299), .B(n_325), .Y(n_324) );
AOI31xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_340), .A3(n_363), .B(n_374), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_316), .B1(n_326), .B2(n_329), .C(n_330), .Y(n_302) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g345 ( .A(n_306), .Y(n_345) );
AND2x4_ASAP7_75t_L g360 ( .A(n_306), .B(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g1347 ( .A(n_306), .Y(n_1347) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g704 ( .A(n_307), .Y(n_704) );
INVx1_ASAP7_75t_L g723 ( .A(n_307), .Y(n_723) );
BUFx6f_ASAP7_75t_L g938 ( .A(n_307), .Y(n_938) );
AND2x4_ASAP7_75t_L g1355 ( .A(n_307), .B(n_1356), .Y(n_1355) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_308), .Y(n_358) );
INVx4_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g702 ( .A(n_310), .Y(n_702) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
INVx2_ASAP7_75t_L g502 ( .A(n_311), .Y(n_502) );
INVx1_ASAP7_75t_L g527 ( .A(n_311), .Y(n_527) );
INVx1_ASAP7_75t_L g680 ( .A(n_311), .Y(n_680) );
INVx2_ASAP7_75t_L g1333 ( .A(n_311), .Y(n_1333) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_SL g522 ( .A(n_314), .Y(n_522) );
INVx1_ASAP7_75t_L g681 ( .A(n_314), .Y(n_681) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_314), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g939 ( .A(n_314), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_314), .A2(n_516), .B1(n_766), .B2(n_1028), .C(n_1030), .Y(n_1062) );
OAI221xp5_ASAP7_75t_L g1081 ( .A1(n_314), .A2(n_516), .B1(n_766), .B2(n_1082), .C(n_1083), .Y(n_1081) );
INVx1_ASAP7_75t_L g1358 ( .A(n_315), .Y(n_1358) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g326 ( .A(n_319), .B(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g967 ( .A(n_319), .Y(n_967) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_320), .Y(n_343) );
INVx2_ASAP7_75t_SL g506 ( .A(n_320), .Y(n_506) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_320), .Y(n_565) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_320), .Y(n_665) );
BUFx3_ASAP7_75t_L g706 ( .A(n_320), .Y(n_706) );
BUFx2_ASAP7_75t_L g847 ( .A(n_320), .Y(n_847) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_320), .Y(n_1080) );
AND2x6_ASAP7_75t_L g1335 ( .A(n_320), .B(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g554 ( .A(n_323), .Y(n_554) );
BUFx3_ASAP7_75t_L g816 ( .A(n_323), .Y(n_816) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
INVx2_ASAP7_75t_L g373 ( .A(n_324), .Y(n_373) );
INVx1_ASAP7_75t_L g708 ( .A(n_324), .Y(n_708) );
INVx1_ASAP7_75t_L g960 ( .A(n_324), .Y(n_960) );
INVx1_ASAP7_75t_L g368 ( .A(n_325), .Y(n_368) );
AOI211xp5_ASAP7_75t_L g808 ( .A1(n_326), .A2(n_809), .B(n_810), .C(n_813), .Y(n_808) );
AOI211xp5_ASAP7_75t_SL g1059 ( .A1(n_326), .A2(n_1048), .B(n_1060), .C(n_1061), .Y(n_1059) );
AOI211xp5_ASAP7_75t_SL g1075 ( .A1(n_326), .A2(n_1076), .B(n_1077), .C(n_1079), .Y(n_1075) );
AND2x4_ASAP7_75t_L g357 ( .A(n_327), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g564 ( .A(n_327), .B(n_565), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_327), .A2(n_357), .B1(n_509), .B2(n_642), .C(n_657), .Y(n_656) );
AOI222xp33_ASAP7_75t_L g922 ( .A1(n_327), .A2(n_568), .B1(n_570), .B2(n_899), .C1(n_900), .C2(n_923), .Y(n_922) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g366 ( .A(n_328), .B(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g372 ( .A(n_328), .B(n_373), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_328), .A2(n_501), .B(n_504), .C(n_508), .Y(n_500) );
OR2x2_ASAP7_75t_L g767 ( .A(n_328), .B(n_403), .Y(n_767) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_SL g530 ( .A(n_332), .Y(n_530) );
INVx2_ASAP7_75t_L g811 ( .A(n_332), .Y(n_811) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g713 ( .A(n_334), .Y(n_713) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g1351 ( .A(n_335), .Y(n_1351) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g719 ( .A(n_338), .Y(n_719) );
BUFx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x6_ASAP7_75t_L g1353 ( .A(n_339), .B(n_1337), .Y(n_1353) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_348), .B1(n_356), .B2(n_359), .C(n_360), .Y(n_340) );
BUFx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g815 ( .A(n_343), .Y(n_815) );
BUFx3_ASAP7_75t_L g823 ( .A(n_343), .Y(n_823) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_SL g560 ( .A(n_347), .Y(n_560) );
BUFx3_ASAP7_75t_L g667 ( .A(n_347), .Y(n_667) );
INVx1_ASAP7_75t_L g696 ( .A(n_347), .Y(n_696) );
INVx2_ASAP7_75t_L g951 ( .A(n_347), .Y(n_951) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g934 ( .A(n_351), .Y(n_934) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_355), .Y(n_503) );
INVx2_ASAP7_75t_L g661 ( .A(n_355), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_355), .Y(n_663) );
INVx1_ASAP7_75t_L g924 ( .A(n_355), .Y(n_924) );
AND2x6_ASAP7_75t_L g1344 ( .A(n_355), .B(n_1331), .Y(n_1344) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_356), .A2(n_360), .B1(n_821), .B2(n_822), .C(n_828), .Y(n_820) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_SL g549 ( .A(n_357), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g845 ( .A1(n_357), .A2(n_509), .B1(n_846), .B2(n_848), .C(n_850), .Y(n_845) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_357), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g1084 ( .A1(n_357), .A2(n_509), .B1(n_1085), .B2(n_1086), .C(n_1088), .Y(n_1084) );
BUFx4f_ASAP7_75t_L g507 ( .A(n_358), .Y(n_507) );
AND2x4_ASAP7_75t_L g509 ( .A(n_358), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g679 ( .A(n_358), .Y(n_679) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_358), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_358), .A2(n_565), .B1(n_920), .B2(n_926), .Y(n_925) );
INVx2_ASAP7_75t_SL g931 ( .A(n_358), .Y(n_931) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g812 ( .A(n_362), .B(n_719), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_370), .B2(n_371), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_365), .A2(n_371), .B1(n_831), .B2(n_832), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_365), .A2(n_371), .B1(n_852), .B2(n_853), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_365), .A2(n_371), .B1(n_1051), .B2(n_1053), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_365), .A2(n_371), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
INVx6_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g552 ( .A(n_367), .Y(n_552) );
INVx1_ASAP7_75t_L g660 ( .A(n_367), .Y(n_660) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
AND2x2_ASAP7_75t_L g517 ( .A(n_368), .B(n_369), .Y(n_517) );
INVx4_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g675 ( .A(n_373), .Y(n_675) );
INVx1_ASAP7_75t_L g578 ( .A(n_374), .Y(n_578) );
AOI31xp33_ASAP7_75t_SL g921 ( .A1(n_374), .A2(n_922), .A3(n_927), .B(n_936), .Y(n_921) );
OAI31xp33_ASAP7_75t_L g971 ( .A1(n_374), .A2(n_972), .A3(n_991), .B(n_1005), .Y(n_971) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_375), .A2(n_836), .B1(n_854), .B2(n_855), .Y(n_835) );
NOR2xp67_ASAP7_75t_L g1011 ( .A(n_375), .B(n_1012), .Y(n_1011) );
AOI22xp5_ASAP7_75t_L g1073 ( .A1(n_375), .A2(n_1069), .B1(n_1074), .B2(n_1092), .Y(n_1073) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g425 ( .A(n_376), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g581 ( .A(n_376), .B(n_426), .Y(n_581) );
AND2x2_ASAP7_75t_L g598 ( .A(n_376), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g695 ( .A(n_376), .B(n_696), .Y(n_695) );
OR2x6_ASAP7_75t_L g950 ( .A(n_376), .B(n_951), .Y(n_950) );
BUFx2_ASAP7_75t_L g1438 ( .A(n_376), .Y(n_1438) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x6_ASAP7_75t_L g472 ( .A(n_377), .B(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g536 ( .A(n_377), .Y(n_536) );
AND4x1_ASAP7_75t_L g378 ( .A(n_379), .B(n_395), .C(n_409), .D(n_422), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_384), .B1(n_385), .B2(n_389), .C(n_390), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_380), .A2(n_385), .B1(n_390), .B2(n_538), .C(n_539), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_380), .A2(n_385), .B1(n_390), .B2(n_567), .C(n_569), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_380), .A2(n_390), .B(n_654), .Y(n_688) );
INVx1_ASAP7_75t_L g785 ( .A(n_380), .Y(n_785) );
AOI221xp5_ASAP7_75t_L g898 ( .A1(n_380), .A2(n_385), .B1(n_390), .B2(n_899), .C(n_900), .Y(n_898) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
AND2x2_ASAP7_75t_L g987 ( .A(n_381), .B(n_988), .Y(n_987) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g758 ( .A(n_382), .Y(n_758) );
AND2x4_ASAP7_75t_L g385 ( .A(n_383), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g390 ( .A(n_383), .B(n_391), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_383), .B(n_618), .Y(n_617) );
NAND2x1_ASAP7_75t_SL g866 ( .A(n_383), .B(n_757), .Y(n_866) );
NAND2x1p5_ASAP7_75t_L g869 ( .A(n_383), .B(n_408), .Y(n_869) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_385), .Y(n_782) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_388), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g630 ( .A(n_388), .B(n_471), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g781 ( .A1(n_390), .A2(n_782), .B1(n_783), .B2(n_784), .C(n_786), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_391), .A2(n_412), .B1(n_913), .B2(n_914), .Y(n_912) );
BUFx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx3_ASAP7_75t_L g408 ( .A(n_392), .Y(n_408) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_392), .Y(n_433) );
BUFx3_ASAP7_75t_L g585 ( .A(n_392), .Y(n_585) );
BUFx6f_ASAP7_75t_L g983 ( .A(n_392), .Y(n_983) );
AND2x4_ASAP7_75t_L g1363 ( .A(n_392), .B(n_1364), .Y(n_1363) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_406), .B2(n_407), .Y(n_395) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g687 ( .A(n_398), .Y(n_687) );
BUFx2_ASAP7_75t_L g789 ( .A(n_398), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_398), .A2(n_407), .B1(n_859), .B2(n_860), .Y(n_858) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_398), .Y(n_1027) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
INVx2_ASAP7_75t_L g911 ( .A(n_399), .Y(n_911) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx3_ASAP7_75t_L g462 ( .A(n_400), .Y(n_462) );
BUFx6f_ASAP7_75t_L g749 ( .A(n_400), .Y(n_749) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
INVx1_ASAP7_75t_L g595 ( .A(n_401), .Y(n_595) );
INVx1_ASAP7_75t_L g1376 ( .A(n_401), .Y(n_1376) );
AND2x6_ASAP7_75t_L g407 ( .A(n_402), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g411 ( .A(n_402), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g416 ( .A(n_402), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g488 ( .A(n_402), .B(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g493 ( .A(n_402), .B(n_417), .Y(n_493) );
AND2x2_ASAP7_75t_L g495 ( .A(n_402), .B(n_433), .Y(n_495) );
AND2x2_ASAP7_75t_L g498 ( .A(n_402), .B(n_462), .Y(n_498) );
AND2x2_ASAP7_75t_L g603 ( .A(n_402), .B(n_417), .Y(n_603) );
AND2x2_ASAP7_75t_L g794 ( .A(n_402), .B(n_417), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g909 ( .A1(n_402), .A2(n_598), .B1(n_910), .B2(n_915), .Y(n_909) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g444 ( .A(n_403), .Y(n_444) );
INVx2_ASAP7_75t_L g729 ( .A(n_404), .Y(n_729) );
AND2x2_ASAP7_75t_L g731 ( .A(n_404), .B(n_418), .Y(n_731) );
AND2x4_ASAP7_75t_L g993 ( .A(n_404), .B(n_430), .Y(n_993) );
INVx1_ASAP7_75t_L g446 ( .A(n_405), .Y(n_446) );
INVx1_ASAP7_75t_L g474 ( .A(n_405), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_407), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_407), .A2(n_1026), .B1(n_1027), .B2(n_1028), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_407), .A2(n_789), .B1(n_1082), .B2(n_1096), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_415), .B2(n_416), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_411), .A2(n_602), .B1(n_603), .B2(n_604), .C(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g685 ( .A(n_411), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_411), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_411), .A2(n_794), .B1(n_862), .B2(n_863), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_411), .A2(n_416), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_411), .A2(n_794), .B1(n_1083), .B2(n_1098), .Y(n_1097) );
BUFx3_ASAP7_75t_L g441 ( .A(n_412), .Y(n_441) );
BUFx2_ASAP7_75t_L g583 ( .A(n_412), .Y(n_583) );
INVx1_ASAP7_75t_L g1394 ( .A(n_412), .Y(n_1394) );
INVx2_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g489 ( .A(n_413), .Y(n_489) );
INVx2_ASAP7_75t_L g763 ( .A(n_413), .Y(n_763) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_414), .Y(n_430) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g588 ( .A(n_418), .Y(n_588) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_418), .Y(n_747) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_418), .Y(n_800) );
AND2x4_ASAP7_75t_L g1371 ( .A(n_418), .B(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1423 ( .A(n_418), .Y(n_1423) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g619 ( .A(n_419), .Y(n_619) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI33xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_427), .A3(n_434), .B1(n_437), .B2(n_440), .B3(n_442), .Y(n_422) );
AOI33xp33_ASAP7_75t_L g795 ( .A1(n_423), .A2(n_442), .A3(n_796), .B1(n_798), .B2(n_803), .B3(n_804), .Y(n_795) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g1390 ( .A(n_425), .B(n_1391), .C(n_1392), .Y(n_1390) );
BUFx2_ASAP7_75t_SL g999 ( .A(n_426), .Y(n_999) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g597 ( .A(n_429), .Y(n_597) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g751 ( .A(n_430), .Y(n_751) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g797 ( .A(n_432), .Y(n_797) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx4_ASAP7_75t_L g439 ( .A(n_436), .Y(n_439) );
INVx2_ASAP7_75t_SL g485 ( .A(n_436), .Y(n_485) );
INVx2_ASAP7_75t_SL g802 ( .A(n_436), .Y(n_802) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_439), .A2(n_622), .B1(n_623), .B2(n_626), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_439), .A2(n_1076), .B1(n_1091), .B2(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
INVx2_ASAP7_75t_L g645 ( .A(n_442), .Y(n_645) );
INVx6_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx5_ASAP7_75t_L g889 ( .A(n_443), .Y(n_889) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx2_ASAP7_75t_L g599 ( .A(n_445), .Y(n_599) );
BUFx2_ASAP7_75t_L g984 ( .A(n_445), .Y(n_984) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g1365 ( .A(n_446), .Y(n_1365) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_542), .B2(n_543), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g541 ( .A(n_452), .Y(n_541) );
NAND4xp75_ASAP7_75t_L g452 ( .A(n_453), .B(n_490), .C(n_499), .D(n_537), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_459), .B2(n_460), .Y(n_454) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g635 ( .A(n_457), .Y(n_635) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g483 ( .A(n_458), .Y(n_483) );
INVx1_ASAP7_75t_L g625 ( .A(n_458), .Y(n_625) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g590 ( .A(n_462), .Y(n_590) );
INVx1_ASAP7_75t_L g636 ( .A(n_462), .Y(n_636) );
INVx2_ASAP7_75t_L g880 ( .A(n_462), .Y(n_880) );
INVx2_ASAP7_75t_L g917 ( .A(n_462), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_467), .B2(n_468), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_465), .A2(n_628), .B1(n_629), .B2(n_631), .Y(n_627) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_467), .A2(n_524), .B(n_526), .C(n_528), .Y(n_523) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_468), .A2(n_872), .B1(n_875), .B2(n_876), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g1101 ( .A1(n_468), .A2(n_1039), .B1(n_1102), .B2(n_1103), .Y(n_1101) );
BUFx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g475 ( .A1(n_469), .A2(n_476), .B1(n_477), .B2(n_478), .Y(n_475) );
INVx2_ASAP7_75t_L g644 ( .A(n_469), .Y(n_644) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI33xp33_ASAP7_75t_L g870 ( .A1(n_472), .A2(n_871), .A3(n_877), .B1(n_882), .B2(n_885), .B3(n_888), .Y(n_870) );
OAI33xp33_ASAP7_75t_L g1036 ( .A1(n_472), .A2(n_888), .A3(n_1037), .B1(n_1042), .B2(n_1046), .B3(n_1052), .Y(n_1036) );
OAI33xp33_ASAP7_75t_L g1100 ( .A1(n_472), .A2(n_888), .A3(n_1101), .B1(n_1104), .B2(n_1107), .B3(n_1109), .Y(n_1100) );
INVx1_ASAP7_75t_L g1372 ( .A(n_474), .Y(n_1372) );
OAI22xp33_ASAP7_75t_L g1109 ( .A1(n_476), .A2(n_1085), .B1(n_1090), .B2(n_1110), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_477), .A2(n_484), .B1(n_502), .B2(n_503), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_478), .A2(n_480), .B1(n_505), .B2(n_507), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_484), .B2(n_485), .Y(n_479) );
BUFx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g878 ( .A(n_482), .Y(n_878) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g1432 ( .A(n_483), .Y(n_1432) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g981 ( .A(n_489), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_489), .B(n_988), .Y(n_1012) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_491), .B(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g615 ( .A(n_493), .Y(n_615) );
INVxp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g606 ( .A(n_495), .Y(n_606) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_511), .A3(n_529), .B(n_535), .Y(n_499) );
HB1xp67_ASAP7_75t_L g1443 ( .A(n_502), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_505), .B(n_1459), .Y(n_1458) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_SL g698 ( .A(n_506), .Y(n_698) );
INVx1_ASAP7_75t_L g929 ( .A(n_506), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g1444 ( .A1(n_506), .A2(n_924), .B1(n_1433), .B2(n_1434), .Y(n_1444) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g561 ( .A(n_509), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g927 ( .A1(n_509), .A2(n_928), .B(n_933), .Y(n_927) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_509), .A2(n_1054), .B1(n_1064), .B2(n_1065), .C(n_1066), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
OAI211xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_518), .C(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_517), .Y(n_525) );
INVx2_ASAP7_75t_L g772 ( .A(n_517), .Y(n_772) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_SL g576 ( .A(n_521), .Y(n_576) );
INVx1_ASAP7_75t_L g829 ( .A(n_521), .Y(n_829) );
BUFx2_ASAP7_75t_L g955 ( .A(n_524), .Y(n_955) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_SL g558 ( .A(n_525), .Y(n_558) );
INVx1_ASAP7_75t_L g573 ( .A(n_525), .Y(n_573) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g683 ( .A(n_535), .Y(n_683) );
AOI21x1_ASAP7_75t_L g725 ( .A1(n_535), .A2(n_726), .B(n_745), .Y(n_725) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g1057 ( .A(n_536), .Y(n_1057) );
AND2x4_ASAP7_75t_L g1357 ( .A(n_536), .B(n_1358), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_540), .A2(n_1152), .B1(n_1153), .B2(n_1154), .Y(n_1151) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g608 ( .A(n_545), .Y(n_608) );
NAND4xp75_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .C(n_579), .D(n_601), .Y(n_545) );
OAI31xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_562), .A3(n_577), .B(n_578), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_550) );
OAI221xp5_ASAP7_75t_L g963 ( .A1(n_551), .A2(n_573), .B1(n_964), .B2(n_965), .C(n_966), .Y(n_963) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g766 ( .A(n_552), .Y(n_766) );
INVx2_ASAP7_75t_L g818 ( .A(n_552), .Y(n_818) );
OAI21xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_559), .Y(n_556) );
INVx1_ASAP7_75t_L g827 ( .A(n_560), .Y(n_827) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_564), .A2(n_838), .B1(n_840), .B2(n_841), .C(n_842), .Y(n_837) );
INVx1_ASAP7_75t_L g658 ( .A(n_565), .Y(n_658) );
BUFx2_ASAP7_75t_L g958 ( .A(n_565), .Y(n_958) );
BUFx4f_ASAP7_75t_L g1403 ( .A(n_565), .Y(n_1403) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_569), .B2(n_570), .Y(n_566) );
INVx4_ASAP7_75t_L g653 ( .A(n_568), .Y(n_653) );
INVx2_ASAP7_75t_L g843 ( .A(n_568), .Y(n_843) );
AOI222xp33_ASAP7_75t_SL g648 ( .A1(n_570), .A2(n_649), .B1(n_651), .B2(n_652), .C1(n_654), .C2(n_655), .Y(n_648) );
INVx2_ASAP7_75t_SL g844 ( .A(n_570), .Y(n_844) );
INVx2_ASAP7_75t_L g1078 ( .A(n_570), .Y(n_1078) );
OAI211xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B(n_574), .C(n_575), .Y(n_571) );
BUFx2_ASAP7_75t_L g1447 ( .A(n_576), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_576), .B(n_1459), .Y(n_1461) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_580), .B(n_600), .Y(n_579) );
AOI33xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .A3(n_586), .B1(n_591), .B2(n_596), .B3(n_598), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g901 ( .A1(n_581), .A2(n_902), .B1(n_907), .B2(n_908), .Y(n_901) );
HB1xp67_ASAP7_75t_L g1361 ( .A(n_584), .Y(n_1361) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g753 ( .A(n_585), .B(n_728), .Y(n_753) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g884 ( .A(n_590), .Y(n_884) );
INVx2_ASAP7_75t_L g1050 ( .A(n_590), .Y(n_1050) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_593), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g727 ( .A(n_594), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_SL g752 ( .A(n_599), .Y(n_752) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AO22x2_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_689), .B1(n_690), .B2(n_773), .Y(n_610) );
INVx1_ASAP7_75t_L g773 ( .A(n_611), .Y(n_773) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_646), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_620), .Y(n_613) );
BUFx4f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx4f_ASAP7_75t_L g867 ( .A(n_617), .Y(n_867) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x6_ASAP7_75t_L g760 ( .A(n_619), .B(n_743), .Y(n_760) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g739 ( .A(n_625), .Y(n_739) );
OAI221xp5_ASAP7_75t_SL g662 ( .A1(n_626), .A2(n_631), .B1(n_659), .B2(n_663), .C(n_664), .Y(n_662) );
OR2x6_ASAP7_75t_L g742 ( .A(n_629), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g887 ( .A(n_629), .Y(n_887) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_629), .B(n_743), .Y(n_1004) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx3_ASAP7_75t_L g735 ( .A(n_630), .Y(n_735) );
BUFx2_ASAP7_75t_L g996 ( .A(n_630), .Y(n_996) );
INVx2_ASAP7_75t_L g1110 ( .A(n_630), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_636), .B2(n_637), .Y(n_632) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI22xp5_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_640), .B1(n_642), .B2(n_643), .Y(n_638) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g1052 ( .A1(n_643), .A2(n_1039), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI21xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_682), .B(n_684), .Y(n_646) );
NAND4xp25_ASAP7_75t_SL g647 ( .A(n_648), .B(n_656), .C(n_662), .D(n_668), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_649), .A2(n_907), .B1(n_937), .B2(n_940), .Y(n_936) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g768 ( .A(n_658), .B(n_767), .Y(n_768) );
BUFx2_ASAP7_75t_L g953 ( .A(n_659), .Y(n_953) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g1451 ( .A(n_663), .Y(n_1451) );
BUFx3_ASAP7_75t_L g670 ( .A(n_665), .Y(n_670) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g932 ( .A(n_667), .Y(n_932) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B1(n_672), .B2(n_676), .C(n_677), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g849 ( .A(n_674), .Y(n_849) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI31xp33_ASAP7_75t_L g807 ( .A1(n_683), .A2(n_808), .A3(n_820), .B(n_830), .Y(n_807) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NOR4xp75_ASAP7_75t_L g691 ( .A(n_692), .B(n_725), .C(n_764), .D(n_769), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_710), .Y(n_692) );
AOI33xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_697), .A3(n_699), .B1(n_701), .B2(n_705), .B3(n_709), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g1397 ( .A(n_694), .B(n_1398), .C(n_1399), .Y(n_1397) );
INVx3_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g825 ( .A(n_700), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_700), .B(n_724), .Y(n_1456) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g839 ( .A(n_704), .Y(n_839) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g770 ( .A(n_708), .B(n_767), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g1400 ( .A(n_709), .B(n_1401), .C(n_1402), .Y(n_1400) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_716), .B1(n_717), .B2(n_720), .C(n_721), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_712), .Y(n_970) );
INVx2_ASAP7_75t_L g1454 ( .A(n_712), .Y(n_1454) );
NAND2x1p5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
OR2x6_ASAP7_75t_L g718 ( .A(n_715), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g724 ( .A(n_715), .Y(n_724) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_715), .B(n_719), .Y(n_1455) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g968 ( .A(n_721), .Y(n_968) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI221x1_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_730), .B1(n_731), .B2(n_732), .C(n_733), .Y(n_726) );
INVx3_ASAP7_75t_L g1007 ( .A(n_727), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_727), .A2(n_731), .B1(n_1427), .B2(n_1428), .Y(n_1426) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx3_ASAP7_75t_L g1006 ( .A(n_731), .Y(n_1006) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_738), .B(n_742), .Y(n_733) );
OAI21xp5_ASAP7_75t_SL g734 ( .A1(n_735), .A2(n_736), .B(n_737), .Y(n_734) );
INVx2_ASAP7_75t_L g976 ( .A(n_739), .Y(n_976) );
INVx1_ASAP7_75t_L g759 ( .A(n_743), .Y(n_759) );
INVx1_ASAP7_75t_L g988 ( .A(n_743), .Y(n_988) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI221xp5_ASAP7_75t_SL g745 ( .A1(n_746), .A2(n_750), .B1(n_753), .B2(n_754), .C(n_755), .Y(n_745) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g903 ( .A(n_749), .Y(n_903) );
INVx2_ASAP7_75t_L g1388 ( .A(n_749), .Y(n_1388) );
INVx8_ASAP7_75t_L g973 ( .A(n_753), .Y(n_973) );
NAND2x1p5_ASAP7_75t_L g756 ( .A(n_757), .B(n_759), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
CKINVDCx11_ASAP7_75t_R g990 ( .A(n_760), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
OR2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
OR2x6_ASAP7_75t_L g771 ( .A(n_767), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g1459 ( .A(n_767), .Y(n_1459) );
OAI221xp5_ASAP7_75t_L g817 ( .A1(n_772), .A2(n_790), .B1(n_792), .B2(n_818), .C(n_819), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_1017), .B1(n_1111), .B2(n_1113), .Y(n_774) );
INVx1_ASAP7_75t_L g1113 ( .A(n_775), .Y(n_1113) );
XNOR2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_893), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_833), .B2(n_892), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_805), .Y(n_779) );
AND4x1_ASAP7_75t_L g780 ( .A(n_781), .B(n_787), .C(n_791), .D(n_795), .Y(n_780) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
BUFx3_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI22xp5_ASAP7_75t_SL g1000 ( .A1(n_802), .A2(n_1001), .B1(n_1002), .B2(n_1003), .Y(n_1000) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx3_ASAP7_75t_L g892 ( .A(n_833), .Y(n_892) );
INVx1_ASAP7_75t_L g890 ( .A(n_834), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_856), .Y(n_834) );
NAND3xp33_ASAP7_75t_L g836 ( .A(n_837), .B(n_845), .C(n_851), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_841), .A2(n_853), .B1(n_878), .B2(n_883), .Y(n_882) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_850), .A2(n_852), .B1(n_872), .B2(n_886), .Y(n_885) );
NOR3xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_864), .C(n_870), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_858), .B(n_861), .Y(n_857) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g1034 ( .A(n_866), .Y(n_1034) );
BUFx3_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
BUFx2_ASAP7_75t_L g1035 ( .A(n_869), .Y(n_1035) );
INVx2_ASAP7_75t_SL g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g1039 ( .A(n_873), .Y(n_1039) );
INVx2_ASAP7_75t_SL g873 ( .A(n_874), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B1(n_880), .B2(n_881), .Y(n_877) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_878), .A2(n_1043), .B1(n_1044), .B2(n_1045), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_878), .A2(n_1045), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
CKINVDCx8_ASAP7_75t_R g888 ( .A(n_889), .Y(n_888) );
NAND3xp33_ASAP7_75t_L g1386 ( .A(n_889), .B(n_1387), .C(n_1389), .Y(n_1386) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_945), .B1(n_946), .B2(n_1016), .Y(n_893) );
INVx1_ASAP7_75t_L g1016 ( .A(n_894), .Y(n_1016) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
NAND2xp5_ASAP7_75t_SL g895 ( .A(n_896), .B(n_941), .Y(n_895) );
INVx1_ASAP7_75t_L g943 ( .A(n_897), .Y(n_943) );
NAND3xp33_ASAP7_75t_SL g897 ( .A(n_898), .B(n_901), .C(n_909), .Y(n_897) );
INVx1_ASAP7_75t_L g1045 ( .A(n_903), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_911), .A2(n_1431), .B1(n_1433), .B2(n_1434), .Y(n_1430) );
INVx1_ASAP7_75t_L g978 ( .A(n_916), .Y(n_978) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g942 ( .A(n_921), .Y(n_942) );
INVx1_ASAP7_75t_L g935 ( .A(n_924), .Y(n_935) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g1087 ( .A(n_931), .Y(n_1087) );
NAND3xp33_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .C(n_944), .Y(n_941) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
AND4x1_ASAP7_75t_L g947 ( .A(n_948), .B(n_971), .C(n_1008), .D(n_1013), .Y(n_947) );
NOR3xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_968), .C(n_969), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_952), .B1(n_961), .B2(n_963), .Y(n_949) );
INVx2_ASAP7_75t_L g1445 ( .A(n_950), .Y(n_1445) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_954), .B1(n_955), .B2(n_956), .C(n_957), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g994 ( .A1(n_954), .A2(n_956), .B1(n_995), .B2(n_997), .C(n_999), .Y(n_994) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx4_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
AOI221xp5_ASAP7_75t_L g1441 ( .A1(n_962), .A2(n_1442), .B1(n_1445), .B2(n_1446), .C(n_1452), .Y(n_1441) );
OAI221xp5_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_977), .B1(n_978), .B2(n_979), .C(n_980), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx2_ASAP7_75t_L g1002 ( .A(n_976), .Y(n_1002) );
INVx1_ASAP7_75t_L g1047 ( .A(n_976), .Y(n_1047) );
INVx2_ASAP7_75t_L g1108 ( .A(n_976), .Y(n_1108) );
BUFx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx2_ASAP7_75t_SL g1396 ( .A(n_983), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_987), .B1(n_989), .B2(n_990), .Y(n_985) );
CKINVDCx6p67_ASAP7_75t_R g992 ( .A(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1041 ( .A(n_996), .Y(n_1041) );
INVx2_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1010), .B(n_1440), .Y(n_1439) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1015), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1018), .Y(n_1112) );
AO22x2_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1020), .B1(n_1070), .B2(n_1071), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
XNOR2xp5_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1022), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1055), .Y(n_1022) );
NOR3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1032), .C(n_1036), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1029), .Y(n_1024) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1039), .B1(n_1040), .B2(n_1041), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1048), .B1(n_1049), .B2(n_1051), .Y(n_1046) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
AOI22xp5_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1058), .B1(n_1068), .B2(n_1069), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
NAND3xp33_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1063), .C(n_1067), .Y(n_1058) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1093), .Y(n_1072) );
NAND3xp33_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1084), .C(n_1089), .Y(n_1074) );
NOR3xp33_ASAP7_75t_SL g1093 ( .A(n_1094), .B(n_1099), .C(n_1100), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1097), .Y(n_1094) );
OAI21xp5_ASAP7_75t_SL g1435 ( .A1(n_1110), .A2(n_1436), .B(n_1437), .Y(n_1435) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
OAI221xp5_ASAP7_75t_L g1114 ( .A1(n_1115), .A2(n_1320), .B1(n_1321), .B2(n_1404), .C(n_1409), .Y(n_1114) );
AOI221xp5_ASAP7_75t_L g1115 ( .A1(n_1116), .A2(n_1201), .B1(n_1264), .B2(n_1265), .C(n_1293), .Y(n_1115) );
A2O1A1Ixp33_ASAP7_75t_SL g1116 ( .A1(n_1117), .A2(n_1155), .B(n_1183), .C(n_1194), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1139), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1119), .B(n_1214), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1119), .B(n_1181), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1119), .B(n_1222), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1119), .B(n_1274), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1119), .B(n_1243), .Y(n_1308) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1120), .B(n_1160), .Y(n_1159) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1120), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1120), .B(n_1205), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1120), .B(n_1232), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1120), .B(n_1161), .Y(n_1236) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1120), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1120), .B(n_1140), .Y(n_1289) );
AOI211xp5_ASAP7_75t_L g1296 ( .A1(n_1120), .A2(n_1208), .B(n_1297), .C(n_1298), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1120), .B(n_1239), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1133), .Y(n_1120) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1128), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1124), .B(n_1129), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1127), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1127), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1130 ( .A(n_1128), .B(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1129), .B(n_1132), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1188 ( .A(n_1130), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1466 ( .A(n_1131), .Y(n_1466) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1134), .Y(n_1173) );
BUFx3_ASAP7_75t_L g1195 ( .A(n_1134), .Y(n_1195) );
AND2x4_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1137), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1135), .B(n_1137), .Y(n_1144) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_1136), .B(n_1137), .Y(n_1138) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1138), .Y(n_1175) );
O2A1O1Ixp33_ASAP7_75t_L g1283 ( .A1(n_1139), .A2(n_1246), .B(n_1284), .C(n_1287), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1145), .Y(n_1139) );
NOR2x1_ASAP7_75t_L g1208 ( .A(n_1140), .B(n_1182), .Y(n_1208) );
AOI21xp5_ASAP7_75t_L g1237 ( .A1(n_1140), .A2(n_1238), .B(n_1241), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1243 ( .A(n_1140), .B(n_1146), .Y(n_1243) );
BUFx2_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
BUFx3_ASAP7_75t_L g1160 ( .A(n_1141), .Y(n_1160) );
INVxp67_ASAP7_75t_L g1206 ( .A(n_1141), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1141), .B(n_1250), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1145), .B(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1145), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1150), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g1266 ( .A1(n_1146), .A2(n_1267), .B1(n_1271), .B2(n_1273), .Y(n_1266) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1147), .B(n_1150), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1147), .B(n_1182), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1147), .B(n_1160), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1147), .B(n_1150), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1315 ( .A(n_1147), .B(n_1160), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1149), .Y(n_1147) );
INVx2_ASAP7_75t_SL g1182 ( .A(n_1150), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1150), .B(n_1160), .Y(n_1232) );
BUFx6f_ASAP7_75t_L g1167 ( .A(n_1152), .Y(n_1167) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1154), .Y(n_1170) );
AOI21xp5_ASAP7_75t_L g1155 ( .A1(n_1156), .A2(n_1162), .B(n_1177), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1161), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1282 ( .A(n_1159), .B(n_1251), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1160), .B(n_1181), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1160), .B(n_1256), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1160), .B(n_1257), .Y(n_1297) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1161), .Y(n_1256) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1161), .B(n_1289), .Y(n_1288) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1163), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_1163), .A2(n_1227), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1163), .B(n_1178), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1163), .B(n_1301), .Y(n_1300) );
INVx2_ASAP7_75t_SL g1163 ( .A(n_1164), .Y(n_1163) );
AND2x4_ASAP7_75t_L g1227 ( .A(n_1164), .B(n_1223), .Y(n_1227) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1164), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1248 ( .A(n_1164), .B(n_1249), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1164), .B(n_1218), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1164), .B(n_1191), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g1281 ( .A(n_1164), .Y(n_1281) );
CKINVDCx5p33_ASAP7_75t_R g1164 ( .A(n_1165), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1165), .B(n_1191), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1165), .B(n_1223), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1172), .Y(n_1165) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1168), .B1(n_1169), .B2(n_1171), .Y(n_1166) );
BUFx3_ASAP7_75t_L g1198 ( .A(n_1167), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1200 ( .A(n_1169), .Y(n_1200) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_1173), .A2(n_1174), .B1(n_1175), .B2(n_1176), .Y(n_1172) );
INVx2_ASAP7_75t_L g1190 ( .A(n_1175), .Y(n_1190) );
NOR2xp33_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1179), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1178), .B(n_1221), .Y(n_1220) );
O2A1O1Ixp33_ASAP7_75t_L g1224 ( .A1(n_1178), .A2(n_1182), .B(n_1225), .C(n_1226), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1178), .B(n_1250), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1178), .B(n_1227), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1178), .B(n_1232), .Y(n_1292) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1180), .B(n_1249), .Y(n_1306) );
OAI21xp5_ASAP7_75t_L g1312 ( .A1(n_1180), .A2(n_1240), .B(n_1292), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1181), .B(n_1206), .Y(n_1230) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1181), .Y(n_1269) );
OAI32xp33_ASAP7_75t_L g1215 ( .A1(n_1182), .A2(n_1216), .A3(n_1217), .B1(n_1219), .B2(n_1222), .Y(n_1215) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1191), .Y(n_1184) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1185), .Y(n_1212) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1185), .Y(n_1218) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1186), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1263 ( .A(n_1186), .B(n_1191), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1186), .B(n_1223), .Y(n_1286) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1186), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1189), .Y(n_1186) );
INVx3_ASAP7_75t_L g1223 ( .A(n_1191), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1193), .Y(n_1191) );
INVx3_ASAP7_75t_L g1252 ( .A(n_1194), .Y(n_1252) );
OAI21xp5_ASAP7_75t_L g1303 ( .A1(n_1194), .A2(n_1274), .B(n_1304), .Y(n_1303) );
OAI22xp33_ASAP7_75t_L g1196 ( .A1(n_1197), .A2(n_1198), .B1(n_1199), .B2(n_1200), .Y(n_1196) );
BUFx2_ASAP7_75t_SL g1320 ( .A(n_1200), .Y(n_1320) );
NAND5xp2_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1207), .C(n_1228), .D(n_1237), .E(n_1253), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1205), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1206), .B(n_1236), .Y(n_1235) );
AOI211xp5_ASAP7_75t_L g1207 ( .A1(n_1208), .A2(n_1209), .B(n_1215), .C(n_1224), .Y(n_1207) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1210), .B(n_1255), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1213), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1212), .Y(n_1245) );
O2A1O1Ixp33_ASAP7_75t_L g1299 ( .A1(n_1212), .A2(n_1235), .B(n_1300), .C(n_1302), .Y(n_1299) );
OAI22xp5_ASAP7_75t_SL g1260 ( .A1(n_1213), .A2(n_1261), .B1(n_1262), .B2(n_1263), .Y(n_1260) );
A2O1A1Ixp33_ASAP7_75t_L g1287 ( .A1(n_1213), .A2(n_1288), .B(n_1290), .C(n_1291), .Y(n_1287) );
A2O1A1Ixp33_ASAP7_75t_L g1310 ( .A1(n_1213), .A2(n_1282), .B(n_1311), .C(n_1312), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1213 ( .A(n_1214), .Y(n_1213) );
AOI22xp5_ASAP7_75t_L g1228 ( .A1(n_1217), .A2(n_1229), .B1(n_1233), .B2(n_1235), .Y(n_1228) );
OAI211xp5_ASAP7_75t_SL g1265 ( .A1(n_1217), .A2(n_1266), .B(n_1275), .C(n_1283), .Y(n_1265) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1218), .B(n_1227), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1218), .B(n_1234), .Y(n_1304) );
OAI322xp33_ASAP7_75t_L g1313 ( .A1(n_1219), .A2(n_1226), .A3(n_1262), .B1(n_1263), .B2(n_1314), .C1(n_1316), .C2(n_1318), .Y(n_1313) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1221), .Y(n_1262) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
NAND3xp33_ASAP7_75t_L g1247 ( .A(n_1223), .B(n_1248), .C(n_1250), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1223), .B(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx2_ASAP7_75t_L g1277 ( .A(n_1230), .Y(n_1277) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1234), .B(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1238), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1240), .Y(n_1238) );
OAI211xp5_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1244), .B(n_1247), .C(n_1252), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1246), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1250), .B(n_1289), .Y(n_1301) );
NOR2xp33_ASAP7_75t_SL g1314 ( .A(n_1250), .B(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1252), .Y(n_1264) );
O2A1O1Ixp33_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1257), .B(n_1258), .C(n_1260), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
OAI21xp5_ASAP7_75t_L g1307 ( .A1(n_1257), .A2(n_1298), .B(n_1308), .Y(n_1307) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1270), .Y(n_1268) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
O2A1O1Ixp33_ASAP7_75t_L g1275 ( .A1(n_1276), .A2(n_1277), .B(n_1278), .C(n_1280), .Y(n_1275) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1276), .Y(n_1290) );
OAI21xp5_ASAP7_75t_L g1291 ( .A1(n_1277), .A2(n_1286), .B(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1282), .Y(n_1280) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
OAI211xp5_ASAP7_75t_SL g1293 ( .A1(n_1294), .A2(n_1296), .B(n_1299), .C(n_1309), .Y(n_1293) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1301), .Y(n_1311) );
OAI21xp5_ASAP7_75t_L g1302 ( .A1(n_1303), .A2(n_1305), .B(n_1307), .Y(n_1302) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
NOR3xp33_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1313), .C(n_1319), .Y(n_1309) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVxp67_ASAP7_75t_SL g1321 ( .A(n_1322), .Y(n_1321) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
AOI221xp5_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1357), .B1(n_1359), .B2(n_1383), .C(n_1385), .Y(n_1326) );
NAND4xp25_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1338), .C(n_1345), .D(n_1354), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_1329), .A2(n_1330), .B1(n_1334), .B2(n_1335), .Y(n_1328) );
AND2x4_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1333), .Y(n_1330) );
INVx1_ASAP7_75t_SL g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1336), .Y(n_1356) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_1339), .A2(n_1340), .B1(n_1343), .B2(n_1344), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_1339), .A2(n_1379), .B1(n_1380), .B2(n_1381), .Y(n_1378) );
AND2x2_ASAP7_75t_SL g1349 ( .A(n_1341), .B(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
AOI222xp33_ASAP7_75t_L g1345 ( .A1(n_1346), .A2(n_1347), .B1(n_1348), .B2(n_1349), .C1(n_1352), .C2(n_1353), .Y(n_1345) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
CKINVDCx8_ASAP7_75t_R g1354 ( .A(n_1355), .Y(n_1354) );
NAND3xp33_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1370), .C(n_1378), .Y(n_1359) );
AOI211xp5_ASAP7_75t_L g1360 ( .A1(n_1361), .A2(n_1362), .B(n_1363), .C(n_1366), .Y(n_1360) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_1371), .A2(n_1373), .B1(n_1374), .B2(n_1377), .Y(n_1370) );
AND2x4_ASAP7_75t_L g1374 ( .A(n_1372), .B(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx5_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
CKINVDCx16_ASAP7_75t_R g1383 ( .A(n_1384), .Y(n_1383) );
NAND4xp25_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1390), .C(n_1397), .D(n_1400), .Y(n_1385) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx2_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1403), .Y(n_1449) );
CKINVDCx5p33_ASAP7_75t_R g1404 ( .A(n_1405), .Y(n_1404) );
BUFx2_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
OAI21xp5_ASAP7_75t_L g1465 ( .A1(n_1411), .A2(n_1466), .B(n_1467), .Y(n_1465) );
INVxp33_ASAP7_75t_SL g1412 ( .A(n_1413), .Y(n_1412) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
HB1xp67_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
NAND4xp25_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1439), .C(n_1441), .D(n_1457), .Y(n_1417) );
OAI21xp5_ASAP7_75t_SL g1418 ( .A1(n_1419), .A2(n_1429), .B(n_1438), .Y(n_1418) );
AOI21xp5_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1424), .B(n_1425), .Y(n_1420) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
OAI22xp5_ASAP7_75t_L g1448 ( .A1(n_1427), .A2(n_1428), .B1(n_1449), .B2(n_1450), .Y(n_1448) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g1457 ( .A1(n_1458), .A2(n_1460), .B1(n_1461), .B2(n_1462), .C(n_1463), .Y(n_1457) );
HB1xp67_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
endmodule