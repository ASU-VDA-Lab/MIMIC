module real_aes_12343_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_552;
wire n_602;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_0), .A2(n_21), .B1(n_551), .B2(n_556), .Y(n_550) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_0), .A2(n_38), .B1(n_700), .B2(n_704), .Y(n_699) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_1), .A2(n_42), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g165 ( .A(n_1), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_2), .B(n_143), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_3), .A2(n_72), .B1(n_563), .B2(n_566), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_3), .A2(n_708), .B(n_709), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_4), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_5), .B(n_188), .Y(n_204) );
BUFx3_ASAP7_75t_L g526 ( .A(n_6), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_7), .B(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g627 ( .A(n_8), .Y(n_627) );
INVx1_ASAP7_75t_L g523 ( .A(n_9), .Y(n_523) );
INVx2_ASAP7_75t_L g643 ( .A(n_9), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_10), .B(n_162), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_11), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_12), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_13), .Y(n_229) );
INVx1_ASAP7_75t_L g95 ( .A(n_14), .Y(n_95) );
BUFx3_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_15), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g500 ( .A(n_15), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_16), .A2(n_48), .B1(n_584), .B2(n_587), .Y(n_583) );
INVx1_ASAP7_75t_L g650 ( .A(n_16), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_17), .Y(n_198) );
BUFx10_ASAP7_75t_L g521 ( .A(n_18), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_19), .B(n_117), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_20), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_21), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_22), .B(n_143), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_23), .A2(n_47), .B1(n_596), .B2(n_597), .Y(n_595) );
INVxp67_ASAP7_75t_SL g638 ( .A(n_23), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_24), .B(n_117), .Y(n_127) );
AND2x2_ASAP7_75t_L g574 ( .A(n_25), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g582 ( .A(n_25), .B(n_35), .Y(n_582) );
INVx1_ASAP7_75t_L g607 ( .A(n_25), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_26), .B(n_129), .Y(n_265) );
INVx1_ASAP7_75t_L g545 ( .A(n_26), .Y(n_545) );
NAND2xp33_ASAP7_75t_L g150 ( .A(n_27), .B(n_121), .Y(n_150) );
INVx1_ASAP7_75t_L g85 ( .A(n_28), .Y(n_85) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_29), .A2(n_218), .B(n_220), .C(n_222), .Y(n_217) );
INVx2_ASAP7_75t_L g555 ( .A(n_30), .Y(n_555) );
OAI21xp33_ASAP7_75t_L g577 ( .A1(n_31), .A2(n_566), .B(n_578), .Y(n_577) );
INVxp33_ASAP7_75t_SL g669 ( .A(n_31), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_32), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_33), .B(n_93), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_34), .B(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g575 ( .A(n_35), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_35), .B(n_607), .Y(n_606) );
AO221x1_ASAP7_75t_L g157 ( .A1(n_36), .A2(n_65), .B1(n_117), .B2(n_124), .C(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_37), .B(n_182), .Y(n_200) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_38), .A2(n_57), .B1(n_617), .B2(n_618), .C(n_621), .Y(n_616) );
AND2x4_ASAP7_75t_L g84 ( .A(n_39), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_39), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g269 ( .A(n_40), .B(n_222), .C(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g637 ( .A(n_41), .Y(n_637) );
INVx1_ASAP7_75t_L g645 ( .A(n_41), .Y(n_645) );
INVx1_ASAP7_75t_L g166 ( .A(n_42), .Y(n_166) );
INVx1_ASAP7_75t_L g113 ( .A(n_43), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_44), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_45), .A2(n_235), .B(n_236), .C(n_238), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_46), .A2(n_546), .B1(n_718), .B2(n_728), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_46), .Y(n_728) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_47), .Y(n_661) );
INVx1_ASAP7_75t_L g675 ( .A(n_48), .Y(n_675) );
INVx2_ASAP7_75t_L g237 ( .A(n_49), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_50), .B(n_111), .Y(n_206) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_51), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_52), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_53), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g615 ( .A(n_54), .Y(n_615) );
AND2x2_ASAP7_75t_L g191 ( .A(n_55), .B(n_111), .Y(n_191) );
INVx1_ASAP7_75t_L g169 ( .A(n_56), .Y(n_169) );
AOI211xp5_ASAP7_75t_L g680 ( .A1(n_57), .A2(n_681), .B(n_685), .C(n_691), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_58), .A2(n_63), .B1(n_505), .B2(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_58), .Y(n_505) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_59), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g161 ( .A1(n_60), .A2(n_62), .B1(n_143), .B2(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_61), .B(n_222), .Y(n_267) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_61), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_63), .Y(n_506) );
AOI21xp33_ASAP7_75t_L g599 ( .A1(n_64), .A2(n_600), .B(n_605), .Y(n_599) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_64), .Y(n_660) );
AND2x2_ASAP7_75t_L g244 ( .A(n_66), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g89 ( .A(n_67), .Y(n_89) );
BUFx3_ASAP7_75t_L g125 ( .A(n_67), .Y(n_125) );
INVx1_ASAP7_75t_L g146 ( .A(n_67), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g108 ( .A(n_68), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_69), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g554 ( .A(n_70), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g561 ( .A(n_70), .Y(n_561) );
INVxp67_ASAP7_75t_SL g603 ( .A(n_70), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_71), .B(n_182), .Y(n_264) );
INVx1_ASAP7_75t_L g686 ( .A(n_72), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_73), .B(n_111), .Y(n_153) );
INVx2_ASAP7_75t_L g528 ( .A(n_74), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_75), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_76), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_96), .B(n_492), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
BUFx2_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx3_ASAP7_75t_L g132 ( .A(n_84), .Y(n_132) );
BUFx6f_ASAP7_75t_SL g205 ( .A(n_84), .Y(n_205) );
INVx2_ASAP7_75t_L g215 ( .A(n_84), .Y(n_215) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_85), .Y(n_517) );
INVxp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AO21x2_ASAP7_75t_L g730 ( .A1(n_87), .A2(n_724), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_90), .Y(n_87) );
AOI21xp5_ASAP7_75t_SL g178 ( .A1(n_88), .A2(n_179), .B(n_180), .Y(n_178) );
BUFx3_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g190 ( .A(n_89), .Y(n_190) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g203 ( .A(n_94), .Y(n_203) );
INVx1_ASAP7_75t_L g227 ( .A(n_94), .Y(n_227) );
INVx2_ASAP7_75t_L g270 ( .A(n_94), .Y(n_270) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g118 ( .A(n_95), .Y(n_118) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NAND3x1_ASAP7_75t_L g97 ( .A(n_98), .B(n_380), .C(n_455), .Y(n_97) );
NOR2x1_ASAP7_75t_L g98 ( .A(n_99), .B(n_327), .Y(n_98) );
NAND3xp33_ASAP7_75t_L g99 ( .A(n_100), .B(n_297), .C(n_317), .Y(n_99) );
AOI221xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_171), .B1(n_249), .B2(n_258), .C(n_275), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_154), .Y(n_102) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_133), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g350 ( .A(n_105), .Y(n_350) );
AND2x2_ASAP7_75t_L g404 ( .A(n_105), .B(n_396), .Y(n_404) );
AND2x2_ASAP7_75t_L g485 ( .A(n_105), .B(n_156), .Y(n_485) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_106), .B(n_260), .Y(n_293) );
AND2x2_ASAP7_75t_L g427 ( .A(n_106), .B(n_156), .Y(n_427) );
INVx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g274 ( .A(n_107), .B(n_134), .Y(n_274) );
AND2x2_ASAP7_75t_L g278 ( .A(n_107), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g306 ( .A(n_107), .B(n_156), .Y(n_306) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_107), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_107), .B(n_134), .Y(n_361) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_114), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_111), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g136 ( .A(n_111), .Y(n_136) );
INVx2_ASAP7_75t_L g177 ( .A(n_111), .Y(n_177) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g195 ( .A(n_112), .Y(n_195) );
INVx1_ASAP7_75t_L g246 ( .A(n_112), .Y(n_246) );
INVx1_ASAP7_75t_L g167 ( .A(n_113), .Y(n_167) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_126), .B(n_131), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_119), .B(n_123), .Y(n_115) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx3_ASAP7_75t_L g149 ( .A(n_118), .Y(n_149) );
INVx2_ASAP7_75t_L g268 ( .A(n_120), .Y(n_268) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g129 ( .A(n_121), .Y(n_129) );
INVx3_ASAP7_75t_L g158 ( .A(n_121), .Y(n_158) );
INVx2_ASAP7_75t_L g188 ( .A(n_121), .Y(n_188) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_122), .Y(n_141) );
INVx2_ASAP7_75t_L g144 ( .A(n_122), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_123), .A2(n_225), .B(n_228), .Y(n_224) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g130 ( .A(n_125), .Y(n_130) );
INVx2_ASAP7_75t_L g222 ( .A(n_125), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B(n_130), .Y(n_126) );
O2A1O1Ixp5_ASAP7_75t_L g197 ( .A1(n_130), .A2(n_198), .B(n_199), .C(n_200), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_130), .A2(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
NOR2xp33_ASAP7_75t_R g163 ( .A(n_132), .B(n_164), .Y(n_163) );
OR2x2_ASAP7_75t_L g326 ( .A(n_133), .B(n_281), .Y(n_326) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g279 ( .A(n_134), .Y(n_279) );
INVx1_ASAP7_75t_L g291 ( .A(n_134), .Y(n_291) );
INVx1_ASAP7_75t_L g316 ( .A(n_134), .Y(n_316) );
AND2x2_ASAP7_75t_L g374 ( .A(n_134), .B(n_261), .Y(n_374) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_137), .B(n_153), .Y(n_134) );
INVx1_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_147), .B(n_152), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_142), .B(n_145), .Y(n_138) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g162 ( .A(n_141), .Y(n_162) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
INVx2_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
INVx2_ASAP7_75t_L g160 ( .A(n_145), .Y(n_160) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g151 ( .A(n_146), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_150), .B(n_151), .Y(n_147) );
INVx2_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
INVx2_ASAP7_75t_L g219 ( .A(n_149), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_149), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g238 ( .A(n_151), .Y(n_238) );
AND2x4_ASAP7_75t_L g176 ( .A(n_152), .B(n_177), .Y(n_176) );
AOI21xp33_ASAP7_75t_L g247 ( .A1(n_152), .A2(n_244), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g335 ( .A(n_154), .Y(n_335) );
OR2x2_ASAP7_75t_L g364 ( .A(n_154), .B(n_326), .Y(n_364) );
OR2x2_ASAP7_75t_L g383 ( .A(n_154), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g345 ( .A(n_155), .Y(n_345) );
AND2x2_ASAP7_75t_L g392 ( .A(n_155), .B(n_283), .Y(n_392) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_155), .Y(n_462) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g259 ( .A(n_156), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g280 ( .A(n_156), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g348 ( .A(n_156), .B(n_279), .Y(n_348) );
INVx2_ASAP7_75t_SL g396 ( .A(n_156), .Y(n_396) );
AO31x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .A3(n_163), .B(n_168), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_162), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
AOI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_167), .Y(n_164) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_166), .B(n_167), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVxp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_207), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_173), .B(n_332), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_173), .A2(n_367), .B1(n_374), .B2(n_375), .Y(n_373) );
AND2x2_ASAP7_75t_L g458 ( .A(n_173), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_192), .Y(n_173) );
INVx2_ASAP7_75t_L g253 ( .A(n_174), .Y(n_253) );
INVx1_ASAP7_75t_L g310 ( .A(n_174), .Y(n_310) );
OR2x2_ASAP7_75t_L g321 ( .A(n_174), .B(n_233), .Y(n_321) );
AND2x2_ASAP7_75t_L g416 ( .A(n_174), .B(n_193), .Y(n_416) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_175), .B(n_183), .Y(n_174) );
NAND2x1_ASAP7_75t_L g175 ( .A(n_176), .B(n_178), .Y(n_175) );
AOI21x1_ASAP7_75t_L g183 ( .A1(n_176), .A2(n_184), .B(n_191), .Y(n_183) );
O2A1O1Ixp5_ASAP7_75t_L g262 ( .A1(n_176), .A2(n_263), .B(n_266), .C(n_271), .Y(n_262) );
INVx2_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_187), .B(n_189), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_189), .A2(n_202), .B(n_204), .Y(n_201) );
INVx1_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
BUFx10_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g287 ( .A(n_192), .Y(n_287) );
INVx1_ASAP7_75t_L g301 ( .A(n_192), .Y(n_301) );
INVx1_ASAP7_75t_L g311 ( .A(n_192), .Y(n_311) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVxp33_ASAP7_75t_L g399 ( .A(n_193), .Y(n_399) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .B(n_206), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVxp67_ASAP7_75t_L g248 ( .A(n_195), .Y(n_248) );
OAI21x1_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_201), .B(n_205), .Y(n_196) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_207), .Y(n_329) );
INVx1_ASAP7_75t_L g428 ( .A(n_207), .Y(n_428) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_209), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g442 ( .A(n_209), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_232), .Y(n_209) );
INVx3_ASAP7_75t_L g257 ( .A(n_210), .Y(n_257) );
AND2x2_ASAP7_75t_L g341 ( .A(n_210), .B(n_287), .Y(n_341) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_216), .B(n_223), .Y(n_210) );
AO21x1_ASAP7_75t_SL g284 ( .A1(n_211), .A2(n_216), .B(n_223), .Y(n_284) );
INVxp67_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
OAI21x1_ASAP7_75t_SL g223 ( .A1(n_212), .A2(n_224), .B(n_230), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
INVx2_ASAP7_75t_L g231 ( .A(n_213), .Y(n_231) );
INVx2_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_L g235 ( .A(n_227), .Y(n_235) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g254 ( .A(n_233), .Y(n_254) );
INVx2_ASAP7_75t_L g286 ( .A(n_233), .Y(n_286) );
AND2x2_ASAP7_75t_L g296 ( .A(n_233), .B(n_253), .Y(n_296) );
AND2x2_ASAP7_75t_L g332 ( .A(n_233), .B(n_257), .Y(n_332) );
AND2x2_ASAP7_75t_L g412 ( .A(n_233), .B(n_252), .Y(n_412) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_239), .B(n_247), .Y(n_233) );
NOR2xp67_ASAP7_75t_L g236 ( .A(n_235), .B(n_237), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_243), .B(n_244), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_248), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
OR2x2_ASAP7_75t_L g480 ( .A(n_251), .B(n_301), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
OR2x2_ASAP7_75t_L g358 ( .A(n_252), .B(n_287), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_252), .B(n_256), .Y(n_489) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g365 ( .A(n_255), .Y(n_365) );
BUFx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g398 ( .A(n_257), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g405 ( .A(n_257), .B(n_286), .Y(n_405) );
OR2x2_ASAP7_75t_L g421 ( .A(n_257), .B(n_286), .Y(n_421) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_273), .Y(n_258) );
AND2x4_ASAP7_75t_L g360 ( .A(n_259), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g379 ( .A(n_259), .B(n_278), .Y(n_379) );
INVx2_ASAP7_75t_L g281 ( .A(n_260), .Y(n_281) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g305 ( .A(n_261), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_261), .B(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_SL g337 ( .A(n_261), .Y(n_337) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g393 ( .A(n_273), .Y(n_393) );
BUFx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g336 ( .A(n_274), .B(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_SL g410 ( .A(n_274), .B(n_396), .Y(n_410) );
AND2x2_ASAP7_75t_L g471 ( .A(n_274), .B(n_305), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_282), .B1(n_288), .B2(n_294), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_281), .B(n_451), .C(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g484 ( .A(n_281), .Y(n_484) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g295 ( .A(n_283), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g318 ( .A(n_283), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_SL g377 ( .A(n_283), .B(n_369), .Y(n_377) );
INVx5_ASAP7_75t_L g431 ( .A(n_283), .Y(n_431) );
AND2x4_ASAP7_75t_L g470 ( .A(n_283), .B(n_412), .Y(n_470) );
AND2x2_ASAP7_75t_L g474 ( .A(n_283), .B(n_357), .Y(n_474) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVxp67_ASAP7_75t_L g459 ( .A(n_284), .Y(n_459) );
NOR2x1_ASAP7_75t_L g488 ( .A(n_285), .B(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g353 ( .A(n_286), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_288), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g461 ( .A(n_289), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_291), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g394 ( .A(n_293), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g436 ( .A(n_293), .B(n_348), .Y(n_436) );
INVx2_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g302 ( .A(n_296), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_296), .B(n_341), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B(n_307), .Y(n_297) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_298), .A2(n_479), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2x1_ASAP7_75t_SL g299 ( .A(n_300), .B(n_302), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_301), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_301), .B(n_405), .Y(n_434) );
INVx2_ASAP7_75t_L g443 ( .A(n_301), .Y(n_443) );
AND2x4_ASAP7_75t_SL g448 ( .A(n_301), .B(n_390), .Y(n_448) );
NOR2x1_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_305), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g368 ( .A(n_305), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g375 ( .A(n_305), .Y(n_375) );
OR2x2_ASAP7_75t_L g314 ( .A(n_306), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g369 ( .A(n_306), .Y(n_369) );
INVx1_ASAP7_75t_L g446 ( .A(n_306), .Y(n_446) );
AOI21xp33_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_312), .B(n_314), .Y(n_307) );
AOI32xp33_ASAP7_75t_L g437 ( .A1(n_308), .A2(n_405), .A3(n_438), .B1(n_439), .B2(n_444), .Y(n_437) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx3_ASAP7_75t_L g367 ( .A(n_310), .Y(n_367) );
OR2x2_ASAP7_75t_L g320 ( .A(n_311), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g408 ( .A(n_311), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_312), .A2(n_373), .B1(n_376), .B2(n_378), .Y(n_372) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp33_ASAP7_75t_L g435 ( .A(n_314), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
BUFx2_ASAP7_75t_L g424 ( .A(n_315), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_319), .A2(n_353), .B1(n_382), .B2(n_385), .C(n_388), .Y(n_381) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
INVx1_ASAP7_75t_L g390 ( .A(n_321), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_323), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g429 ( .A(n_323), .B(n_351), .Y(n_429) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x6_ASAP7_75t_L g475 ( .A(n_326), .B(n_476), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_338), .C(n_362), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B(n_333), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_331), .A2(n_364), .B1(n_464), .B2(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx2_ASAP7_75t_L g477 ( .A(n_336), .Y(n_477) );
OR2x2_ASAP7_75t_L g347 ( .A(n_337), .B(n_348), .Y(n_347) );
NOR2x1_ASAP7_75t_SL g387 ( .A(n_337), .B(n_348), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_346), .B2(n_352), .C(n_354), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g352 ( .A(n_341), .B(n_353), .Y(n_352) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g491 ( .A(n_344), .B(n_350), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx1_ASAP7_75t_L g452 ( .A(n_350), .Y(n_452) );
AND2x2_ASAP7_75t_L g403 ( .A(n_351), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g438 ( .A(n_351), .B(n_427), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B(n_359), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_355), .A2(n_473), .B1(n_475), .B2(n_477), .Y(n_472) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_356), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g432 ( .A(n_358), .Y(n_432) );
OR2x2_ASAP7_75t_L g464 ( .A(n_358), .B(n_431), .Y(n_464) );
INVx4_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI321xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .A3(n_366), .B1(n_368), .B2(n_370), .C(n_372), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_SL g384 ( .A(n_374), .Y(n_384) );
AND2x4_ASAP7_75t_L g426 ( .A(n_374), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_374), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx4_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND5x1_ASAP7_75t_L g380 ( .A(n_381), .B(n_400), .C(n_425), .D(n_437), .E(n_447), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_383), .A2(n_414), .B1(n_417), .B2(n_422), .Y(n_413) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI32xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .A3(n_393), .B1(n_394), .B2(n_397), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g468 ( .A(n_398), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_413), .Y(n_400) );
OAI32xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .A3(n_406), .B1(n_409), .B2(n_411), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g476 ( .A(n_404), .Y(n_476) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_409), .A2(n_421), .B(n_468), .C(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVxp33_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_412), .B(n_443), .Y(n_454) );
AND2x2_ASAP7_75t_L g460 ( .A(n_412), .B(n_431), .Y(n_460) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx4_ASAP7_75t_L g419 ( .A(n_416), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_418), .A2(n_426), .A3(n_428), .B1(n_429), .B2(n_430), .C1(n_433), .C2(n_435), .Y(n_425) );
INVx6_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g465 ( .A(n_426), .Y(n_465) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g451 ( .A(n_431), .Y(n_451) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_438), .A2(n_448), .B1(n_449), .B2(n_453), .Y(n_447) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g487 ( .A(n_440), .Y(n_487) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI31xp33_ASAP7_75t_L g486 ( .A1(n_448), .A2(n_487), .A3(n_488), .B(n_490), .Y(n_486) );
INVx2_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
AND4x1_ASAP7_75t_L g455 ( .A(n_456), .B(n_466), .C(n_478), .D(n_486), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_460), .B(n_461), .C(n_463), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_SL g466 ( .A(n_467), .B(n_472), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_546), .B1(n_714), .B2(n_718), .C(n_719), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_509), .B1(n_538), .B2(n_544), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_494), .A2(n_544), .B1(n_716), .B2(n_717), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_501), .B2(n_508), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g508 ( .A(n_501), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B1(n_504), .B2(n_507), .Y(n_501) );
INVx1_ASAP7_75t_L g507 ( .A(n_502), .Y(n_507) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx5_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx5_ASAP7_75t_L g716 ( .A(n_512), .Y(n_716) );
AND2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_529), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .Y(n_513) );
INVxp67_ASAP7_75t_L g542 ( .A(n_514), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g725 ( .A(n_515), .Y(n_725) );
INVx1_ASAP7_75t_L g732 ( .A(n_516), .Y(n_732) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g724 ( .A(n_517), .Y(n_724) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_519), .B(n_533), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .C(n_524), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
CKINVDCx11_ASAP7_75t_R g531 ( .A(n_521), .Y(n_531) );
AND2x4_ASAP7_75t_L g534 ( .A(n_522), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g636 ( .A(n_523), .B(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_523), .Y(n_649) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g537 ( .A(n_526), .B(n_527), .Y(n_537) );
OR2x6_ASAP7_75t_L g659 ( .A(n_526), .B(n_528), .Y(n_659) );
INVx1_ASAP7_75t_L g695 ( .A(n_526), .Y(n_695) );
AND2x4_ASAP7_75t_L g713 ( .A(n_526), .B(n_694), .Y(n_713) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g694 ( .A(n_528), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g633 ( .A(n_537), .B(n_634), .Y(n_633) );
CKINVDCx14_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx3_ASAP7_75t_L g717 ( .A(n_540), .Y(n_717) );
INVx4_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g718 ( .A(n_546), .Y(n_718) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI211x1_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_623), .B(n_628), .C(n_667), .Y(n_547) );
NAND4xp25_ASAP7_75t_SL g548 ( .A(n_549), .B(n_576), .C(n_591), .D(n_608), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_562), .B(n_572), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx3_ASAP7_75t_L g596 ( .A(n_553), .Y(n_596) );
BUFx4f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g611 ( .A(n_554), .Y(n_611) );
INVx2_ASAP7_75t_L g560 ( .A(n_555), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_555), .B(n_561), .Y(n_565) );
INVx2_ASAP7_75t_L g571 ( .A(n_555), .Y(n_571) );
INVx4_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx4_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_558), .Y(n_598) );
INVx4_ASAP7_75t_L g614 ( .A(n_558), .Y(n_614) );
INVx5_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g604 ( .A(n_560), .Y(n_604) );
INVx2_ASAP7_75t_L g570 ( .A(n_561), .Y(n_570) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g579 ( .A(n_564), .Y(n_579) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx12f_ASAP7_75t_L g594 ( .A(n_569), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g590 ( .A(n_570), .Y(n_590) );
AND2x4_ASAP7_75t_L g620 ( .A(n_570), .B(n_571), .Y(n_620) );
BUFx3_ASAP7_75t_L g586 ( .A(n_571), .Y(n_586) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g622 ( .A(n_575), .B(n_607), .Y(n_622) );
AOI21xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_580), .B(n_583), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g585 ( .A(n_582), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g588 ( .A(n_582), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI211xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_595), .C(n_599), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_592), .A2(n_647), .B1(n_650), .B2(n_651), .Y(n_646) );
BUFx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx5_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g617 ( .A(n_602), .Y(n_617) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
BUFx4_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B1(n_613), .B2(n_615), .C(n_616), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_612), .A2(n_686), .B1(n_687), .B2(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g709 ( .A1(n_615), .A2(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx4_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x6_ASAP7_75t_L g692 ( .A(n_626), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g634 ( .A(n_627), .Y(n_634) );
OR2x2_ASAP7_75t_L g658 ( .A(n_627), .B(n_659), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_646), .C(n_655), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_638), .B(n_639), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x4_ASAP7_75t_L g639 ( .A(n_633), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g647 ( .A(n_633), .B(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g651 ( .A(n_633), .B(n_652), .Y(n_651) );
AND2x6_ASAP7_75t_L g712 ( .A(n_634), .B(n_713), .Y(n_712) );
OR2x6_ASAP7_75t_L g657 ( .A(n_635), .B(n_658), .Y(n_657) );
INVx8_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g654 ( .A(n_637), .Y(n_654) );
AND2x4_ASAP7_75t_L g674 ( .A(n_637), .B(n_642), .Y(n_674) );
INVx2_ASAP7_75t_L g698 ( .A(n_640), .Y(n_698) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_641), .Y(n_678) );
AND2x4_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g665 ( .A(n_643), .B(n_644), .Y(n_665) );
AND2x2_ASAP7_75t_L g684 ( .A(n_643), .B(n_645), .Y(n_684) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g666 ( .A(n_658), .Y(n_666) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx5_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g690 ( .A(n_664), .Y(n_690) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_665), .Y(n_706) );
AND2x4_ASAP7_75t_L g670 ( .A(n_666), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g676 ( .A(n_666), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_679), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_675), .B2(n_676), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_674), .Y(n_688) );
INVx4_ASAP7_75t_L g703 ( .A(n_674), .Y(n_703) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_696), .B1(n_699), .B2(n_707), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx4f_ASAP7_75t_L g711 ( .A(n_683), .Y(n_711) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g708 ( .A(n_698), .Y(n_708) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx3_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_726), .B1(n_729), .B2(n_730), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g731 ( .A(n_725), .B(n_732), .Y(n_731) );
INVxp33_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
endmodule