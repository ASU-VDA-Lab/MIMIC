module fake_jpeg_3393_n_101 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_0),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_32),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_20),
.Y(n_26)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_2),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_18),
.A2(n_0),
.B(n_7),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_8),
.Y(n_41)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_40),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_22),
.B1(n_17),
.B2(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_45),
.B1(n_50),
.B2(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_17),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_21),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_21),
.B1(n_12),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_23),
.B1(n_13),
.B2(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_48),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_59),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_27),
.B1(n_21),
.B2(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_47),
.B1(n_38),
.B2(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_10),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_39),
.B1(n_38),
.B2(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_40),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_44),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_71),
.B1(n_63),
.B2(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_53),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_74),
.A2(n_79),
.B1(n_68),
.B2(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_66),
.B(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

AOI322xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_42),
.A3(n_43),
.B1(n_54),
.B2(n_62),
.C1(n_65),
.C2(n_73),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_81),
.C(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_87),
.C(n_77),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_75),
.C(n_74),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_85),
.CI(n_86),
.CON(n_93),
.SN(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_94),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_92),
.C(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_97),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_93),
.Y(n_101)
);


endmodule