module fake_netlist_6_515_n_1896 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1896);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1896;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1669;
wire n_1403;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx3_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_178),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_6),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_45),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_15),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_173),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_5),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_14),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_3),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_24),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_1),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_112),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_96),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_68),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_35),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_62),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_76),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_75),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_113),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_73),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_114),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_62),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_43),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_74),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_134),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_18),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_79),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_45),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_141),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_138),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_43),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_102),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_111),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_67),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_28),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_127),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_49),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_90),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_23),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_84),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_166),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_27),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_103),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_20),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_32),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_9),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_163),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_58),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_87),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_85),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_118),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_64),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_107),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_93),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_157),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_37),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_1),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_176),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_56),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_51),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_94),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_165),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_133),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_158),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_146),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_81),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_40),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_50),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_142),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_71),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_91),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_137),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_50),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_97),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_123),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_57),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_15),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_29),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_162),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_54),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_106),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_52),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_144),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_149),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_23),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_59),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_21),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_117),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_24),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_77),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_110),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_30),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_88),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_13),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_22),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_17),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_70),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_108),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_95),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_168),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_109),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_21),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_28),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_92),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_5),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_57),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_169),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_78),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_52),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_65),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_151),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_172),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_125),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_152),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_14),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_154),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_89),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_29),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_46),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_116),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_69),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_13),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_129),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_40),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_55),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_61),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_32),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_60),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_56),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_30),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_9),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_0),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_101),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_27),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_44),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_31),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_160),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_82),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_51),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_83),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_55),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_53),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_48),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_26),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_39),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_2),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_60),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_100),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_47),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_31),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_72),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_122),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_35),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_11),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_131),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_53),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_98),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_0),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_209),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_209),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_184),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_189),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_209),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_278),
.B(n_320),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_197),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_199),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_258),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_198),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_198),
.B(n_2),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_252),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_209),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_239),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_209),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_252),
.B(n_4),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_259),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_259),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_200),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_203),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_207),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_212),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_216),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_180),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_270),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_180),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_226),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_264),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_260),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_219),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_186),
.B(n_192),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_220),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_259),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_259),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_222),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_206),
.B(n_4),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_182),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_230),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_259),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_208),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_183),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_226),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_231),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_208),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_232),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_192),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_237),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_238),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_283),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_240),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_283),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_286),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_244),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_226),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_286),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_190),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_193),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_185),
.B(n_6),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_193),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_260),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_185),
.B(n_7),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_202),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_202),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_217),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_217),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_221),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_221),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_330),
.B(n_7),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_241),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_206),
.B(n_8),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_241),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_275),
.B(n_8),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_274),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_274),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_277),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_277),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_281),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_293),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_293),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_246),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_297),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_297),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_306),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_247),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_275),
.B(n_10),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_248),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_269),
.B(n_10),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_362),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_376),
.B(n_181),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_360),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_361),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_364),
.B(n_309),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_373),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_363),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_375),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_377),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_366),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_377),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_378),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_400),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_368),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_365),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_397),
.B(n_309),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_431),
.B(n_312),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_403),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_385),
.B(n_387),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_312),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_371),
.B(n_187),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_420),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_403),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_415),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_415),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_421),
.B(n_349),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_370),
.B(n_349),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_369),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_380),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_381),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_415),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_423),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_401),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_382),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_R g502 ( 
.A(n_383),
.B(n_250),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_384),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_R g505 ( 
.A(n_393),
.B(n_253),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_399),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_386),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_404),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_408),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_SL g511 ( 
.A(n_433),
.B(n_330),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_414),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_423),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_419),
.B(n_254),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_422),
.B(n_262),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_R g516 ( 
.A(n_374),
.B(n_359),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_396),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_406),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_409),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_429),
.B(n_187),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_411),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_441),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_372),
.B(n_188),
.Y(n_524)
);

BUFx8_ASAP7_75t_L g525 ( 
.A(n_392),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_424),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_481),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_470),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

NAND3xp33_ASAP7_75t_L g531 ( 
.A(n_451),
.B(n_402),
.C(n_398),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_477),
.A2(n_479),
.B1(n_451),
.B2(n_486),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_525),
.B(n_486),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_455),
.B(n_191),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_484),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_226),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_470),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_484),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_482),
.B(n_205),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_475),
.A2(n_447),
.B1(n_445),
.B2(n_389),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_485),
.B(n_367),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_485),
.B(n_379),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_455),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_487),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_487),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_525),
.B(n_446),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_525),
.B(n_191),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_476),
.Y(n_549)
);

AND3x2_ASAP7_75t_L g550 ( 
.A(n_475),
.B(n_211),
.C(n_204),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_525),
.B(n_482),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_476),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_477),
.B(n_263),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_477),
.B(n_265),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_477),
.B(n_266),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_495),
.B(n_188),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_502),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_477),
.A2(n_346),
.B1(n_214),
.B2(n_201),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_450),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_498),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_525),
.B(n_204),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_470),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_493),
.A2(n_417),
.B1(n_187),
.B2(n_276),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_498),
.Y(n_565)
);

AND2x6_ASAP7_75t_L g566 ( 
.A(n_479),
.B(n_211),
.Y(n_566)
);

BUFx4f_ASAP7_75t_L g567 ( 
.A(n_479),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_479),
.B(n_514),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_479),
.B(n_515),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_515),
.B(n_267),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_483),
.B(n_272),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_455),
.B(n_213),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_L g573 ( 
.A(n_493),
.B(n_430),
.C(n_407),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_470),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_499),
.Y(n_575)
);

NOR2x1p5_ASAP7_75t_L g576 ( 
.A(n_495),
.B(n_201),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_520),
.B(n_434),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_520),
.A2(n_288),
.B1(n_325),
.B2(n_323),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_499),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_502),
.Y(n_580)
);

BUFx4f_ASAP7_75t_L g581 ( 
.A(n_524),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_455),
.B(n_213),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_455),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_483),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_483),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_492),
.B(n_215),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_513),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_492),
.B(n_424),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_493),
.B(n_392),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_513),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_527),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_524),
.B(n_215),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_524),
.B(n_346),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_495),
.B(n_425),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_449),
.B(n_285),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_504),
.B(n_425),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_527),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_516),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_504),
.B(n_218),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_488),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_504),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_511),
.B(n_210),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_459),
.B(n_426),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_478),
.Y(n_605)
);

BUFx6f_ASAP7_75t_SL g606 ( 
.A(n_517),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_511),
.B(n_426),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_449),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_452),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_505),
.B(n_463),
.Y(n_610)
);

CKINVDCx16_ASAP7_75t_R g611 ( 
.A(n_494),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_516),
.A2(n_496),
.B1(n_501),
.B2(n_474),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_503),
.B(n_427),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_505),
.B(n_218),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_500),
.A2(n_214),
.B1(n_327),
.B2(n_332),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_507),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_452),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_453),
.B(n_291),
.Y(n_618)
);

AND2x6_ASAP7_75t_L g619 ( 
.A(n_488),
.B(n_223),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_509),
.A2(n_287),
.B1(n_319),
.B2(n_310),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_478),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_510),
.B(n_223),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_512),
.B(n_427),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_480),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_453),
.B(n_428),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_488),
.B(n_224),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_454),
.B(n_292),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_488),
.B(n_224),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_480),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_454),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_456),
.B(n_298),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_518),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_488),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_519),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_489),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_489),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_456),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_489),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_458),
.Y(n_640)
);

AND2x2_ASAP7_75t_SL g641 ( 
.A(n_506),
.B(n_225),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_458),
.B(n_428),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_460),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_489),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_523),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_494),
.Y(n_646)
);

AND2x6_ASAP7_75t_L g647 ( 
.A(n_480),
.B(n_225),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_460),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_521),
.B(n_432),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_461),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_500),
.A2(n_316),
.B1(n_306),
.B2(n_326),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_461),
.B(n_300),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_489),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_491),
.Y(n_654)
);

AO22x2_ASAP7_75t_L g655 ( 
.A1(n_462),
.A2(n_332),
.B1(n_342),
.B2(n_344),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_462),
.B(n_302),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_523),
.B(n_227),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_SL g658 ( 
.A1(n_464),
.A2(n_228),
.B(n_227),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_526),
.B(n_435),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_464),
.B(n_308),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_523),
.B(n_228),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_466),
.B(n_313),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_466),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_467),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_490),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_523),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_467),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_490),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_490),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_506),
.B(n_435),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_468),
.B(n_436),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_490),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_491),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_549),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_R g675 ( 
.A(n_633),
.B(n_522),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_585),
.B(n_448),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_544),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_584),
.B(n_194),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_549),
.Y(n_679)
);

O2A1O1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_593),
.A2(n_342),
.B(n_326),
.C(n_327),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_584),
.B(n_195),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_544),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_583),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_532),
.B(n_490),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_604),
.B(n_196),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_583),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_528),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_552),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_568),
.B(n_569),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_590),
.A2(n_344),
.B1(n_316),
.B2(n_354),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_612),
.B(n_448),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_604),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_581),
.B(n_226),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_613),
.B(n_229),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_602),
.B(n_354),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_649),
.B(n_436),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g697 ( 
.A(n_541),
.B(n_236),
.C(n_234),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_570),
.B(n_468),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_581),
.A2(n_317),
.B1(n_339),
.B2(n_341),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_590),
.A2(n_358),
.B1(n_338),
.B2(n_321),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_530),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_589),
.B(n_437),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_595),
.B(n_469),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_577),
.A2(n_315),
.B1(n_353),
.B2(n_356),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_535),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_567),
.B(n_226),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_595),
.B(n_469),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_597),
.B(n_472),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_597),
.B(n_472),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_613),
.B(n_242),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_567),
.B(n_226),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_653),
.B(n_491),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_600),
.B(n_226),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_594),
.A2(n_334),
.B(n_251),
.C(n_324),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_577),
.B(n_497),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_638),
.B(n_497),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_558),
.B(n_251),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_638),
.B(n_497),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_580),
.B(n_255),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_555),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_640),
.B(n_500),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_555),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_640),
.B(n_500),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_539),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_545),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_560),
.B(n_508),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_546),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_624),
.B(n_438),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_624),
.B(n_226),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_561),
.B(n_500),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_565),
.B(n_523),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_540),
.B(n_233),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_533),
.A2(n_314),
.B1(n_318),
.B2(n_322),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_537),
.A2(n_271),
.B1(n_324),
.B2(n_311),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_636),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_639),
.B(n_235),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_575),
.B(n_579),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_587),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_588),
.B(n_523),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_587),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_591),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_605),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_557),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_639),
.B(n_294),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_639),
.B(n_255),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_665),
.B(n_271),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_L g748 ( 
.A(n_621),
.B(n_256),
.C(n_257),
.Y(n_748)
);

AND2x2_ASAP7_75t_SL g749 ( 
.A(n_537),
.B(n_273),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_605),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_542),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_641),
.A2(n_273),
.B1(n_311),
.B2(n_305),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_622),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_641),
.A2(n_280),
.B1(n_334),
.B2(n_305),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_533),
.A2(n_289),
.B1(n_280),
.B2(n_282),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_665),
.B(n_282),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_592),
.B(n_598),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_571),
.B(n_523),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_608),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_599),
.B(n_506),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_531),
.B(n_345),
.C(n_243),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_609),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_553),
.A2(n_284),
.B1(n_289),
.B2(n_299),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_623),
.B(n_245),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_622),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_646),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_625),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_534),
.B(n_299),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_617),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_534),
.B(n_301),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_631),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_543),
.B(n_438),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_551),
.A2(n_301),
.B1(n_352),
.B2(n_276),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_607),
.A2(n_352),
.B1(n_261),
.B2(n_268),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_593),
.A2(n_440),
.B1(n_444),
.B2(n_442),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_625),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_594),
.A2(n_348),
.B1(n_279),
.B2(n_290),
.C(n_295),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_630),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_643),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_L g781 ( 
.A(n_564),
.B(n_351),
.C(n_296),
.Y(n_781)
);

NOR3x1_ASAP7_75t_L g782 ( 
.A(n_573),
.B(n_444),
.C(n_442),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_554),
.A2(n_350),
.B1(n_303),
.B2(n_304),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_616),
.B(n_439),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_534),
.B(n_526),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_630),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_572),
.B(n_439),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_572),
.B(n_457),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_648),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_572),
.B(n_457),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_654),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_582),
.B(n_457),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_665),
.B(n_187),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_654),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_556),
.A2(n_465),
.B(n_473),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_623),
.B(n_307),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_672),
.B(n_249),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_576),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_SL g799 ( 
.A1(n_611),
.A2(n_508),
.B1(n_343),
.B2(n_340),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_559),
.B(n_355),
.C(n_328),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_650),
.B(n_443),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_663),
.B(n_473),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_619),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_616),
.B(n_443),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_664),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_616),
.B(n_440),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_667),
.B(n_473),
.Y(n_807)
);

NAND2x1_ASAP7_75t_L g808 ( 
.A(n_672),
.B(n_471),
.Y(n_808)
);

BUFx5_ASAP7_75t_L g809 ( 
.A(n_619),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_636),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_586),
.B(n_335),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_586),
.B(n_336),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_637),
.B(n_249),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_637),
.B(n_471),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_637),
.B(n_347),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_603),
.B(n_331),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_614),
.B(n_333),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_644),
.B(n_357),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_596),
.B(n_337),
.Y(n_819)
);

NAND2x1_ASAP7_75t_L g820 ( 
.A(n_644),
.B(n_416),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_644),
.B(n_413),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_618),
.B(n_628),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_668),
.B(n_412),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_668),
.B(n_276),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_659),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_632),
.B(n_276),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_551),
.A2(n_249),
.B1(n_410),
.B2(n_177),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_610),
.B(n_410),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_658),
.A2(n_249),
.B(n_12),
.C(n_16),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_668),
.B(n_171),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_669),
.B(n_161),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_652),
.B(n_11),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_669),
.B(n_153),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_578),
.B(n_12),
.C(n_16),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_656),
.B(n_19),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_687),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_677),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_677),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_677),
.Y(n_839)
);

CKINVDCx8_ASAP7_75t_R g840 ( 
.A(n_718),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_689),
.A2(n_660),
.B(n_662),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_684),
.A2(n_536),
.B(n_601),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_736),
.Y(n_843)
);

O2A1O1Ixp5_ASAP7_75t_L g844 ( 
.A1(n_706),
.A2(n_548),
.B(n_562),
.C(n_547),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_822),
.B(n_600),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_692),
.A2(n_547),
.B1(n_562),
.B2(n_548),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_758),
.A2(n_536),
.B(n_601),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_766),
.B(n_633),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_785),
.A2(n_536),
.B(n_601),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_822),
.B(n_600),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_736),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_752),
.A2(n_754),
.B1(n_755),
.B2(n_682),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_729),
.B(n_600),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_701),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_716),
.A2(n_634),
.B(n_620),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_705),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_685),
.B(n_635),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_804),
.B(n_635),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_776),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_722),
.A2(n_634),
.B(n_563),
.Y(n_860)
);

NAND2xp33_ASAP7_75t_L g861 ( 
.A(n_752),
.B(n_566),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_808),
.A2(n_661),
.B(n_657),
.Y(n_862)
);

O2A1O1Ixp5_ASAP7_75t_L g863 ( 
.A1(n_706),
.A2(n_661),
.B(n_657),
.C(n_563),
.Y(n_863)
);

AOI21x1_ASAP7_75t_L g864 ( 
.A1(n_693),
.A2(n_673),
.B(n_670),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_806),
.B(n_550),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_787),
.B(n_566),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_725),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_772),
.Y(n_868)
);

OAI21xp33_ASAP7_75t_L g869 ( 
.A1(n_694),
.A2(n_615),
.B(n_651),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_694),
.B(n_606),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_SL g871 ( 
.A(n_710),
.B(n_671),
.C(n_642),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_795),
.A2(n_673),
.B(n_626),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_787),
.B(n_801),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_710),
.B(n_566),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_712),
.A2(n_529),
.B(n_538),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_788),
.A2(n_529),
.B(n_538),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_760),
.B(n_642),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_698),
.B(n_626),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_790),
.A2(n_529),
.B(n_538),
.Y(n_879)
);

AO21x1_ASAP7_75t_L g880 ( 
.A1(n_730),
.A2(n_655),
.B(n_647),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_819),
.B(n_574),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_819),
.B(n_574),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_792),
.A2(n_574),
.B(n_645),
.Y(n_883)
);

BUFx12f_ASAP7_75t_L g884 ( 
.A(n_744),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_SL g885 ( 
.A(n_727),
.B(n_606),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_677),
.B(n_574),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_801),
.B(n_645),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_703),
.B(n_655),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_798),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_826),
.A2(n_629),
.B1(n_627),
.B2(n_619),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_707),
.B(n_647),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_708),
.B(n_647),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_709),
.B(n_645),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_751),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_717),
.A2(n_645),
.B(n_666),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_816),
.B(n_19),
.Y(n_896)
);

BUFx12f_ASAP7_75t_L g897 ( 
.A(n_696),
.Y(n_897)
);

NOR2x1_ASAP7_75t_L g898 ( 
.A(n_834),
.B(n_629),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_724),
.A2(n_666),
.B(n_629),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_726),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_702),
.B(n_627),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_693),
.A2(n_666),
.B(n_627),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_754),
.A2(n_666),
.B1(n_627),
.B2(n_619),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_828),
.B(n_627),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_825),
.B(n_20),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_719),
.A2(n_150),
.B(n_147),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_810),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_734),
.B(n_139),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_676),
.B(n_25),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_728),
.B(n_99),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_711),
.A2(n_136),
.B(n_132),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_682),
.A2(n_128),
.B1(n_126),
.B2(n_119),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_683),
.A2(n_115),
.B1(n_86),
.B2(n_80),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_683),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_742),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_810),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_764),
.A2(n_25),
.B(n_26),
.C(n_33),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_695),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_711),
.A2(n_66),
.B(n_34),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_731),
.A2(n_33),
.B(n_34),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_732),
.A2(n_36),
.B(n_37),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_816),
.B(n_678),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_740),
.A2(n_36),
.B(n_38),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_811),
.B(n_812),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_686),
.A2(n_63),
.B1(n_39),
.B2(n_41),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_814),
.A2(n_38),
.B(n_41),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_764),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_927)
);

INVx11_ASAP7_75t_L g928 ( 
.A(n_675),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_811),
.B(n_42),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_675),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_759),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_674),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_796),
.A2(n_63),
.B(n_48),
.C(n_49),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_695),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_812),
.B(n_47),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_762),
.B(n_54),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_738),
.A2(n_58),
.B(n_61),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_769),
.B(n_771),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_718),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_774),
.A2(n_733),
.B(n_715),
.C(n_730),
.Y(n_940)
);

OAI21xp33_ASAP7_75t_L g941 ( 
.A1(n_796),
.A2(n_778),
.B(n_690),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_817),
.B(n_686),
.Y(n_942)
);

NOR2x1p5_ASAP7_75t_SL g943 ( 
.A(n_809),
.B(n_679),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_757),
.A2(n_756),
.B(n_746),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_774),
.A2(n_733),
.B(n_715),
.C(n_829),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_749),
.A2(n_746),
.B(n_747),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_747),
.A2(n_756),
.B(n_815),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_695),
.B(n_678),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_780),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_789),
.B(n_805),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_681),
.B(n_718),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_817),
.B(n_681),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_832),
.B(n_835),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_818),
.A2(n_745),
.B(n_737),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_821),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_832),
.B(n_835),
.Y(n_956)
);

INVxp67_ASAP7_75t_L g957 ( 
.A(n_720),
.Y(n_957)
);

BUFx4f_ASAP7_75t_L g958 ( 
.A(n_720),
.Y(n_958)
);

NAND2x1p5_ASAP7_75t_L g959 ( 
.A(n_803),
.B(n_830),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_813),
.A2(n_824),
.B1(n_749),
.B2(n_773),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_782),
.B(n_720),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_737),
.A2(n_745),
.B(n_807),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_688),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_802),
.A2(n_768),
.B(n_770),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_735),
.B(n_690),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_735),
.A2(n_827),
.B1(n_793),
.B2(n_797),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_700),
.B(n_823),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_713),
.B(n_779),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_697),
.B(n_761),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_793),
.A2(n_797),
.B(n_714),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_L g971 ( 
.A(n_748),
.B(n_781),
.C(n_704),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_699),
.B(n_691),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_721),
.B(n_791),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_723),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_831),
.A2(n_833),
.B(n_824),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_813),
.A2(n_786),
.B(n_739),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_783),
.B(n_799),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_741),
.B(n_777),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_803),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_743),
.B(n_794),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_680),
.A2(n_763),
.B(n_800),
.C(n_820),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_750),
.B(n_753),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_765),
.A2(n_767),
.B(n_830),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_775),
.B(n_829),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_775),
.B(n_803),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_809),
.B(n_689),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_809),
.A2(n_689),
.B(n_684),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_809),
.A2(n_689),
.B(n_684),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_809),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_689),
.B(n_822),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_822),
.A2(n_694),
.B(n_710),
.C(n_685),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_822),
.A2(n_694),
.B1(n_710),
.B2(n_685),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_689),
.B(n_822),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_677),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_R g995 ( 
.A(n_727),
.B(n_633),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_689),
.B(n_822),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_689),
.A2(n_684),
.B(n_567),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_687),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_736),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_689),
.B(n_822),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_689),
.A2(n_684),
.B(n_567),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_692),
.B(n_599),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_729),
.B(n_784),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_685),
.B(n_710),
.C(n_694),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_677),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_736),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_689),
.A2(n_684),
.B(n_567),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_784),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_729),
.B(n_784),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_689),
.A2(n_532),
.B1(n_692),
.B2(n_752),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_677),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_689),
.A2(n_684),
.B(n_569),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_687),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_689),
.A2(n_684),
.B(n_567),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_990),
.A2(n_996),
.B(n_993),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_836),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_979),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_1000),
.A2(n_986),
.B(n_1012),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_992),
.B(n_922),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_942),
.A2(n_882),
.B(n_881),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_842),
.A2(n_987),
.B(n_997),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_842),
.A2(n_872),
.B(n_864),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_987),
.A2(n_983),
.B(n_847),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_983),
.A2(n_847),
.B(n_997),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_861),
.A2(n_1007),
.B(n_1001),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_991),
.A2(n_941),
.B(n_924),
.C(n_896),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_848),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1004),
.A2(n_857),
.B1(n_952),
.B2(n_1003),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_838),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_866),
.B(n_873),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_854),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_SL g1032 ( 
.A1(n_988),
.A2(n_852),
.B(n_850),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1014),
.A2(n_970),
.B(n_845),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_838),
.Y(n_1034)
);

OA22x2_ASAP7_75t_L g1035 ( 
.A1(n_868),
.A2(n_927),
.B1(n_953),
.B2(n_956),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_SL g1036 ( 
.A1(n_929),
.A2(n_935),
.B1(n_945),
.B2(n_888),
.C(n_1010),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_884),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_SL g1038 ( 
.A1(n_880),
.A2(n_919),
.B(n_911),
.Y(n_1038)
);

INVx3_ASAP7_75t_SL g1039 ( 
.A(n_930),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_L g1040 ( 
.A(n_977),
.B(n_1009),
.C(n_1002),
.Y(n_1040)
);

AOI21x1_ASAP7_75t_L g1041 ( 
.A1(n_970),
.A2(n_954),
.B(n_947),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_846),
.B(n_960),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_878),
.B(n_877),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_894),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_860),
.A2(n_975),
.B(n_902),
.Y(n_1045)
);

AOI221xp5_ASAP7_75t_SL g1046 ( 
.A1(n_869),
.A2(n_905),
.B1(n_917),
.B2(n_933),
.C(n_936),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_965),
.A2(n_940),
.B(n_984),
.C(n_946),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_944),
.A2(n_841),
.B(n_863),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_SL g1049 ( 
.A(n_961),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_897),
.B(n_1008),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_853),
.B(n_874),
.Y(n_1051)
);

OA21x2_ASAP7_75t_L g1052 ( 
.A1(n_855),
.A2(n_975),
.B(n_844),
.Y(n_1052)
);

INVx3_ASAP7_75t_SL g1053 ( 
.A(n_909),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_865),
.B(n_858),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_995),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_944),
.A2(n_841),
.B(n_964),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_889),
.Y(n_1057)
);

AO31x2_ASAP7_75t_L g1058 ( 
.A1(n_966),
.A2(n_947),
.A3(n_962),
.B(n_954),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_856),
.Y(n_1059)
);

AOI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_971),
.A2(n_951),
.B(n_870),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_962),
.A2(n_964),
.A3(n_891),
.B(n_892),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_932),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_867),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_963),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_849),
.A2(n_976),
.B(n_899),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_899),
.A2(n_862),
.B(n_876),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_974),
.Y(n_1067)
);

BUFx12f_ASAP7_75t_L g1068 ( 
.A(n_939),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_893),
.A2(n_883),
.B(n_886),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_879),
.A2(n_875),
.B(n_959),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_904),
.A2(n_901),
.B(n_989),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_838),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_900),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_839),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_955),
.B(n_938),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_915),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_839),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_931),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_948),
.B(n_1013),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_895),
.A2(n_898),
.B(n_906),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_979),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_994),
.B(n_839),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_950),
.B(n_998),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_843),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_851),
.Y(n_1085)
);

BUFx12f_ASAP7_75t_L g1086 ( 
.A(n_961),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_981),
.A2(n_921),
.A3(n_923),
.B(n_926),
.Y(n_1087)
);

INVx4_ASAP7_75t_L g1088 ( 
.A(n_1005),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_949),
.B(n_871),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_1005),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_967),
.A2(n_914),
.B1(n_985),
.B2(n_887),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_937),
.A2(n_919),
.B(n_920),
.C(n_926),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_840),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_SL g1094 ( 
.A(n_979),
.B(n_1005),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_866),
.A2(n_914),
.B(n_887),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_994),
.B(n_837),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_968),
.A2(n_973),
.B(n_978),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_980),
.A2(n_982),
.B(n_903),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_972),
.A2(n_859),
.B(n_1006),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_1011),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_873),
.B(n_918),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_907),
.A2(n_999),
.B(n_916),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_912),
.A2(n_913),
.B(n_923),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_957),
.B(n_934),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_928),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_910),
.A2(n_908),
.B(n_890),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_921),
.A2(n_920),
.B(n_937),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_969),
.B(n_885),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_910),
.A2(n_958),
.B(n_943),
.Y(n_1109)
);

NOR2xp67_ASAP7_75t_L g1110 ( 
.A(n_925),
.B(n_958),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_848),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_990),
.B(n_993),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_897),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_990),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_990),
.B(n_993),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_991),
.A2(n_992),
.B(n_924),
.Y(n_1116)
);

AOI221x1_ASAP7_75t_L g1117 ( 
.A1(n_991),
.A2(n_1004),
.B1(n_956),
.B2(n_953),
.C(n_896),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_990),
.B(n_993),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_848),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_991),
.A2(n_992),
.B(n_924),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_838),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_979),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_842),
.A2(n_872),
.B(n_864),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_990),
.A2(n_689),
.B(n_567),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_992),
.A2(n_990),
.B(n_996),
.C(n_993),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_842),
.A2(n_872),
.B(n_864),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_990),
.B(n_993),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_991),
.A2(n_992),
.B(n_924),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_SL g1129 ( 
.A1(n_880),
.A2(n_919),
.B(n_911),
.Y(n_1129)
);

AOI21xp33_ASAP7_75t_L g1130 ( 
.A1(n_992),
.A2(n_924),
.B(n_991),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_942),
.A2(n_882),
.B(n_881),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_932),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_991),
.A2(n_992),
.B(n_924),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_990),
.B(n_993),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_992),
.B(n_990),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_990),
.B(n_993),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_880),
.A2(n_991),
.A3(n_966),
.B(n_997),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_992),
.B(n_692),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1003),
.B(n_1009),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_868),
.B(n_646),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_990),
.A2(n_689),
.B(n_567),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_836),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_990),
.A2(n_689),
.B(n_567),
.Y(n_1143)
);

NAND2x1_ASAP7_75t_L g1144 ( 
.A(n_994),
.B(n_914),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_897),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_884),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_842),
.A2(n_872),
.B(n_864),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_866),
.B(n_873),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_848),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_842),
.A2(n_872),
.B(n_864),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_897),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_990),
.B(n_993),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_990),
.B(n_993),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_932),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_988),
.A2(n_855),
.B(n_997),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_991),
.A2(n_992),
.B(n_924),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_SL g1157 ( 
.A(n_992),
.B(n_991),
.C(n_857),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1003),
.B(n_1009),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_991),
.A2(n_992),
.B(n_924),
.Y(n_1159)
);

AOI22x1_ASAP7_75t_L g1160 ( 
.A1(n_841),
.A2(n_964),
.B1(n_970),
.B2(n_954),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_836),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_990),
.A2(n_689),
.B(n_567),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_992),
.A2(n_990),
.B1(n_996),
.B2(n_993),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_990),
.B(n_993),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_836),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_992),
.A2(n_990),
.B(n_996),
.C(n_993),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_838),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1017),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1030),
.B(n_1148),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1017),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1019),
.B(n_1027),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1016),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1030),
.B(n_1148),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1017),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1031),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1112),
.B(n_1115),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1111),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1124),
.A2(n_1143),
.B(n_1141),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1119),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1139),
.B(n_1158),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1149),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1118),
.B(n_1127),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1134),
.B(n_1136),
.Y(n_1183)
);

OAI21xp33_ASAP7_75t_L g1184 ( 
.A1(n_1138),
.A2(n_1153),
.B(n_1152),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1138),
.B(n_1054),
.Y(n_1185)
);

INVx3_ASAP7_75t_SL g1186 ( 
.A(n_1105),
.Y(n_1186)
);

CKINVDCx6p67_ASAP7_75t_R g1187 ( 
.A(n_1039),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1081),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1157),
.A2(n_1108),
.B1(n_1079),
.B2(n_1028),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_SL g1190 ( 
.A1(n_1026),
.A2(n_1042),
.B(n_1130),
.C(n_1166),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1059),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1164),
.B(n_1163),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1081),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1063),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1073),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1108),
.A2(n_1060),
.B1(n_1040),
.B2(n_1135),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1026),
.A2(n_1042),
.B(n_1116),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1056),
.A2(n_1162),
.B(n_1133),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1076),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1120),
.A2(n_1128),
.B(n_1156),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1068),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1125),
.B(n_1166),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1030),
.B(n_1148),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1101),
.B(n_1053),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1078),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1125),
.B(n_1015),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1135),
.B(n_1114),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1053),
.B(n_1104),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_1081),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1043),
.B(n_1159),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1018),
.A2(n_1032),
.B(n_1033),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1025),
.A2(n_1048),
.B(n_1106),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1051),
.A2(n_1047),
.B(n_1160),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1055),
.B(n_1039),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1081),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1047),
.A2(n_1155),
.B(n_1024),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1142),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1140),
.B(n_1075),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1110),
.B(n_1057),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1161),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1165),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1044),
.B(n_1083),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1035),
.A2(n_1089),
.B1(n_1049),
.B2(n_1086),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1050),
.B(n_1109),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1062),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1105),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1117),
.B(n_1036),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1050),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1050),
.Y(n_1229)
);

CKINVDCx14_ASAP7_75t_R g1230 ( 
.A(n_1113),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1068),
.Y(n_1231)
);

INVx5_ASAP7_75t_L g1232 ( 
.A(n_1122),
.Y(n_1232)
);

OR2x6_ASAP7_75t_L g1233 ( 
.A(n_1086),
.B(n_1095),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1122),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1145),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1046),
.B(n_1064),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1035),
.B(n_1064),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1067),
.B(n_1132),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1093),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1155),
.A2(n_1071),
.B(n_1097),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1067),
.Y(n_1241)
);

CKINVDCx16_ASAP7_75t_R g1242 ( 
.A(n_1093),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1049),
.B(n_1091),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_SL g1244 ( 
.A(n_1037),
.B(n_1146),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1088),
.B(n_1121),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1132),
.B(n_1154),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1084),
.B(n_1085),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1052),
.A2(n_1092),
.B(n_1023),
.Y(n_1248)
);

AOI221x1_ASAP7_75t_L g1249 ( 
.A1(n_1038),
.A2(n_1129),
.B1(n_1099),
.B2(n_1102),
.C(n_1137),
.Y(n_1249)
);

OAI321xp33_ASAP7_75t_L g1250 ( 
.A1(n_1041),
.A2(n_1021),
.A3(n_1020),
.B1(n_1131),
.B2(n_1069),
.C(n_1085),
.Y(n_1250)
);

INVx8_ASAP7_75t_L g1251 ( 
.A(n_1122),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1151),
.B(n_1121),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1100),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1137),
.B(n_1100),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1122),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1037),
.Y(n_1256)
);

AOI21xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1167),
.A2(n_1090),
.B(n_1082),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1137),
.B(n_1061),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1088),
.B(n_1029),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1137),
.B(n_1061),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1146),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1061),
.B(n_1087),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1029),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1061),
.B(n_1087),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1088),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1090),
.B(n_1167),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1034),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1034),
.B(n_1074),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1072),
.B(n_1077),
.Y(n_1269)
);

OAI21xp33_ASAP7_75t_L g1270 ( 
.A1(n_1107),
.A2(n_1103),
.B(n_1082),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1087),
.B(n_1077),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1072),
.B(n_1074),
.Y(n_1272)
);

BUFx12f_ASAP7_75t_L g1273 ( 
.A(n_1096),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1144),
.B(n_1096),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1107),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1087),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1094),
.B(n_1058),
.Y(n_1277)
);

CKINVDCx8_ASAP7_75t_R g1278 ( 
.A(n_1058),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1058),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1098),
.B(n_1080),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1022),
.A2(n_1123),
.B(n_1150),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1080),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1103),
.B(n_1070),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1022),
.B(n_1126),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1065),
.B(n_1045),
.Y(n_1285)
);

INVx5_ASAP7_75t_L g1286 ( 
.A(n_1066),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1066),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1147),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1138),
.B(n_692),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1112),
.B(n_990),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1044),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1068),
.Y(n_1292)
);

BUFx10_ASAP7_75t_L g1293 ( 
.A(n_1108),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1016),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1016),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1016),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1112),
.A2(n_992),
.B1(n_993),
.B2(n_990),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1111),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1016),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1124),
.A2(n_993),
.B(n_990),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_SL g1301 ( 
.A1(n_1109),
.A2(n_880),
.B(n_1106),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1057),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1112),
.B(n_990),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1139),
.B(n_1158),
.Y(n_1304)
);

NOR2x1_ASAP7_75t_SL g1305 ( 
.A(n_1091),
.B(n_838),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1016),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1028),
.B(n_992),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1017),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1042),
.A2(n_993),
.B(n_990),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1111),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1157),
.A2(n_1004),
.B1(n_941),
.B2(n_992),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1016),
.Y(n_1312)
);

NAND2x1_ASAP7_75t_L g1313 ( 
.A(n_1088),
.B(n_994),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1112),
.B(n_990),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1016),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1030),
.B(n_1148),
.Y(n_1316)
);

OR2x6_ASAP7_75t_L g1317 ( 
.A(n_1109),
.B(n_1050),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1177),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1307),
.A2(n_1311),
.B1(n_1200),
.B2(n_1289),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1243),
.A2(n_1184),
.B1(n_1189),
.B2(n_1196),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1176),
.A2(n_1182),
.B1(n_1183),
.B2(n_1314),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1239),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1186),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1271),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1176),
.B(n_1182),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_SL g1326 ( 
.A1(n_1301),
.A2(n_1305),
.B(n_1309),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1183),
.B(n_1290),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1191),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1185),
.B(n_1180),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1291),
.Y(n_1330)
);

AO21x1_ASAP7_75t_L g1331 ( 
.A1(n_1197),
.A2(n_1227),
.B(n_1202),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1194),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1290),
.B(n_1303),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1199),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_R g1335 ( 
.A1(n_1171),
.A2(n_1218),
.B1(n_1296),
.B2(n_1295),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1205),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1179),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1223),
.A2(n_1297),
.B(n_1192),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1237),
.B(n_1303),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1304),
.B(n_1293),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1220),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1181),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1314),
.B(n_1297),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1293),
.A2(n_1192),
.B1(n_1224),
.B2(n_1210),
.Y(n_1344)
);

BUFx2_ASAP7_75t_R g1345 ( 
.A(n_1226),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1294),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1209),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1271),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1276),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1254),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1277),
.Y(n_1351)
);

INVxp67_ASAP7_75t_SL g1352 ( 
.A(n_1247),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1298),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1238),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1224),
.A2(n_1210),
.B1(n_1207),
.B2(n_1317),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1207),
.B(n_1202),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1209),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1310),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1251),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1300),
.A2(n_1198),
.B(n_1212),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1208),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1219),
.A2(n_1204),
.B1(n_1214),
.B2(n_1317),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1222),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1317),
.A2(n_1279),
.B1(n_1219),
.B2(n_1233),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1251),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1198),
.A2(n_1206),
.B(n_1190),
.Y(n_1366)
);

CKINVDCx6p67_ASAP7_75t_R g1367 ( 
.A(n_1187),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1306),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1225),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1315),
.Y(n_1370)
);

BUFx8_ASAP7_75t_L g1371 ( 
.A(n_1231),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1241),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1172),
.B(n_1175),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1251),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1246),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1169),
.B(n_1173),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1244),
.A2(n_1242),
.B1(n_1229),
.B2(n_1228),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1232),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1195),
.Y(n_1379)
);

BUFx2_ASAP7_75t_SL g1380 ( 
.A(n_1232),
.Y(n_1380)
);

AO21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1227),
.A2(n_1260),
.B(n_1258),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1248),
.A2(n_1216),
.B(n_1249),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1169),
.A2(n_1316),
.B1(n_1173),
.B2(n_1203),
.Y(n_1383)
);

AO21x1_ASAP7_75t_L g1384 ( 
.A1(n_1213),
.A2(n_1211),
.B(n_1240),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1217),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1233),
.B(n_1178),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1233),
.A2(n_1203),
.B1(n_1316),
.B2(n_1292),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1221),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1299),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1230),
.A2(n_1201),
.B1(n_1312),
.B2(n_1235),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_1236),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1252),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1245),
.B(n_1259),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1253),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1236),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1267),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1282),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1261),
.A2(n_1273),
.B1(n_1256),
.B2(n_1302),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1270),
.A2(n_1263),
.B1(n_1264),
.B2(n_1262),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1255),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1250),
.A2(n_1275),
.B(n_1283),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1269),
.Y(n_1402)
);

BUFx8_ASAP7_75t_SL g1403 ( 
.A(n_1168),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1232),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1286),
.B(n_1287),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1262),
.A2(n_1264),
.B1(n_1266),
.B2(n_1268),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1170),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1280),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1284),
.B(n_1285),
.Y(n_1409)
);

BUFx4_ASAP7_75t_SL g1410 ( 
.A(n_1232),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1193),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1250),
.A2(n_1286),
.B(n_1281),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1193),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1265),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1215),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1215),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1234),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1234),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1272),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1265),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1288),
.A2(n_1313),
.B(n_1274),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1286),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1278),
.Y(n_1423)
);

INVx4_ASAP7_75t_L g1424 ( 
.A(n_1168),
.Y(n_1424)
);

BUFx2_ASAP7_75t_SL g1425 ( 
.A(n_1174),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1188),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1308),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1308),
.Y(n_1428)
);

INVx4_ASAP7_75t_L g1429 ( 
.A(n_1257),
.Y(n_1429)
);

BUFx4f_ASAP7_75t_SL g1430 ( 
.A(n_1187),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1291),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1191),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1185),
.B(n_1311),
.Y(n_1433)
);

BUFx2_ASAP7_75t_SL g1434 ( 
.A(n_1209),
.Y(n_1434)
);

CKINVDCx6p67_ASAP7_75t_R g1435 ( 
.A(n_1186),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1307),
.A2(n_1004),
.B1(n_1157),
.B2(n_941),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1209),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1291),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1191),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1184),
.B(n_993),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1251),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1289),
.B(n_857),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1251),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1412),
.A2(n_1360),
.B(n_1384),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1409),
.B(n_1324),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1349),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1349),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1361),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1339),
.B(n_1343),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1397),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1339),
.B(n_1343),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1351),
.B(n_1324),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1442),
.A2(n_1319),
.B1(n_1436),
.B2(n_1320),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1386),
.B(n_1422),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1363),
.Y(n_1455)
);

AO21x2_ASAP7_75t_L g1456 ( 
.A1(n_1326),
.A2(n_1366),
.B(n_1401),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1330),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1356),
.B(n_1321),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1351),
.B(n_1348),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1431),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1421),
.B(n_1423),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1386),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1433),
.B(n_1350),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1356),
.B(n_1391),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1386),
.A2(n_1325),
.B(n_1382),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1327),
.B(n_1333),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1433),
.B(n_1350),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1408),
.Y(n_1468)
);

INVx5_ASAP7_75t_L g1469 ( 
.A(n_1386),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1409),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1381),
.B(n_1423),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1397),
.Y(n_1472)
);

INVx4_ASAP7_75t_L g1473 ( 
.A(n_1347),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1399),
.B(n_1354),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1331),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1405),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1405),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1329),
.B(n_1340),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1381),
.B(n_1385),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1369),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1369),
.B(n_1372),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1392),
.B(n_1322),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1395),
.B(n_1354),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1379),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1373),
.B(n_1388),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1373),
.B(n_1389),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1394),
.B(n_1375),
.Y(n_1487)
);

BUFx2_ASAP7_75t_SL g1488 ( 
.A(n_1429),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1364),
.B(n_1383),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1338),
.A2(n_1440),
.B(n_1344),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1406),
.B(n_1400),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1347),
.Y(n_1492)
);

BUFx2_ASAP7_75t_SL g1493 ( 
.A(n_1429),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1328),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1332),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1355),
.A2(n_1396),
.B(n_1378),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1380),
.B(n_1434),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1334),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1322),
.B(n_1376),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1438),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1336),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1341),
.B(n_1370),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1352),
.B(n_1362),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1346),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1402),
.B(n_1432),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1368),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1439),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1410),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1335),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1407),
.A2(n_1411),
.B(n_1415),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1342),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1353),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1413),
.A2(n_1416),
.B(n_1417),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1418),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1419),
.B(n_1393),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1335),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1429),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1377),
.B(n_1387),
.C(n_1390),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1393),
.B(n_1426),
.Y(n_1519)
);

INVx4_ASAP7_75t_SL g1520 ( 
.A(n_1347),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1470),
.B(n_1445),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1512),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1464),
.B(n_1458),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1449),
.B(n_1451),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1449),
.B(n_1427),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1509),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1464),
.B(n_1358),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1451),
.B(n_1470),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1463),
.B(n_1427),
.Y(n_1529)
);

NOR2x1_ASAP7_75t_L g1530 ( 
.A(n_1488),
.B(n_1380),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1446),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1463),
.B(n_1428),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1458),
.B(n_1318),
.Y(n_1533)
);

BUFx4f_ASAP7_75t_L g1534 ( 
.A(n_1497),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1445),
.B(n_1318),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1446),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1467),
.B(n_1428),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1447),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1472),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1447),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1467),
.B(n_1428),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1444),
.B(n_1424),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1479),
.B(n_1452),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1472),
.B(n_1337),
.Y(n_1545)
);

OAI211xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1453),
.A2(n_1398),
.B(n_1323),
.C(n_1443),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1462),
.B(n_1434),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1509),
.B(n_1337),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1357),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1516),
.Y(n_1550)
);

NOR2x1_ASAP7_75t_L g1551 ( 
.A(n_1488),
.B(n_1404),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1454),
.B(n_1469),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1454),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1490),
.A2(n_1323),
.B1(n_1435),
.B2(n_1367),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1469),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1510),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1479),
.B(n_1424),
.Y(n_1557)
);

INVxp33_ASAP7_75t_L g1558 ( 
.A(n_1482),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1452),
.B(n_1425),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1516),
.B(n_1435),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1461),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1450),
.B(n_1367),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1450),
.B(n_1420),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1462),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1513),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1465),
.B(n_1420),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1459),
.B(n_1471),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1471),
.B(n_1420),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1485),
.B(n_1414),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1485),
.B(n_1414),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1486),
.B(n_1414),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1462),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1554),
.A2(n_1518),
.B1(n_1489),
.B2(n_1503),
.Y(n_1573)
);

NAND3xp33_ASAP7_75t_L g1574 ( 
.A(n_1549),
.B(n_1490),
.C(n_1466),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1526),
.Y(n_1575)
);

NAND4xp25_ASAP7_75t_L g1576 ( 
.A(n_1554),
.B(n_1478),
.C(n_1448),
.D(n_1511),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1544),
.B(n_1475),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1462),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1544),
.B(n_1524),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1523),
.B(n_1503),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1524),
.B(n_1475),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1528),
.B(n_1465),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1523),
.B(n_1448),
.Y(n_1583)
);

OAI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1546),
.A2(n_1499),
.B1(n_1455),
.B2(n_1500),
.C(n_1460),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1546),
.A2(n_1489),
.B1(n_1491),
.B2(n_1515),
.Y(n_1585)
);

NAND4xp25_ASAP7_75t_L g1586 ( 
.A(n_1533),
.B(n_1511),
.C(n_1505),
.D(n_1491),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1560),
.A2(n_1489),
.B1(n_1474),
.B2(n_1508),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1527),
.B(n_1457),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1528),
.B(n_1456),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1527),
.B(n_1474),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1533),
.B(n_1484),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1592)
);

OAI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1560),
.A2(n_1461),
.B1(n_1505),
.B2(n_1517),
.C(n_1508),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1562),
.A2(n_1489),
.B1(n_1522),
.B2(n_1548),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1567),
.B(n_1456),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1550),
.B(n_1486),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1521),
.B(n_1539),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1456),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1550),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1553),
.B(n_1456),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1535),
.B(n_1481),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1535),
.B(n_1481),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1553),
.B(n_1477),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1558),
.A2(n_1496),
.B(n_1517),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1521),
.B(n_1481),
.Y(n_1605)
);

NAND3xp33_ASAP7_75t_L g1606 ( 
.A(n_1548),
.B(n_1504),
.C(n_1494),
.Y(n_1606)
);

OAI221xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1566),
.A2(n_1483),
.B1(n_1517),
.B2(n_1495),
.C(n_1507),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1525),
.B(n_1529),
.Y(n_1608)
);

OAI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1545),
.A2(n_1483),
.B(n_1502),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1525),
.B(n_1481),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1529),
.B(n_1498),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1532),
.B(n_1498),
.Y(n_1612)
);

NAND3xp33_ASAP7_75t_L g1613 ( 
.A(n_1545),
.B(n_1504),
.C(n_1506),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1566),
.A2(n_1501),
.B1(n_1506),
.B2(n_1507),
.C(n_1495),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1553),
.B(n_1532),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1562),
.B(n_1519),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1552),
.A2(n_1462),
.B(n_1461),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1553),
.B(n_1477),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1537),
.B(n_1498),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1537),
.B(n_1468),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1541),
.B(n_1477),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1541),
.B(n_1468),
.Y(n_1622)
);

OAI221xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1542),
.A2(n_1501),
.B1(n_1494),
.B2(n_1497),
.C(n_1476),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1569),
.B(n_1468),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_L g1625 ( 
.A(n_1551),
.B(n_1473),
.C(n_1496),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1531),
.Y(n_1626)
);

OAI211xp5_ASAP7_75t_L g1627 ( 
.A1(n_1542),
.A2(n_1502),
.B(n_1487),
.C(n_1480),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1542),
.B(n_1444),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_SL g1629 ( 
.A1(n_1552),
.A2(n_1462),
.B(n_1515),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1543),
.B(n_1476),
.C(n_1514),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1597),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1626),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1615),
.B(n_1552),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1626),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1615),
.B(n_1552),
.Y(n_1635)
);

INVx5_ASAP7_75t_SL g1636 ( 
.A(n_1578),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1582),
.B(n_1543),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1590),
.B(n_1539),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1583),
.B(n_1570),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1599),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1580),
.B(n_1570),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1588),
.B(n_1430),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1597),
.Y(n_1643)
);

NOR2xp67_ASAP7_75t_L g1644 ( 
.A(n_1606),
.B(n_1555),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1582),
.B(n_1543),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1575),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1592),
.Y(n_1647)
);

NAND4xp25_ASAP7_75t_L g1648 ( 
.A(n_1574),
.B(n_1563),
.C(n_1561),
.D(n_1487),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1613),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1589),
.B(n_1444),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1589),
.B(n_1565),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1574),
.A2(n_1571),
.B1(n_1538),
.B2(n_1536),
.C(n_1540),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1581),
.B(n_1564),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1628),
.B(n_1565),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1591),
.B(n_1571),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1613),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1628),
.B(n_1556),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1606),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1601),
.B(n_1563),
.Y(n_1659)
);

NAND4xp25_ASAP7_75t_SL g1660 ( 
.A(n_1585),
.B(n_1530),
.C(n_1557),
.D(n_1551),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1603),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1602),
.B(n_1605),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1603),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1581),
.B(n_1564),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1609),
.B(n_1568),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1618),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1609),
.B(n_1568),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1595),
.B(n_1556),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1596),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1618),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1595),
.B(n_1564),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1612),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1619),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1611),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1625),
.B(n_1561),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1598),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1647),
.B(n_1579),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1579),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1663),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1669),
.B(n_1621),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1649),
.B(n_1621),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1632),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1640),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_R g1684 ( 
.A(n_1660),
.B(n_1371),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1656),
.B(n_1598),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1663),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1654),
.B(n_1608),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1654),
.B(n_1586),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1637),
.B(n_1577),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1653),
.Y(n_1690)
);

AND2x4_ASAP7_75t_SL g1691 ( 
.A(n_1675),
.B(n_1547),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1634),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1646),
.Y(n_1693)
);

NAND2x1_ASAP7_75t_L g1694 ( 
.A(n_1644),
.B(n_1630),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1643),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1658),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1674),
.B(n_1577),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1651),
.B(n_1630),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1637),
.B(n_1617),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1645),
.B(n_1629),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1658),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1672),
.B(n_1610),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1651),
.B(n_1620),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1631),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1631),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1673),
.B(n_1616),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1657),
.B(n_1622),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1657),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1645),
.B(n_1600),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1638),
.B(n_1624),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1668),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1659),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1661),
.B(n_1600),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1642),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1636),
.A2(n_1585),
.B1(n_1584),
.B2(n_1573),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1714),
.B(n_1576),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1714),
.B(n_1345),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1699),
.B(n_1633),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1699),
.B(n_1633),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1715),
.A2(n_1578),
.B(n_1652),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1679),
.Y(n_1721)
);

NOR2x1p5_ASAP7_75t_L g1722 ( 
.A(n_1694),
.B(n_1648),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1696),
.B(n_1650),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1682),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1682),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1692),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1683),
.B(n_1665),
.Y(n_1727)
);

AOI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1684),
.A2(n_1594),
.B(n_1593),
.C(n_1587),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1700),
.B(n_1635),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1700),
.B(n_1635),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1694),
.Y(n_1731)
);

NOR2xp67_ASAP7_75t_L g1732 ( 
.A(n_1698),
.B(n_1661),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1701),
.B(n_1650),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1712),
.B(n_1667),
.Y(n_1734)
);

NAND3xp33_ASAP7_75t_L g1735 ( 
.A(n_1693),
.B(n_1604),
.C(n_1623),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1679),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1686),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1692),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1688),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1695),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1688),
.A2(n_1675),
.B(n_1641),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1685),
.B(n_1668),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1708),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1676),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1681),
.B(n_1671),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1689),
.B(n_1636),
.Y(n_1746)
);

INVxp67_ASAP7_75t_SL g1747 ( 
.A(n_1704),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1689),
.B(n_1636),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1708),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1706),
.B(n_1671),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1677),
.B(n_1662),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1691),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1691),
.B(n_1636),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1655),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1705),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1710),
.B(n_1675),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1711),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1690),
.B(n_1661),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1724),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1721),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1729),
.B(n_1709),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1758),
.Y(n_1762)
);

CKINVDCx16_ASAP7_75t_R g1763 ( 
.A(n_1717),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1722),
.A2(n_1720),
.B1(n_1716),
.B2(n_1735),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1739),
.B(n_1687),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1755),
.B(n_1678),
.Y(n_1766)
);

CKINVDCx16_ASAP7_75t_R g1767 ( 
.A(n_1731),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1741),
.A2(n_1702),
.B1(n_1680),
.B2(n_1697),
.C(n_1690),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1728),
.A2(n_1627),
.B1(n_1547),
.B2(n_1519),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1751),
.B(n_1687),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1731),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1721),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1729),
.B(n_1709),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1703),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1730),
.B(n_1713),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1730),
.B(n_1713),
.Y(n_1776)
);

AOI222xp33_ASAP7_75t_L g1777 ( 
.A1(n_1756),
.A2(n_1686),
.B1(n_1639),
.B2(n_1534),
.C1(n_1371),
.C2(n_1664),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1752),
.B(n_1727),
.Y(n_1778)
);

CKINVDCx16_ASAP7_75t_R g1779 ( 
.A(n_1753),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1734),
.B(n_1750),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1753),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1724),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1746),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1725),
.Y(n_1784)
);

AOI222xp33_ASAP7_75t_L g1785 ( 
.A1(n_1732),
.A2(n_1534),
.B1(n_1371),
.B2(n_1653),
.C1(n_1664),
.C2(n_1559),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1744),
.B(n_1754),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1736),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1746),
.A2(n_1607),
.B1(n_1703),
.B2(n_1707),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1718),
.B(n_1707),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1725),
.Y(n_1790)
);

INVxp67_ASAP7_75t_SL g1791 ( 
.A(n_1748),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1740),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1726),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1718),
.B(n_1666),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1791),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1779),
.B(n_1719),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1792),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1767),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1779),
.B(n_1719),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1764),
.B(n_1740),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1778),
.A2(n_1757),
.B1(n_1743),
.B2(n_1749),
.C(n_1726),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1783),
.B(n_1781),
.Y(n_1802)
);

NOR2x1_ASAP7_75t_L g1803 ( 
.A(n_1781),
.B(n_1738),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1763),
.B(n_1748),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1759),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1759),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1763),
.B(n_1754),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1781),
.B(n_1743),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1762),
.Y(n_1809)
);

BUFx2_ASAP7_75t_SL g1810 ( 
.A(n_1771),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1769),
.A2(n_1767),
.B1(n_1777),
.B2(n_1788),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1762),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1780),
.B(n_1745),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1769),
.B(n_1758),
.Y(n_1814)
);

AOI21xp33_ASAP7_75t_L g1815 ( 
.A1(n_1765),
.A2(n_1757),
.B(n_1749),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1782),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1765),
.B(n_1758),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1782),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1784),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1775),
.B(n_1744),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1810),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1805),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1806),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1807),
.B(n_1771),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1795),
.B(n_1786),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1816),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1804),
.B(n_1786),
.Y(n_1827)
);

INVxp67_ASAP7_75t_SL g1828 ( 
.A(n_1804),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1796),
.B(n_1775),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1818),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1796),
.B(n_1776),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1819),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1798),
.B(n_1770),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1802),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1797),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1799),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1799),
.B(n_1776),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1800),
.B(n_1774),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1803),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1812),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_SL g1841 ( 
.A(n_1821),
.B(n_1811),
.C(n_1801),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1836),
.B(n_1817),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1825),
.B(n_1817),
.Y(n_1843)
);

AOI311xp33_ASAP7_75t_L g1844 ( 
.A1(n_1827),
.A2(n_1809),
.A3(n_1815),
.B(n_1808),
.C(n_1813),
.Y(n_1844)
);

AOI211xp5_ASAP7_75t_L g1845 ( 
.A1(n_1828),
.A2(n_1814),
.B(n_1812),
.C(n_1820),
.Y(n_1845)
);

NAND4xp25_ASAP7_75t_L g1846 ( 
.A(n_1833),
.B(n_1814),
.C(n_1820),
.D(n_1785),
.Y(n_1846)
);

OAI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1839),
.A2(n_1784),
.B(n_1793),
.C(n_1790),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_L g1848 ( 
.A(n_1834),
.B(n_1824),
.C(n_1825),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1838),
.A2(n_1834),
.B(n_1831),
.Y(n_1849)
);

OAI32xp33_ASAP7_75t_L g1850 ( 
.A1(n_1838),
.A2(n_1793),
.A3(n_1790),
.B1(n_1766),
.B2(n_1789),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1829),
.B(n_1794),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1840),
.Y(n_1852)
);

NOR2x1_ASAP7_75t_SL g1853 ( 
.A(n_1842),
.B(n_1840),
.Y(n_1853)
);

NAND4xp75_ASAP7_75t_L g1854 ( 
.A(n_1849),
.B(n_1835),
.C(n_1837),
.D(n_1831),
.Y(n_1854)
);

NAND3xp33_ASAP7_75t_SL g1855 ( 
.A(n_1845),
.B(n_1837),
.C(n_1829),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_L g1856 ( 
.A(n_1844),
.B(n_1823),
.C(n_1822),
.Y(n_1856)
);

OAI322xp33_ASAP7_75t_L g1857 ( 
.A1(n_1843),
.A2(n_1830),
.A3(n_1826),
.B1(n_1832),
.B2(n_1760),
.C1(n_1787),
.C2(n_1772),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1852),
.B(n_1832),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1851),
.B(n_1761),
.Y(n_1859)
);

NOR4xp75_ASAP7_75t_L g1860 ( 
.A(n_1841),
.B(n_1768),
.C(n_1761),
.D(n_1773),
.Y(n_1860)
);

OAI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1848),
.A2(n_1772),
.B(n_1760),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1847),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1853),
.A2(n_1846),
.B(n_1850),
.Y(n_1863)
);

AND4x1_ASAP7_75t_L g1864 ( 
.A(n_1856),
.B(n_1773),
.C(n_1794),
.D(n_1738),
.Y(n_1864)
);

NAND4xp75_ASAP7_75t_L g1865 ( 
.A(n_1862),
.B(n_1858),
.C(n_1861),
.D(n_1859),
.Y(n_1865)
);

NOR2x1_ASAP7_75t_L g1866 ( 
.A(n_1854),
.B(n_1787),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1855),
.B(n_1736),
.Y(n_1867)
);

OAI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1860),
.A2(n_1733),
.B(n_1723),
.C(n_1737),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1867),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1863),
.A2(n_1737),
.B1(n_1733),
.B2(n_1723),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1864),
.B(n_1742),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1865),
.B(n_1857),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1868),
.A2(n_1742),
.B1(n_1493),
.B2(n_1534),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1866),
.A2(n_1493),
.B1(n_1534),
.B2(n_1557),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1867),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1863),
.A2(n_1547),
.B1(n_1572),
.B2(n_1564),
.Y(n_1876)
);

NAND4xp25_ASAP7_75t_SL g1877 ( 
.A(n_1872),
.B(n_1403),
.C(n_1670),
.D(n_1559),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1869),
.Y(n_1878)
);

INVxp67_ASAP7_75t_SL g1879 ( 
.A(n_1870),
.Y(n_1879)
);

OA22x2_ASAP7_75t_L g1880 ( 
.A1(n_1873),
.A2(n_1497),
.B1(n_1547),
.B2(n_1666),
.Y(n_1880)
);

NOR2x1_ASAP7_75t_L g1881 ( 
.A(n_1875),
.B(n_1365),
.Y(n_1881)
);

NAND3x1_ASAP7_75t_L g1882 ( 
.A(n_1881),
.B(n_1876),
.C(n_1871),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1879),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1878),
.B(n_1874),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1883),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1885),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1886),
.Y(n_1887)
);

NOR4xp75_ASAP7_75t_L g1888 ( 
.A(n_1886),
.B(n_1882),
.C(n_1884),
.D(n_1877),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1887),
.Y(n_1889)
);

OA21x2_ASAP7_75t_L g1890 ( 
.A1(n_1888),
.A2(n_1880),
.B(n_1359),
.Y(n_1890)
);

NOR2xp67_ASAP7_75t_L g1891 ( 
.A(n_1889),
.B(n_1359),
.Y(n_1891)
);

NAND2x1p5_ASAP7_75t_L g1892 ( 
.A(n_1890),
.B(n_1365),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1892),
.A2(n_1891),
.B(n_1890),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1893),
.A2(n_1890),
.B1(n_1403),
.B2(n_1374),
.Y(n_1894)
);

OAI221xp5_ASAP7_75t_R g1895 ( 
.A1(n_1894),
.A2(n_1374),
.B1(n_1441),
.B2(n_1520),
.C(n_1614),
.Y(n_1895)
);

AOI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1895),
.A2(n_1357),
.B(n_1437),
.C(n_1492),
.Y(n_1896)
);


endmodule