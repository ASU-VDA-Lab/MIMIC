module fake_jpeg_27777_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_23),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_31)
);

NAND2x1_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_24),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_25),
.C(n_27),
.Y(n_39)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_43),
.B(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_22),
.B1(n_16),
.B2(n_15),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_44),
.B1(n_46),
.B2(n_43),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_15),
.B1(n_16),
.B2(n_13),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_30),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_30),
.A2(n_27),
.B1(n_19),
.B2(n_17),
.Y(n_46)
);

CKINVDCx9p33_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_63),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_58),
.B1(n_64),
.B2(n_71),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_32),
.C(n_25),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_71),
.C(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_26),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_68),
.B1(n_38),
.B2(n_35),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_14),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_14),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_25),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_25),
.B(n_21),
.C(n_32),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_33),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_36),
.B(n_29),
.C(n_37),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_50),
.B1(n_47),
.B2(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_53),
.B(n_35),
.C(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_70),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_59),
.B1(n_21),
.B2(n_18),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_72),
.C(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_65),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_93),
.C(n_76),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_76),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_32),
.C(n_73),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_96),
.B1(n_101),
.B2(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_2),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_87),
.C(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_11),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_93),
.B1(n_95),
.B2(n_101),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_105),
.B1(n_82),
.B2(n_88),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_4),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_76),
.C(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_111),
.Y(n_119)
);

AO221x1_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_82),
.B1(n_83),
.B2(n_88),
.C(n_3),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_116),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_102),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_114),
.B(n_115),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_18),
.C(n_23),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_120),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_109),
.B(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_116),
.Y(n_122)
);

AOI211xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_123),
.B(n_11),
.C(n_5),
.Y(n_127)
);

AOI31xp33_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_104),
.A3(n_5),
.B(n_4),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_6),
.C(n_10),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_6),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_123),
.B(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_126),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_129),
.Y(n_131)
);


endmodule