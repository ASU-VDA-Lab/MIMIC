module fake_netlist_1_2065_n_33 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_7;
wire n_27;
INVxp67_ASAP7_75t_SL g7 ( .A(n_6), .Y(n_7) );
INVx3_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
CKINVDCx16_ASAP7_75t_R g9 ( .A(n_5), .Y(n_9) );
NAND2xp33_ASAP7_75t_L g10 ( .A(n_5), .B(n_0), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_9), .Y(n_13) );
BUFx12f_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_9), .B(n_0), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_8), .B(n_1), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
AOI222xp33_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_7), .B1(n_10), .B2(n_12), .C1(n_8), .C2(n_3), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_15), .B(n_8), .Y(n_19) );
NAND3xp33_ASAP7_75t_L g20 ( .A(n_16), .B(n_12), .C(n_8), .Y(n_20) );
NOR3xp33_ASAP7_75t_SL g21 ( .A(n_13), .B(n_7), .C(n_2), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_19), .B(n_14), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_19), .B(n_14), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
OAI222xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_12), .B1(n_21), .B2(n_17), .C1(n_14), .C2(n_4), .Y(n_26) );
NAND4xp25_ASAP7_75t_L g27 ( .A(n_25), .B(n_23), .C(n_20), .D(n_24), .Y(n_27) );
NOR2xp33_ASAP7_75t_SL g28 ( .A(n_26), .B(n_17), .Y(n_28) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_28), .Y(n_29) );
INVxp67_ASAP7_75t_SL g30 ( .A(n_27), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_29), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_17), .B1(n_1), .B2(n_3), .Y(n_32) );
OAI21xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_30), .B(n_31), .Y(n_33) );
endmodule