module fake_jpeg_12250_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_17),
.C(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_64),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_52),
.B1(n_43),
.B2(n_42),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_62),
.B1(n_65),
.B2(n_54),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_70),
.B1(n_52),
.B2(n_59),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_71),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_1),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_67),
.B1(n_12),
.B2(n_10),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_58),
.B(n_48),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_50),
.C(n_49),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_18),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_7),
.B(n_9),
.Y(n_98)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_6),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_92),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

OAI221xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_67),
.B1(n_11),
.B2(n_12),
.C(n_10),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_85),
.B1(n_79),
.B2(n_84),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_26),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_100),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_13),
.B(n_14),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_29),
.B(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_105),
.B(n_102),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_115),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_120),
.B(n_111),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_100),
.C(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_112),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_117),
.B1(n_113),
.B2(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_122),
.B(n_123),
.Y(n_124)
);

NAND2x1p5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_119),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_105),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_103),
.A3(n_116),
.B1(n_97),
.B2(n_109),
.C1(n_33),
.C2(n_38),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_34),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_116),
.Y(n_129)
);


endmodule