module real_aes_16897_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_855, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_855;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
AND2x4_ASAP7_75t_L g849 ( .A(n_0), .B(n_850), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_1), .A2(n_32), .B1(n_151), .B2(n_188), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_2), .A2(n_9), .B1(n_535), .B2(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g850 ( .A(n_3), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_4), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_5), .A2(n_10), .B1(n_571), .B2(n_572), .Y(n_570) );
OR2x2_ASAP7_75t_L g113 ( .A(n_6), .B(n_28), .Y(n_113) );
BUFx2_ASAP7_75t_L g843 ( .A(n_6), .Y(n_843) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_7), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_8), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_11), .B(n_172), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_12), .A2(n_95), .B1(n_244), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_13), .A2(n_29), .B1(n_552), .B2(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_14), .B(n_172), .Y(n_549) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_15), .A2(n_43), .B(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_16), .B(n_219), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_17), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_18), .A2(n_84), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_18), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_19), .A2(n_36), .B1(n_150), .B2(n_249), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_20), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_21), .A2(n_41), .B1(n_150), .B2(n_535), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_22), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_23), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_24), .B(n_182), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_25), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_26), .B(n_159), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_27), .Y(n_243) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_28), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_30), .A2(n_79), .B1(n_151), .B2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_31), .A2(n_35), .B1(n_151), .B2(n_548), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_33), .A2(n_46), .B1(n_535), .B2(n_537), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_34), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_37), .B(n_172), .Y(n_203) );
INVx2_ASAP7_75t_L g502 ( .A(n_38), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_39), .B(n_207), .Y(n_214) );
INVx1_ASAP7_75t_L g111 ( .A(n_40), .Y(n_111) );
BUFx3_ASAP7_75t_L g511 ( .A(n_40), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_42), .B(n_154), .Y(n_222) );
AND2x2_ASAP7_75t_L g153 ( .A(n_44), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_45), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_47), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_48), .B(n_249), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_49), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_50), .A2(n_67), .B1(n_249), .B2(n_537), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_51), .A2(n_70), .B1(n_151), .B2(n_548), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_52), .B(n_187), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_53), .A2(n_136), .B(n_138), .C(n_141), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_54), .B(n_829), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_55), .A2(n_92), .B1(n_535), .B2(n_572), .Y(n_612) );
INVx1_ASAP7_75t_L g129 ( .A(n_56), .Y(n_129) );
AND2x4_ASAP7_75t_L g132 ( .A(n_57), .B(n_133), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_58), .A2(n_59), .B1(n_150), .B2(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_60), .B(n_159), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_61), .B(n_154), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_62), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_63), .B(n_150), .Y(n_206) );
INVx1_ASAP7_75t_L g133 ( .A(n_64), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_65), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_66), .B(n_159), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_68), .B(n_151), .Y(n_180) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_69), .B(n_188), .C(n_207), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_71), .B(n_151), .Y(n_163) );
INVx2_ASAP7_75t_L g143 ( .A(n_72), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_73), .B(n_172), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_74), .B(n_221), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_75), .B(n_168), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_76), .A2(n_91), .B1(n_136), .B2(n_150), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_77), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_78), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_80), .A2(n_86), .B1(n_182), .B2(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_81), .B(n_172), .Y(n_245) );
NAND2xp33_ASAP7_75t_SL g276 ( .A(n_82), .B(n_165), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_83), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g492 ( .A(n_84), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_84), .B(n_115), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_85), .B(n_159), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_87), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_88), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g520 ( .A(n_88), .Y(n_520) );
NAND2xp33_ASAP7_75t_L g553 ( .A(n_89), .B(n_172), .Y(n_553) );
NAND2xp33_ASAP7_75t_L g164 ( .A(n_90), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_93), .B(n_154), .Y(n_190) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_94), .B(n_165), .C(n_221), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g100 ( .A1(n_96), .A2(n_101), .B1(n_839), .B2(n_853), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_97), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_98), .B(n_151), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_99), .B(n_182), .Y(n_185) );
OR2x6_ASAP7_75t_L g101 ( .A(n_102), .B(n_493), .Y(n_101) );
NAND3x1_ASAP7_75t_L g102 ( .A(n_103), .B(n_503), .C(n_836), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_498), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_114), .B(n_493), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx5_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx8_ASAP7_75t_R g497 ( .A(n_108), .Y(n_497) );
AND2x6_ASAP7_75t_SL g108 ( .A(n_109), .B(n_112), .Y(n_108) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_111), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_112), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NOR2x1_ASAP7_75t_L g835 ( .A(n_113), .B(n_511), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_116), .B1(n_489), .B2(n_490), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_116), .A2(n_492), .B(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_377), .Y(n_116) );
NOR4xp75_ASAP7_75t_L g117 ( .A(n_118), .B(n_316), .C(n_340), .D(n_359), .Y(n_117) );
NAND3x1_ASAP7_75t_L g118 ( .A(n_119), .B(n_256), .C(n_307), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_191), .B1(n_234), .B2(n_252), .Y(n_119) );
AND2x2_ASAP7_75t_L g438 ( .A(n_120), .B(n_313), .Y(n_438) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_156), .Y(n_120) );
AND2x2_ASAP7_75t_L g388 ( .A(n_121), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_121), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g415 ( .A(n_121), .Y(n_415) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g260 ( .A(n_122), .Y(n_260) );
INVx2_ASAP7_75t_L g282 ( .A(n_122), .Y(n_282) );
AND2x2_ASAP7_75t_L g376 ( .A(n_122), .B(n_339), .Y(n_376) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g255 ( .A(n_123), .Y(n_255) );
AND2x2_ASAP7_75t_L g355 ( .A(n_123), .B(n_267), .Y(n_355) );
AOI21x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_134), .B(n_153), .Y(n_123) );
NOR2xp67_ASAP7_75t_SL g124 ( .A(n_125), .B(n_130), .Y(n_124) );
INVx2_ASAP7_75t_L g538 ( .A(n_125), .Y(n_538) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_126), .A2(n_131), .A3(n_225), .B(n_231), .Y(n_224) );
NOR2xp33_ASAP7_75t_SL g576 ( .A(n_126), .B(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_126), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx2_ASAP7_75t_L g233 ( .A(n_127), .Y(n_233) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
INVx1_ASAP7_75t_L g532 ( .A(n_130), .Y(n_532) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AO31x2_ASAP7_75t_L g558 ( .A1(n_131), .A2(n_559), .A3(n_562), .B(n_563), .Y(n_558) );
AO31x2_ASAP7_75t_L g568 ( .A1(n_131), .A2(n_569), .A3(n_575), .B(n_576), .Y(n_568) );
AO31x2_ASAP7_75t_L g579 ( .A1(n_131), .A2(n_580), .A3(n_585), .B(n_586), .Y(n_579) );
BUFx10_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx10_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
INVx1_ASAP7_75t_L g555 ( .A(n_132), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_144), .Y(n_134) );
INVx1_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g140 ( .A(n_137), .Y(n_140) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_137), .Y(n_151) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
INVx1_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_137), .Y(n_188) );
INVx1_ASAP7_75t_L g202 ( .A(n_137), .Y(n_202) );
INVx1_ASAP7_75t_L g230 ( .A(n_137), .Y(n_230) );
INVx1_ASAP7_75t_L g275 ( .A(n_137), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
INVx2_ASAP7_75t_SL g593 ( .A(n_140), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_141), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_141), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_141), .A2(n_201), .B(n_203), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_141), .A2(n_274), .B(n_276), .Y(n_273) );
BUFx4f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g147 ( .A(n_143), .Y(n_147) );
BUFx8_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
INVx1_ASAP7_75t_L g221 ( .A(n_143), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_148), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_145), .A2(n_226), .B1(n_228), .B2(n_229), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_145), .A2(n_228), .B1(n_534), .B2(n_536), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_145), .A2(n_228), .B1(n_560), .B2(n_561), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_145), .A2(n_228), .B1(n_581), .B2(n_583), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_145), .A2(n_228), .B1(n_631), .B2(n_632), .Y(n_630) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g169 ( .A(n_147), .Y(n_169) );
OAI22xp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B1(n_151), .B2(n_152), .Y(n_148) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_150), .A2(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g227 ( .A(n_150), .Y(n_227) );
INVx1_ASAP7_75t_L g537 ( .A(n_151), .Y(n_537) );
INVx4_ASAP7_75t_L g548 ( .A(n_151), .Y(n_548) );
INVx1_ASAP7_75t_L g572 ( .A(n_151), .Y(n_572) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_155), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_155), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g308 ( .A(n_156), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g423 ( .A(n_156), .Y(n_423) );
AND2x2_ASAP7_75t_L g429 ( .A(n_156), .B(n_293), .Y(n_429) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_175), .Y(n_156) );
INVx1_ASAP7_75t_L g265 ( .A(n_157), .Y(n_265) );
INVx4_ASAP7_75t_L g286 ( .A(n_157), .Y(n_286) );
OR2x2_ASAP7_75t_L g335 ( .A(n_157), .B(n_315), .Y(n_335) );
BUFx2_ASAP7_75t_L g404 ( .A(n_157), .Y(n_404) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_161), .Y(n_157) );
INVx2_ASAP7_75t_L g562 ( .A(n_159), .Y(n_562) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_SL g173 ( .A(n_160), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g198 ( .A(n_160), .Y(n_198) );
INVx1_ASAP7_75t_SL g268 ( .A(n_160), .Y(n_268) );
INVx2_ASAP7_75t_SL g544 ( .A(n_160), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_160), .B(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g585 ( .A(n_160), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_160), .B(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_160), .B(n_615), .Y(n_614) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_166), .B(n_173), .Y(n_161) );
INVx2_ASAP7_75t_L g249 ( .A(n_165), .Y(n_249) );
INVx1_ASAP7_75t_L g552 ( .A(n_165), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_168), .A2(n_247), .B(n_248), .Y(n_246) );
INVx2_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g219 ( .A(n_172), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_172), .A2(n_271), .B(n_272), .Y(n_270) );
INVx3_ASAP7_75t_L g535 ( .A(n_172), .Y(n_535) );
OAI21x1_ASAP7_75t_L g178 ( .A1(n_174), .A2(n_179), .B(n_184), .Y(n_178) );
OAI21x1_ASAP7_75t_L g199 ( .A1(n_174), .A2(n_200), .B(n_204), .Y(n_199) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_174), .A2(n_213), .B(n_216), .Y(n_212) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_174), .A2(n_242), .B(n_246), .Y(n_241) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_174), .A2(n_270), .B(n_273), .Y(n_269) );
AND2x2_ASAP7_75t_L g254 ( .A(n_175), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g357 ( .A(n_175), .Y(n_357) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g281 ( .A(n_176), .Y(n_281) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_190), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_177), .A2(n_241), .B(n_250), .Y(n_240) );
OAI21xp33_ASAP7_75t_SL g295 ( .A1(n_177), .A2(n_178), .B(n_190), .Y(n_295) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_177), .A2(n_241), .B(n_250), .Y(n_306) );
INVx1_ASAP7_75t_L g571 ( .A(n_182), .Y(n_571) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_189), .Y(n_184) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2x1_ASAP7_75t_L g426 ( .A(n_193), .B(n_366), .Y(n_426) );
AND2x4_ASAP7_75t_L g193 ( .A(n_194), .B(n_209), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OR2x2_ASAP7_75t_L g311 ( .A(n_195), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g331 ( .A(n_195), .B(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_195), .Y(n_365) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g321 ( .A(n_196), .B(n_211), .Y(n_321) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_196), .B(n_210), .Y(n_476) );
BUFx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g398 ( .A(n_197), .Y(n_398) );
OAI21x1_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_208), .Y(n_197) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_198), .A2(n_212), .B(n_222), .Y(n_211) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_198), .A2(n_199), .B(n_208), .Y(n_238) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_198), .A2(n_212), .B(n_222), .Y(n_251) );
INVx2_ASAP7_75t_L g244 ( .A(n_202), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
INVx6_ASAP7_75t_L g228 ( .A(n_207), .Y(n_228) );
O2A1O1Ixp5_ASAP7_75t_L g242 ( .A1(n_207), .A2(n_243), .B(n_244), .C(n_245), .Y(n_242) );
O2A1O1Ixp5_ASAP7_75t_L g546 ( .A1(n_207), .A2(n_547), .B(n_548), .C(n_549), .Y(n_546) );
INVx2_ASAP7_75t_L g419 ( .A(n_209), .Y(n_419) );
AND2x4_ASAP7_75t_L g457 ( .A(n_209), .B(n_396), .Y(n_457) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_223), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g297 ( .A(n_211), .Y(n_297) );
AND2x2_ASAP7_75t_L g332 ( .A(n_211), .B(n_224), .Y(n_332) );
AND2x2_ASAP7_75t_L g455 ( .A(n_211), .B(n_305), .Y(n_455) );
AND2x2_ASAP7_75t_L g466 ( .A(n_211), .B(n_240), .Y(n_466) );
AOI21x1_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_220), .Y(n_216) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_SL g574 ( .A(n_221), .Y(n_574) );
INVx1_ASAP7_75t_L g595 ( .A(n_221), .Y(n_595) );
AND2x2_ASAP7_75t_L g324 ( .A(n_223), .B(n_238), .Y(n_324) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g237 ( .A(n_224), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g298 ( .A(n_224), .B(n_238), .Y(n_298) );
OR2x2_ASAP7_75t_L g312 ( .A(n_224), .B(n_251), .Y(n_312) );
AND2x2_ASAP7_75t_L g397 ( .A(n_224), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_224), .B(n_251), .Y(n_408) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_224), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_228), .A2(n_551), .B(n_553), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_228), .A2(n_570), .B1(n_573), .B2(n_574), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_228), .A2(n_592), .B1(n_594), .B2(n_595), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_228), .A2(n_574), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g584 ( .A(n_230), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
BUFx2_ASAP7_75t_L g575 ( .A(n_233), .Y(n_575) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_239), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g346 ( .A(n_237), .Y(n_346) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_237), .B(n_454), .C(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g290 ( .A(n_238), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_239), .B(n_298), .Y(n_420) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_251), .Y(n_239) );
INVx1_ASAP7_75t_L g263 ( .A(n_240), .Y(n_263) );
AND2x2_ASAP7_75t_L g469 ( .A(n_251), .B(n_305), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_252), .Y(n_472) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g451 ( .A(n_253), .B(n_284), .Y(n_451) );
OR2x2_ASAP7_75t_L g462 ( .A(n_253), .B(n_335), .Y(n_462) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g338 ( .A(n_254), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g486 ( .A(n_254), .B(n_264), .Y(n_486) );
AND2x2_ASAP7_75t_L g294 ( .A(n_255), .B(n_295), .Y(n_294) );
A2O1A1O1Ixp25_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_261), .B(n_278), .C(n_287), .D(n_291), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g372 ( .A(n_259), .B(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g309 ( .A(n_260), .Y(n_309) );
INVx1_ASAP7_75t_L g344 ( .A(n_261), .Y(n_344) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g323 ( .A(n_262), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g314 ( .A(n_263), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g343 ( .A(n_264), .Y(n_343) );
AND2x2_ASAP7_75t_L g414 ( .A(n_264), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g460 ( .A(n_264), .B(n_294), .Y(n_460) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g285 ( .A(n_266), .Y(n_285) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_266), .Y(n_293) );
INVx2_ASAP7_75t_L g339 ( .A(n_266), .Y(n_339) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g315 ( .A(n_267), .Y(n_315) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_277), .Y(n_267) );
INVx1_ASAP7_75t_L g582 ( .A(n_275), .Y(n_582) );
INVx1_ASAP7_75t_L g410 ( .A(n_278), .Y(n_410) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_283), .Y(n_278) );
OAI21xp33_ASAP7_75t_L g334 ( .A1(n_279), .A2(n_284), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
AND2x2_ASAP7_75t_L g300 ( .A(n_280), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g405 ( .A(n_280), .B(n_355), .Y(n_405) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g337 ( .A(n_281), .B(n_315), .Y(n_337) );
AND2x2_ASAP7_75t_L g361 ( .A(n_282), .B(n_286), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_282), .B(n_301), .Y(n_445) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_SL g389 ( .A(n_284), .Y(n_389) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx2_ASAP7_75t_L g301 ( .A(n_286), .Y(n_301) );
NAND2x1_ASAP7_75t_L g356 ( .A(n_286), .B(n_357), .Y(n_356) );
OAI32xp33_ASAP7_75t_L g477 ( .A1(n_287), .A2(n_353), .A3(n_461), .B1(n_478), .B2(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g351 ( .A(n_289), .Y(n_351) );
AND2x2_ASAP7_75t_L g374 ( .A(n_289), .B(n_332), .Y(n_374) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g371 ( .A(n_290), .B(n_305), .Y(n_371) );
OAI22xp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_296), .B1(n_299), .B2(n_302), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g328 ( .A(n_294), .B(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g347 ( .A(n_295), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx2_ASAP7_75t_L g461 ( .A(n_297), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_298), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g440 ( .A(n_298), .Y(n_440) );
AND2x2_ASAP7_75t_L g468 ( .A(n_298), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g375 ( .A(n_300), .B(n_376), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g424 ( .A1(n_300), .A2(n_355), .B(n_425), .C(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
AND2x2_ASAP7_75t_L g373 ( .A(n_301), .B(n_339), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_303), .B(n_324), .Y(n_342) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_305), .Y(n_320) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_305), .Y(n_367) );
INVx1_ASAP7_75t_L g396 ( .A(n_305), .Y(n_396) );
BUFx3_ASAP7_75t_L g409 ( .A(n_305), .Y(n_409) );
INVx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND3xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .C(n_313), .Y(n_307) );
INVx1_ASAP7_75t_L g431 ( .A(n_308), .Y(n_431) );
OR2x2_ASAP7_75t_L g358 ( .A(n_309), .B(n_343), .Y(n_358) );
OR2x2_ASAP7_75t_L g322 ( .A(n_310), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_311), .A2(n_349), .B1(n_353), .B2(n_358), .Y(n_348) );
INVx2_ASAP7_75t_L g352 ( .A(n_312), .Y(n_352) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_312), .Y(n_364) );
INVx1_ASAP7_75t_L g383 ( .A(n_312), .Y(n_383) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVxp67_ASAP7_75t_L g327 ( .A(n_315), .Y(n_327) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_315), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_325), .B1(n_330), .B2(n_333), .Y(n_316) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_324), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g393 ( .A(n_326), .Y(n_393) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI221x1_ASAP7_75t_L g379 ( .A1(n_328), .A2(n_380), .B1(n_384), .B2(n_386), .C(n_390), .Y(n_379) );
BUFx2_ASAP7_75t_L g482 ( .A(n_329), .Y(n_482) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_332), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_332), .B(n_409), .Y(n_434) );
AND2x2_ASAP7_75t_L g488 ( .A(n_332), .B(n_367), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_338), .Y(n_333) );
AOI211xp5_ASAP7_75t_L g470 ( .A1(n_335), .A2(n_471), .B(n_477), .C(n_480), .Y(n_470) );
OAI222xp33_ASAP7_75t_L g458 ( .A1(n_336), .A2(n_459), .B1(n_461), .B2(n_462), .C1(n_463), .C2(n_467), .Y(n_458) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AO21x1_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_347), .B(n_348), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_344), .B2(n_345), .Y(n_341) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g484 ( .A(n_347), .Y(n_484) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x2_ASAP7_75t_L g385 ( .A(n_352), .B(n_371), .Y(n_385) );
INVx1_ASAP7_75t_L g411 ( .A(n_352), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_353), .A2(n_407), .B1(n_410), .B2(n_411), .Y(n_406) );
INVx1_ASAP7_75t_L g437 ( .A(n_353), .Y(n_437) );
OR2x6_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g483 ( .A(n_354), .Y(n_483) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g444 ( .A(n_357), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_357), .B(n_373), .Y(n_478) );
OAI21xp33_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_362), .B(n_368), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NOR3x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .C(n_366), .Y(n_363) );
BUFx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B1(n_374), .B2(n_375), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_371), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g456 ( .A(n_371), .Y(n_456) );
INVx2_ASAP7_75t_L g430 ( .A(n_374), .Y(n_430) );
INVx3_ASAP7_75t_L g391 ( .A(n_375), .Y(n_391) );
NOR2x1_ASAP7_75t_L g377 ( .A(n_378), .B(n_435), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_399), .C(n_424), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g447 ( .A(n_396), .Y(n_447) );
BUFx2_ASAP7_75t_L g418 ( .A(n_398), .Y(n_418) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_403), .B(n_406), .C(n_412), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_409), .B(n_476), .Y(n_475) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_416), .B1(n_420), .B2(n_421), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
AND2x2_ASAP7_75t_L g464 ( .A(n_417), .B(n_455), .Y(n_464) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g465 ( .A(n_418), .B(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_441), .C(n_470), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_458), .Y(n_441) );
OAI22xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_446), .B1(n_451), .B2(n_452), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NOR2xp67_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .Y(n_452) );
INVx2_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx2_ASAP7_75t_L g479 ( .A(n_465), .Y(n_479) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI21xp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_485), .B(n_487), .Y(n_480) );
NAND3x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .C(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR2x1_ASAP7_75t_R g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g508 ( .A(n_502), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_502), .B(n_833), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_512), .B(n_521), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_505), .A2(n_522), .B(n_828), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_506), .B(n_838), .Y(n_837) );
INVx5_ASAP7_75t_L g838 ( .A(n_507), .Y(n_838) );
AND2x6_ASAP7_75t_SL g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND3xp33_ASAP7_75t_SL g836 ( .A(n_513), .B(n_522), .C(n_837), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx4_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx12f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
BUFx8_ASAP7_75t_SL g827 ( .A(n_519), .Y(n_827) );
AND2x2_ASAP7_75t_L g834 ( .A(n_519), .B(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g852 ( .A(n_520), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_827), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_730), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_525), .B(n_654), .C(n_685), .D(n_714), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_621), .Y(n_525) );
OAI322xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_565), .A3(n_588), .B1(n_599), .B2(n_607), .C1(n_616), .C2(n_618), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_528), .B(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_541), .Y(n_528) );
AND2x2_ASAP7_75t_L g651 ( .A(n_529), .B(n_652), .Y(n_651) );
INVx4_ASAP7_75t_L g687 ( .A(n_529), .Y(n_687) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g662 ( .A(n_530), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g665 ( .A(n_530), .B(n_567), .Y(n_665) );
AND2x2_ASAP7_75t_L g682 ( .A(n_530), .B(n_579), .Y(n_682) );
AND2x2_ASAP7_75t_L g780 ( .A(n_530), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g603 ( .A(n_531), .Y(n_603) );
AND2x4_ASAP7_75t_L g786 ( .A(n_531), .B(n_781), .Y(n_786) );
AO31x2_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .A3(n_538), .B(n_539), .Y(n_531) );
AO31x2_ASAP7_75t_L g610 ( .A1(n_532), .A2(n_575), .A3(n_611), .B(n_614), .Y(n_610) );
AO31x2_ASAP7_75t_L g629 ( .A1(n_538), .A2(n_596), .A3(n_630), .B(n_633), .Y(n_629) );
AND2x4_ASAP7_75t_L g791 ( .A(n_541), .B(n_692), .Y(n_791) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g620 ( .A(n_542), .Y(n_620) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_542), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_557), .Y(n_542) );
AND2x2_ASAP7_75t_L g608 ( .A(n_543), .B(n_558), .Y(n_608) );
INVx1_ASAP7_75t_L g649 ( .A(n_543), .Y(n_649) );
OAI21x1_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B(n_556), .Y(n_543) );
OAI21x1_ASAP7_75t_L g644 ( .A1(n_544), .A2(n_545), .B(n_556), .Y(n_644) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_550), .B(n_554), .Y(n_545) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g596 ( .A(n_555), .Y(n_596) );
INVx2_ASAP7_75t_L g640 ( .A(n_557), .Y(n_640) );
AND2x2_ASAP7_75t_L g704 ( .A(n_557), .B(n_643), .Y(n_704) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g658 ( .A(n_558), .Y(n_658) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_558), .Y(n_711) );
OR2x2_ASAP7_75t_L g782 ( .A(n_558), .B(n_590), .Y(n_782) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_565), .B(n_661), .C(n_664), .D(n_666), .Y(n_660) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g798 ( .A(n_566), .B(n_786), .Y(n_798) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_578), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_567), .B(n_627), .Y(n_626) );
AND2x4_ASAP7_75t_L g652 ( .A(n_567), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g672 ( .A(n_567), .Y(n_672) );
INVx1_ASAP7_75t_L g689 ( .A(n_567), .Y(n_689) );
INVx1_ASAP7_75t_L g697 ( .A(n_567), .Y(n_697) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_567), .Y(n_811) );
INVx4_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_568), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g729 ( .A(n_568), .B(n_629), .Y(n_729) );
AND2x2_ASAP7_75t_L g737 ( .A(n_568), .B(n_579), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_568), .B(n_760), .Y(n_759) );
BUFx2_ASAP7_75t_L g802 ( .A(n_568), .Y(n_802) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g606 ( .A(n_579), .Y(n_606) );
OR2x2_ASAP7_75t_L g667 ( .A(n_579), .B(n_629), .Y(n_667) );
INVx2_ASAP7_75t_L g674 ( .A(n_579), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_579), .B(n_627), .Y(n_698) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_579), .Y(n_785) );
AO31x2_ASAP7_75t_L g590 ( .A1(n_585), .A2(n_591), .A3(n_596), .B(n_597), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_588), .B(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g609 ( .A(n_590), .B(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g619 ( .A(n_590), .Y(n_619) );
INVx2_ASAP7_75t_L g637 ( .A(n_590), .Y(n_637) );
AND2x4_ASAP7_75t_L g669 ( .A(n_590), .B(n_641), .Y(n_669) );
OR2x2_ASAP7_75t_L g749 ( .A(n_590), .B(n_649), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_604), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_601), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g666 ( .A(n_601), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_601), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_602), .B(n_672), .Y(n_680) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g625 ( .A(n_603), .Y(n_625) );
OR2x2_ASAP7_75t_L g718 ( .A(n_603), .B(n_628), .Y(n_718) );
INVx1_ASAP7_75t_L g645 ( .A(n_604), .Y(n_645) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g617 ( .A(n_605), .Y(n_617) );
INVx1_ASAP7_75t_L g653 ( .A(n_606), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
OAI322xp33_ASAP7_75t_L g621 ( .A1(n_608), .A2(n_622), .A3(n_635), .B1(n_638), .B2(n_645), .C1(n_646), .C2(n_650), .Y(n_621) );
AND2x4_ASAP7_75t_L g668 ( .A(n_608), .B(n_669), .Y(n_668) );
AOI211xp5_ASAP7_75t_SL g699 ( .A1(n_608), .A2(n_700), .B(n_701), .C(n_705), .Y(n_699) );
AND2x2_ASAP7_75t_L g719 ( .A(n_608), .B(n_609), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_608), .B(n_636), .Y(n_725) );
AND2x4_ASAP7_75t_SL g647 ( .A(n_609), .B(n_648), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_609), .B(n_665), .C(n_693), .Y(n_738) );
AND2x2_ASAP7_75t_L g769 ( .A(n_609), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g636 ( .A(n_610), .B(n_637), .Y(n_636) );
INVx3_ASAP7_75t_L g641 ( .A(n_610), .Y(n_641) );
BUFx2_ASAP7_75t_L g709 ( .A(n_610), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_619), .B(n_643), .Y(n_642) );
NAND2x1_ASAP7_75t_L g683 ( .A(n_619), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g702 ( .A(n_619), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_620), .B(n_636), .Y(n_767) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g710 ( .A(n_625), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_629), .Y(n_663) );
AND2x4_ASAP7_75t_L g673 ( .A(n_629), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g760 ( .A(n_629), .Y(n_760) );
INVx2_ASAP7_75t_L g781 ( .A(n_629), .Y(n_781) );
OAI22xp33_ASAP7_75t_L g793 ( .A1(n_635), .A2(n_794), .B1(n_796), .B2(n_797), .Y(n_793) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g705 ( .A(n_636), .B(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g659 ( .A(n_637), .B(n_643), .Y(n_659) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .Y(n_638) );
INVx1_ASAP7_75t_L g678 ( .A(n_639), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x4_ASAP7_75t_L g648 ( .A(n_640), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g770 ( .A(n_640), .Y(n_770) );
INVx2_ASAP7_75t_L g656 ( .A(n_641), .Y(n_656) );
AND2x2_ASAP7_75t_L g684 ( .A(n_641), .B(n_643), .Y(n_684) );
INVx3_ASAP7_75t_L g692 ( .A(n_641), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_641), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g677 ( .A(n_642), .Y(n_677) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g693 ( .A(n_644), .Y(n_693) );
OAI222xp33_ASAP7_75t_L g816 ( .A1(n_646), .A2(n_806), .B1(n_817), .B2(n_820), .C1(n_822), .C2(n_824), .Y(n_816) );
INVx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g757 ( .A(n_648), .Y(n_757) );
AND2x2_ASAP7_75t_L g821 ( .A(n_648), .B(n_691), .Y(n_821) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_651), .B(n_742), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_660), .B1(n_668), .B2(n_670), .C(n_675), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g743 ( .A(n_656), .Y(n_743) );
INVx2_ASAP7_75t_L g805 ( .A(n_657), .Y(n_805) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_L g706 ( .A(n_658), .Y(n_706) );
AND2x2_ASAP7_75t_L g742 ( .A(n_658), .B(n_743), .Y(n_742) );
AND2x4_ASAP7_75t_L g708 ( .A(n_659), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g734 ( .A(n_659), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g823 ( .A(n_659), .Y(n_823) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g772 ( .A(n_663), .Y(n_772) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g795 ( .A(n_665), .B(n_673), .Y(n_795) );
AND2x2_ASAP7_75t_L g818 ( .A(n_665), .B(n_819), .Y(n_818) );
OR2x2_ASAP7_75t_L g679 ( .A(n_667), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g814 ( .A(n_667), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_668), .A2(n_722), .B1(n_756), .B2(n_758), .Y(n_755) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_668), .A2(n_784), .B(n_787), .Y(n_783) );
INVxp67_ASAP7_75t_L g700 ( .A(n_669), .Y(n_700) );
INVx2_ASAP7_75t_SL g804 ( .A(n_669), .Y(n_804) );
AND2x4_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
OR2x2_ASAP7_75t_L g717 ( .A(n_671), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g815 ( .A(n_671), .B(n_814), .Y(n_815) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g688 ( .A(n_673), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_673), .B(n_697), .Y(n_713) );
INVx2_ASAP7_75t_L g740 ( .A(n_673), .Y(n_740) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B1(n_681), .B2(n_683), .Y(n_675) );
NOR2xp33_ASAP7_75t_SL g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_677), .A2(n_751), .B1(n_764), .B2(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g773 ( .A(n_682), .B(n_774), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_690), .B(n_694), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_L g754 ( .A(n_687), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_687), .B(n_737), .Y(n_765) );
INVx1_ASAP7_75t_L g723 ( .A(n_689), .Y(n_723) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_691), .B(n_704), .Y(n_796) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI21xp33_ASAP7_75t_L g809 ( .A1(n_692), .A2(n_810), .B(n_812), .Y(n_809) );
OAI21xp5_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_699), .B(n_707), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g753 ( .A(n_698), .Y(n_753) );
INVx1_ASAP7_75t_L g819 ( .A(n_698), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g792 ( .A(n_702), .Y(n_792) );
OR2x2_ASAP7_75t_L g803 ( .A(n_703), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .C(n_712), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_708), .A2(n_769), .B1(n_771), .B2(n_773), .Y(n_768) );
INVx1_ASAP7_75t_L g735 ( .A(n_709), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_710), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g748 ( .A(n_711), .Y(n_748) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_713), .B(n_717), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_713), .A2(n_776), .B1(n_779), .B2(n_782), .C(n_783), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_719), .B(n_720), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g724 ( .A(n_718), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_725), .B1(n_726), .B2(n_855), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x4_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
AND2x4_ASAP7_75t_L g807 ( .A(n_729), .B(n_785), .Y(n_807) );
NAND4xp25_ASAP7_75t_L g730 ( .A(n_731), .B(n_761), .C(n_788), .D(n_808), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_744), .Y(n_731) );
OAI221xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_736), .B1(n_738), .B2(n_739), .C(n_741), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_734), .A2(n_791), .B1(n_813), .B2(n_815), .Y(n_812) );
INVx1_ASAP7_75t_L g787 ( .A(n_736), .Y(n_787) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g771 ( .A(n_737), .B(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_737), .B(n_780), .Y(n_779) );
NAND2x1_ASAP7_75t_L g824 ( .A(n_737), .B(n_825), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_739), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g746 ( .A(n_743), .B(n_747), .Y(n_746) );
OAI21xp33_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_750), .B(n_755), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g774 ( .A(n_760), .Y(n_774) );
AOI211xp5_ASAP7_75t_L g788 ( .A1(n_760), .A2(n_789), .B(n_793), .C(n_799), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_775), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_763), .B(n_768), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OR2x2_ASAP7_75t_L g822 ( .A(n_770), .B(n_823), .Y(n_822) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AND2x4_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx3_ASAP7_75t_L g826 ( .A(n_786), .Y(n_826) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND2x1p5_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI22xp33_ASAP7_75t_R g799 ( .A1(n_800), .A2(n_803), .B1(n_805), .B2(n_806), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AND2x4_ASAP7_75t_L g813 ( .A(n_802), .B(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_816), .Y(n_808) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx10_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_841), .B(n_846), .Y(n_840) );
OR2x6_ASAP7_75t_L g853 ( .A(n_841), .B(n_846), .Y(n_853) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
INVxp33_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NOR3xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_851), .C(n_852), .Y(n_847) );
INVx2_ASAP7_75t_SL g848 ( .A(n_849), .Y(n_848) );
endmodule