module fake_aes_7195_n_692 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_692, n_648);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_692;
output n_648;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g80 ( .A(n_31), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_7), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_53), .Y(n_82) );
INVxp33_ASAP7_75t_L g83 ( .A(n_61), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_2), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_13), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_79), .Y(n_86) );
CKINVDCx14_ASAP7_75t_R g87 ( .A(n_59), .Y(n_87) );
CKINVDCx16_ASAP7_75t_R g88 ( .A(n_7), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_72), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_65), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_66), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_62), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_56), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_25), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_19), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_67), .Y(n_97) );
INVx4_ASAP7_75t_R g98 ( .A(n_30), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_60), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_36), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_9), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_76), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_27), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_9), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_11), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_16), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_46), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_55), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_40), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_16), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_57), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_14), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_0), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_68), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_1), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_11), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_35), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_48), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_42), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_3), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_78), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_33), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_54), .Y(n_126) );
INVxp33_ASAP7_75t_SL g127 ( .A(n_64), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_26), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_21), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_91), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_90), .A2(n_34), .B(n_75), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_93), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_92), .B(n_0), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_126), .B(n_1), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_104), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_105), .B(n_3), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_94), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_129), .B(n_4), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_88), .B(n_4), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_94), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_122), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_122), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_125), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_101), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_82), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_85), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_83), .B(n_5), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_125), .B(n_5), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_84), .B(n_6), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_99), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_103), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_107), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_110), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_123), .B(n_6), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_111), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_125), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_113), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_125), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_125), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_96), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_117), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_96), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_112), .B(n_114), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_112), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_101), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_132), .B(n_108), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_153), .B(n_114), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_169), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_153), .B(n_119), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_169), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_140), .B(n_105), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
NAND2xp33_ASAP7_75t_L g182 ( .A(n_131), .B(n_97), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_133), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
OR2x2_ASAP7_75t_L g185 ( .A(n_132), .B(n_119), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_154), .B(n_86), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_169), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_140), .B(n_115), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_172), .B(n_86), .Y(n_190) );
OR2x6_ASAP7_75t_L g191 ( .A(n_145), .B(n_115), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_136), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_152), .B(n_100), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
OAI221xp5_ASAP7_75t_L g196 ( .A1(n_139), .A2(n_106), .B1(n_109), .B2(n_118), .C(n_89), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g197 ( .A(n_173), .B(n_102), .Y(n_197) );
INVxp67_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
AO22x2_ASAP7_75t_L g199 ( .A1(n_131), .A2(n_128), .B1(n_120), .B2(n_121), .Y(n_199) );
AO22x2_ASAP7_75t_L g200 ( .A1(n_146), .A2(n_80), .B1(n_124), .B2(n_102), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_169), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_152), .B(n_100), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_141), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_158), .B(n_97), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_158), .B(n_87), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_171), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_151), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_137), .B(n_101), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_146), .A2(n_127), .B1(n_101), .B2(n_116), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_171), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_155), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_159), .B(n_101), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_151), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_159), .B(n_127), .Y(n_218) );
BUFx10_ASAP7_75t_L g219 ( .A(n_143), .Y(n_219) );
INVx4_ASAP7_75t_L g220 ( .A(n_142), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_133), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_151), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_148), .B(n_8), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_151), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_148), .B(n_8), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_174), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_149), .B(n_98), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_174), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_149), .B(n_41), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_160), .B(n_10), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_160), .B(n_10), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_161), .B(n_43), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_161), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_174), .Y(n_234) );
INVx5_ASAP7_75t_L g235 ( .A(n_133), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_162), .B(n_12), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_162), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_164), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_133), .Y(n_239) );
OR2x6_ASAP7_75t_L g240 ( .A(n_138), .B(n_12), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_223), .Y(n_241) );
AND2x6_ASAP7_75t_L g242 ( .A(n_184), .B(n_170), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_175), .Y(n_243) );
OR2x4_ASAP7_75t_L g244 ( .A(n_185), .B(n_157), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_218), .B(n_170), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_223), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_215), .B(n_166), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_215), .B(n_166), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_240), .B(n_163), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_190), .B(n_215), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_223), .B(n_156), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_176), .B(n_164), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_194), .B(n_174), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_198), .B(n_135), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_240), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_240), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_210), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_204), .B(n_135), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_210), .Y(n_260) );
NOR2x1p5_ASAP7_75t_L g261 ( .A(n_178), .B(n_13), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_225), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_200), .A2(n_168), .B1(n_167), .B2(n_130), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_191), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_225), .A2(n_168), .B1(n_167), .B2(n_130), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_230), .Y(n_266) );
BUFx4f_ASAP7_75t_L g267 ( .A(n_230), .Y(n_267) );
BUFx2_ASAP7_75t_SL g268 ( .A(n_225), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_187), .B(n_168), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_213), .A2(n_167), .B1(n_144), .B2(n_147), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_191), .B(n_15), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_216), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_206), .B(n_147), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_207), .B(n_147), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_202), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_233), .B(n_144), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_177), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_230), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
AND3x1_ASAP7_75t_SL g280 ( .A(n_196), .B(n_15), .C(n_17), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_191), .B(n_17), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_237), .B(n_144), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_180), .B(n_18), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_177), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_179), .Y(n_286) );
CKINVDCx6p67_ASAP7_75t_R g287 ( .A(n_219), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_238), .B(n_134), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_220), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_220), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_180), .B(n_18), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_179), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_186), .B(n_165), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_192), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_193), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_188), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_201), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_188), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_203), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_208), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_205), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_208), .Y(n_302) );
INVx4_ASAP7_75t_L g303 ( .A(n_180), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_189), .B(n_134), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_189), .B(n_165), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_211), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_208), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_182), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_189), .B(n_134), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_199), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
BUFx12f_ASAP7_75t_L g312 ( .A(n_257), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
INVx8_ASAP7_75t_L g314 ( .A(n_271), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_258), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_246), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_247), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_287), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_247), .B(n_200), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_249), .B(n_200), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_248), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_267), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_251), .A2(n_231), .B(n_236), .C(n_212), .Y(n_326) );
NAND2xp33_ASAP7_75t_L g327 ( .A(n_242), .B(n_213), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_249), .B(n_182), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_249), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_294), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_253), .B(n_199), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_271), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_283), .B(n_227), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_258), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_259), .A2(n_227), .B(n_229), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_248), .B(n_197), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_271), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_244), .B(n_219), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_264), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_267), .B(n_214), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_294), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_283), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_283), .Y(n_345) );
XOR2xp5_ASAP7_75t_L g346 ( .A(n_264), .B(n_199), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_294), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_310), .A2(n_214), .B1(n_232), .B2(n_229), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_291), .A2(n_214), .B1(n_232), .B2(n_219), .Y(n_349) );
AOI21x1_ASAP7_75t_L g350 ( .A1(n_293), .A2(n_217), .B(n_209), .Y(n_350) );
INVx4_ASAP7_75t_L g351 ( .A(n_291), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_255), .A2(n_195), .B(n_192), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_289), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_250), .A2(n_192), .B(n_195), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_295), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_297), .Y(n_356) );
NOR2x1_ASAP7_75t_R g357 ( .A(n_257), .B(n_195), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_246), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_260), .Y(n_359) );
INVx4_ASAP7_75t_L g360 ( .A(n_291), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_303), .Y(n_361) );
NAND2xp33_ASAP7_75t_L g362 ( .A(n_242), .B(n_224), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_256), .B(n_224), .Y(n_363) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_250), .A2(n_224), .B(n_228), .Y(n_364) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_246), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_314), .A2(n_250), .B1(n_243), .B2(n_281), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_314), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_315), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_314), .Y(n_370) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_346), .A2(n_263), .B(n_245), .C(n_251), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_314), .A2(n_268), .B1(n_303), .B2(n_266), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_323), .B(n_266), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_327), .A2(n_303), .B1(n_262), .B2(n_278), .Y(n_374) );
BUFx10_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_315), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_355), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_332), .B(n_244), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_327), .A2(n_262), .B1(n_242), .B2(n_241), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g380 ( .A1(n_318), .A2(n_242), .B1(n_246), .B2(n_308), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_311), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_337), .A2(n_273), .B(n_265), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_350), .A2(n_265), .B(n_274), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_356), .Y(n_384) );
INVx6_ASAP7_75t_L g385 ( .A(n_311), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_336), .Y(n_386) );
NAND2xp33_ASAP7_75t_L g387 ( .A(n_344), .B(n_242), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_319), .B(n_272), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
OR2x6_ASAP7_75t_L g390 ( .A(n_351), .B(n_252), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_322), .B(n_289), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_351), .A2(n_252), .B1(n_299), .B2(n_306), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_351), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_330), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_360), .B(n_301), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_360), .A2(n_269), .B1(n_261), .B2(n_304), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_313), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_311), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_336), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g400 ( .A1(n_377), .A2(n_338), .B1(n_340), .B2(n_339), .C1(n_341), .C2(n_312), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_377), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_396), .A2(n_340), .B1(n_334), .B2(n_360), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_396), .A2(n_318), .B1(n_312), .B2(n_345), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g404 ( .A1(n_371), .A2(n_334), .B(n_349), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_378), .A2(n_334), .B1(n_328), .B2(n_329), .Y(n_405) );
BUFx4f_ASAP7_75t_SL g406 ( .A(n_367), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_366), .A2(n_326), .B1(n_349), .B2(n_317), .C(n_325), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_395), .A2(n_363), .B1(n_325), .B2(n_364), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_369), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_367), .A2(n_362), .B1(n_342), .B2(n_320), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_395), .A2(n_361), .B1(n_269), .B2(n_362), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_395), .A2(n_361), .B1(n_354), .B2(n_353), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_384), .A2(n_326), .B1(n_270), .B2(n_352), .C(n_254), .Y(n_414) );
BUFx4f_ASAP7_75t_SL g415 ( .A(n_367), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_373), .A2(n_342), .B1(n_361), .B2(n_280), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_395), .A2(n_353), .B1(n_320), .B2(n_324), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_380), .A2(n_348), .B1(n_359), .B2(n_321), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_388), .A2(n_348), .B1(n_321), .B2(n_359), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_384), .A2(n_309), .B1(n_305), .B2(n_282), .C(n_288), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_394), .A2(n_305), .B1(n_276), .B2(n_280), .C(n_316), .Y(n_421) );
BUFx12f_ASAP7_75t_L g422 ( .A(n_370), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_374), .A2(n_324), .B1(n_365), .B2(n_358), .Y(n_423) );
OAI211xp5_ASAP7_75t_L g424 ( .A1(n_389), .A2(n_293), .B(n_324), .C(n_130), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_393), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_379), .A2(n_321), .B1(n_358), .B2(n_365), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_394), .B(n_300), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_388), .A2(n_321), .B1(n_358), .B2(n_365), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_416), .A2(n_421), .B1(n_412), .B2(n_405), .C(n_404), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_400), .B(n_397), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_401), .Y(n_431) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_409), .Y(n_432) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_419), .A2(n_383), .B(n_382), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_403), .A2(n_392), .B1(n_387), .B2(n_390), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_409), .B(n_369), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_402), .A2(n_390), .B1(n_370), .B2(n_397), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_401), .B(n_369), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_427), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_406), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_404), .A2(n_372), .B1(n_390), .B2(n_393), .C(n_391), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_427), .B(n_376), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_428), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_407), .A2(n_399), .B1(n_376), .B2(n_386), .C(n_307), .Y(n_444) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_415), .A2(n_390), .B1(n_376), .B2(n_399), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_411), .A2(n_399), .B1(n_386), .B2(n_390), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_408), .A2(n_386), .B1(n_398), .B2(n_368), .C(n_381), .Y(n_447) );
NAND2x1_ASAP7_75t_L g448 ( .A(n_428), .B(n_385), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_422), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_422), .A2(n_375), .B1(n_385), .B2(n_381), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_425), .B(n_368), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_419), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_414), .B(n_375), .Y(n_453) );
OAI21x1_ASAP7_75t_L g454 ( .A1(n_426), .A2(n_383), .B(n_382), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_420), .B(n_375), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_413), .A2(n_375), .B1(n_365), .B2(n_358), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_410), .A2(n_398), .B1(n_385), .B2(n_381), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_417), .A2(n_307), .B1(n_300), .B2(n_302), .C(n_381), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_423), .Y(n_460) );
AOI33xp33_ASAP7_75t_L g461 ( .A1(n_424), .A2(n_226), .A3(n_209), .B1(n_217), .B2(n_222), .B3(n_228), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
OR2x6_ASAP7_75t_L g463 ( .A(n_428), .B(n_398), .Y(n_463) );
AOI33xp33_ASAP7_75t_L g464 ( .A1(n_449), .A2(n_226), .A3(n_234), .B1(n_222), .B2(n_302), .B3(n_292), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_431), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_462), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_463), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_442), .B(n_368), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_434), .A2(n_385), .B1(n_368), .B2(n_347), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_431), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_439), .B(n_385), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_463), .B(n_20), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_442), .B(n_165), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_429), .A2(n_347), .B1(n_343), .B2(n_335), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_433), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_437), .B(n_165), .Y(n_477) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_443), .B(n_347), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_463), .Y(n_479) );
NOR2x1p5_ASAP7_75t_L g480 ( .A(n_448), .B(n_347), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_430), .A2(n_343), .B1(n_335), .B2(n_331), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_435), .B(n_165), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_443), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_432), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_435), .B(n_165), .Y(n_485) );
AND3x2_ASAP7_75t_L g486 ( .A(n_440), .B(n_438), .C(n_456), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_438), .B(n_150), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_452), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_451), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_452), .Y(n_490) );
NAND2x1p5_ASAP7_75t_L g491 ( .A(n_448), .B(n_343), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_455), .B(n_150), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_436), .A2(n_343), .B1(n_335), .B2(n_331), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_455), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_453), .B(n_335), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_451), .B(n_150), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_433), .B(n_150), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_433), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_463), .Y(n_500) );
OAI22xp5_ASAP7_75t_SL g501 ( .A1(n_441), .A2(n_331), .B1(n_23), .B2(n_24), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_445), .B(n_331), .Y(n_503) );
AOI222xp33_ASAP7_75t_L g504 ( .A1(n_444), .A2(n_133), .B1(n_150), .B2(n_260), .C1(n_279), .C2(n_275), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_447), .Y(n_505) );
AOI21xp5_ASAP7_75t_SL g506 ( .A1(n_450), .A2(n_459), .B(n_460), .Y(n_506) );
AOI211xp5_ASAP7_75t_SL g507 ( .A1(n_460), .A2(n_22), .B(n_28), .C(n_29), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_454), .B(n_150), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_457), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_458), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_461), .B(n_133), .Y(n_511) );
AOI222xp33_ASAP7_75t_L g512 ( .A1(n_439), .A2(n_275), .B1(n_279), .B2(n_292), .C1(n_286), .C2(n_298), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_442), .B(n_32), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_462), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_466), .B(n_514), .Y(n_515) );
NAND2xp33_ASAP7_75t_L g516 ( .A(n_501), .B(n_279), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_494), .B(n_465), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_494), .B(n_37), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_467), .B(n_38), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_486), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_470), .B(n_39), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_498), .B(n_183), .C(n_221), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_489), .B(n_44), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_476), .Y(n_525) );
OAI22xp5_ASAP7_75t_SL g526 ( .A1(n_501), .A2(n_45), .B1(n_47), .B2(n_49), .Y(n_526) );
OAI31xp33_ASAP7_75t_L g527 ( .A1(n_510), .A2(n_298), .A3(n_296), .B(n_286), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_488), .B(n_50), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_476), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_471), .A2(n_296), .B1(n_285), .B2(n_277), .C(n_235), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_483), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_484), .B(n_51), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_467), .B(n_52), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_484), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_490), .B(n_63), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_490), .A2(n_234), .B1(n_239), .B2(n_221), .C(n_183), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_492), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_473), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_492), .B(n_69), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_510), .B(n_70), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_467), .B(n_71), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_498), .B(n_74), .Y(n_542) );
NAND4xp25_ASAP7_75t_L g543 ( .A(n_510), .B(n_277), .C(n_285), .D(n_77), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_468), .B(n_235), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_468), .B(n_235), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_500), .B(n_235), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_480), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_467), .B(n_183), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_479), .B(n_221), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_479), .B(n_221), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_475), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_480), .Y(n_554) );
NAND2x1_ASAP7_75t_L g555 ( .A(n_472), .B(n_239), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_513), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_497), .B(n_239), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_472), .A2(n_474), .B1(n_510), .B2(n_506), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_479), .B(n_239), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_505), .B(n_275), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_496), .B(n_275), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_496), .B(n_279), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_495), .B(n_509), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_475), .Y(n_564) );
NAND2x1_ASAP7_75t_L g565 ( .A(n_472), .B(n_481), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_477), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_499), .Y(n_567) );
INVx3_ASAP7_75t_L g568 ( .A(n_555), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_534), .Y(n_569) );
INVxp33_ASAP7_75t_L g570 ( .A(n_565), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_556), .B(n_478), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_525), .B(n_509), .Y(n_572) );
OAI211xp5_ASAP7_75t_SL g573 ( .A1(n_515), .A2(n_506), .B(n_507), .C(n_464), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_563), .B(n_481), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_563), .B(n_525), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_517), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_521), .B(n_472), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_529), .B(n_478), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_529), .B(n_477), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_518), .B(n_482), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_531), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_544), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_537), .B(n_482), .Y(n_583) );
INVxp67_ASAP7_75t_SL g584 ( .A(n_565), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_558), .A2(n_478), .B1(n_493), .B2(n_469), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_537), .B(n_485), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_538), .B(n_485), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_567), .Y(n_588) );
INVx1_ASAP7_75t_SL g589 ( .A(n_545), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_546), .B(n_499), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_549), .B(n_502), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_567), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_549), .B(n_508), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_547), .B(n_508), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_557), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_554), .B(n_502), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_554), .B(n_491), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_566), .B(n_493), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_542), .B(n_512), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_542), .B(n_491), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_543), .B(n_511), .Y(n_601) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_555), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_532), .B(n_512), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_532), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_545), .B(n_491), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_528), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_548), .B(n_503), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_528), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_540), .B(n_507), .C(n_504), .D(n_511), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_553), .B(n_504), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_575), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_568), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_589), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_584), .A2(n_516), .B1(n_526), .B2(n_560), .C(n_527), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_569), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_576), .Y(n_616) );
AOI31xp33_ASAP7_75t_SL g617 ( .A1(n_577), .A2(n_524), .A3(n_516), .B(n_564), .Y(n_617) );
XOR2x2_ASAP7_75t_L g618 ( .A(n_577), .B(n_541), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_588), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_573), .B(n_524), .Y(n_620) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_605), .B(n_587), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_581), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_588), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_595), .B(n_523), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_584), .A2(n_539), .B(n_548), .C(n_530), .Y(n_625) );
XOR2x2_ASAP7_75t_L g626 ( .A(n_601), .B(n_541), .Y(n_626) );
OAI32xp33_ASAP7_75t_L g627 ( .A1(n_570), .A2(n_539), .A3(n_522), .B1(n_519), .B2(n_535), .Y(n_627) );
AOI221xp5_ASAP7_75t_SL g628 ( .A1(n_585), .A2(n_522), .B1(n_519), .B2(n_559), .C(n_552), .Y(n_628) );
XOR2x2_ASAP7_75t_L g629 ( .A(n_601), .B(n_520), .Y(n_629) );
XOR2x2_ASAP7_75t_L g630 ( .A(n_599), .B(n_520), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g631 ( .A1(n_604), .A2(n_520), .B1(n_533), .B2(n_541), .C1(n_551), .C2(n_552), .Y(n_631) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_568), .B(n_533), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_600), .Y(n_633) );
BUFx3_ASAP7_75t_L g634 ( .A(n_593), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_570), .A2(n_533), .B1(n_559), .B2(n_550), .C(n_561), .Y(n_635) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_592), .Y(n_636) );
INVx3_ASAP7_75t_L g637 ( .A(n_591), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_591), .A2(n_550), .B(n_561), .Y(n_638) );
AOI211xp5_ASAP7_75t_SL g639 ( .A1(n_602), .A2(n_536), .B(n_562), .C(n_573), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_592), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_590), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g642 ( .A1(n_603), .A2(n_562), .B1(n_608), .B2(n_606), .C1(n_598), .C2(n_607), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_572), .Y(n_643) );
XNOR2x1_ASAP7_75t_L g644 ( .A(n_571), .B(n_594), .Y(n_644) );
INVxp67_ASAP7_75t_SL g645 ( .A(n_602), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_609), .A2(n_574), .B(n_597), .C(n_596), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_596), .B(n_579), .Y(n_647) );
UNKNOWN g648 ( );
AOI32xp33_ASAP7_75t_L g649 ( .A1(n_578), .A2(n_596), .A3(n_610), .B1(n_586), .B2(n_580), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_601), .A2(n_558), .B1(n_577), .B2(n_439), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_582), .Y(n_651) );
OAI21xp33_ASAP7_75t_L g652 ( .A1(n_570), .A2(n_584), .B(n_521), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_575), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_568), .B(n_521), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_577), .B(n_515), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_642), .B(n_646), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_623), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_623), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_641), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_647), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_655), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_649), .B(n_639), .C(n_620), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_619), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_626), .A2(n_629), .B1(n_630), .B2(n_620), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_652), .A2(n_654), .B(n_634), .C(n_628), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_626), .A2(n_629), .B1(n_630), .B2(n_650), .Y(n_666) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_614), .B(n_625), .C(n_645), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_643), .B(n_619), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_645), .A2(n_624), .B(n_640), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_667), .B(n_616), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_668), .Y(n_671) );
AOI221x1_ASAP7_75t_L g672 ( .A1(n_662), .A2(n_612), .B1(n_615), .B2(n_637), .C(n_638), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_656), .B(n_636), .Y(n_673) );
NOR3xp33_ASAP7_75t_L g674 ( .A(n_665), .B(n_612), .C(n_635), .Y(n_674) );
XOR2xp5_ASAP7_75t_L g675 ( .A(n_666), .B(n_618), .Y(n_675) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_664), .A2(n_631), .B(n_635), .C(n_627), .Y(n_676) );
NOR5xp2_ASAP7_75t_L g677 ( .A(n_669), .B(n_648), .C(n_653), .D(n_611), .E(n_617), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_674), .B(n_673), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_672), .B(n_669), .C(n_632), .D(n_661), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_671), .B(n_659), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_676), .B(n_658), .C(n_657), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_675), .A2(n_660), .B1(n_618), .B2(n_663), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_680), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_682), .A2(n_670), .B1(n_651), .B2(n_613), .Y(n_684) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_681), .Y(n_685) );
OR2x2_ASAP7_75t_SL g686 ( .A(n_683), .B(n_678), .Y(n_686) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_684), .B(n_679), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_687), .B(n_685), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_686), .A2(n_637), .B1(n_612), .B2(n_644), .Y(n_689) );
XOR2xp5_ASAP7_75t_L g690 ( .A(n_689), .B(n_621), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_690), .A2(n_688), .B1(n_677), .B2(n_633), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_691), .A2(n_647), .B(n_622), .Y(n_692) );
endmodule