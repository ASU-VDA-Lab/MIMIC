module fake_jpeg_2029_n_23 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_2),
.B(n_4),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_6),
.B(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_SL g10 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_10)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_7),
.B1(n_8),
.B2(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_10),
.B(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_15),
.Y(n_16)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_13),
.C(n_11),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_19),
.B(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_18),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_3),
.C(n_4),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_5),
.C(n_0),
.Y(n_23)
);


endmodule