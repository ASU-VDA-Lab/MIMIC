module fake_jpeg_13229_n_135 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_5),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_28),
.B(n_32),
.Y(n_68)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_7),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_51),
.B1(n_22),
.B2(n_25),
.Y(n_62)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_48),
.Y(n_67)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_1),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_63),
.C(n_64),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_22),
.B(n_11),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_11),
.C(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_13),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_68),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_16),
.B(n_1),
.C(n_3),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_75),
.B1(n_39),
.B2(n_41),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_30),
.A2(n_3),
.B1(n_16),
.B2(n_27),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_3),
.B1(n_29),
.B2(n_44),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_76),
.A2(n_33),
.B1(n_36),
.B2(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_82),
.B1(n_79),
.B2(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_67),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_65),
.B1(n_74),
.B2(n_56),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_76),
.B(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_52),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_77),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_80),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_100),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_78),
.B1(n_61),
.B2(n_90),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_53),
.C(n_57),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_96),
.B1(n_105),
.B2(n_85),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_61),
.B1(n_53),
.B2(n_60),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_60),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_114),
.B1(n_105),
.B2(n_100),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_110),
.B(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_98),
.C(n_99),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_102),
.B1(n_101),
.B2(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_120),
.Y(n_121)
);

NOR2xp67_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_111),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_120),
.C(n_118),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_95),
.B(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_117),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_129),
.B(n_130),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_119),
.A3(n_121),
.B1(n_122),
.B2(n_115),
.C1(n_114),
.C2(n_94),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_98),
.B(n_58),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_131),
.C(n_58),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_60),
.Y(n_135)
);


endmodule