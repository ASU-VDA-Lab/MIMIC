module real_jpeg_5876_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_1),
.A2(n_23),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_52),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_1),
.A2(n_52),
.B1(n_126),
.B2(n_243),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_1),
.A2(n_52),
.B1(n_269),
.B2(n_272),
.Y(n_268)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_3),
.A2(n_22),
.B1(n_123),
.B2(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_39),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_3),
.A2(n_22),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_3),
.A2(n_22),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_3),
.A2(n_222),
.B(n_224),
.C(n_230),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_3),
.B(n_255),
.C(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_3),
.B(n_97),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_3),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_3),
.B(n_111),
.Y(n_299)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_5),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_5),
.Y(n_158)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_5),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_5),
.Y(n_286)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_6),
.Y(n_135)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_8),
.Y(n_136)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_8),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_8),
.Y(n_199)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_9),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_10),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_10),
.A2(n_88),
.B1(n_150),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_10),
.A2(n_88),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_10),
.A2(n_88),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_11),
.A2(n_144),
.B1(n_145),
.B2(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_11),
.Y(n_144)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_211),
.B1(n_323),
.B2(n_324),
.Y(n_13)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_14),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_210),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_177),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_17),
.B(n_177),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.C(n_161),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_18),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_54),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_19),
.B(n_55),
.C(n_99),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_50),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_24),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_22),
.A2(n_225),
.B(n_227),
.Y(n_224)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_24),
.Y(n_137)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_27),
.B(n_51),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_32),
.Y(n_141)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_39),
.B(n_195),
.Y(n_194)
);

AO22x1_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_42),
.Y(n_139)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_44),
.Y(n_133)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_98),
.B1(n_99),
.B2(n_128),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_91),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_83),
.Y(n_57)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_63),
.Y(n_226)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_66),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_66),
.Y(n_232)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_72),
.Y(n_209)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_73),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_77),
.Y(n_245)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_82),
.Y(n_223)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_84),
.B(n_97),
.Y(n_163)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_91),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_92),
.B(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_120),
.B(n_121),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_101),
.B(n_122),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_101),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_101),
.B(n_185),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_111),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_108),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_112),
.B1(n_114),
.B2(n_118),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_110),
.Y(n_229)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_111),
.B(n_242),
.Y(n_259)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_115),
.Y(n_272)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_119),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_119),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_120),
.B(n_121),
.Y(n_240)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_125),
.Y(n_253)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_129),
.A2(n_130),
.B1(n_161),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_142),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_131),
.B(n_142),
.Y(n_191)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.A3(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_152),
.B(n_154),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_176),
.B(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx8_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_153),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_154),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_155),
.A2(n_170),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_155),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_159),
.Y(n_176)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_165),
.B(n_205),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_169),
.B(n_284),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_170),
.Y(n_265)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_173),
.Y(n_271)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_176),
.B(n_267),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_177),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.CI(n_190),
.CON(n_177),
.SN(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_183),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_184),
.B(n_241),
.Y(n_274)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_201),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_211),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_246),
.B(n_322),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_213),
.B(n_216),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.C(n_237),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_217),
.B(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_220),
.A2(n_237),
.B1(n_238),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_220),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_233),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_221),
.A2(n_233),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_221),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_233),
.Y(n_313)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_316),
.B(n_321),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_303),
.B(n_315),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_278),
.B(n_302),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_260),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_250),
.B(n_260),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_258),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_252),
.B1(n_258),
.B2(n_281),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_273),
.Y(n_260)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

INVx3_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_276),
.C(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_288),
.B(n_301),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_282),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_297),
.B(n_300),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_296),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_306),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_310),
.C(n_312),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_320),
.Y(n_321)
);


endmodule