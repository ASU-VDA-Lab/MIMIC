module real_aes_6271_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_98;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_0), .A2(n_102), .B(n_105), .C(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_1), .A2(n_131), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_2), .B(n_161), .Y(n_160) );
AND2x6_ASAP7_75t_L g102 ( .A(n_3), .B(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g493 ( .A(n_3), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_3), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_4), .A2(n_43), .B1(n_461), .B2(n_465), .Y(n_460) );
INVx1_ASAP7_75t_L g198 ( .A(n_5), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_6), .B(n_114), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_7), .B(n_439), .Y(n_438) );
AO22x2_ASAP7_75t_L g410 ( .A1(n_8), .A2(n_27), .B1(n_411), .B2(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g94 ( .A(n_9), .Y(n_94) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_10), .A2(n_139), .B(n_220), .C(n_222), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_11), .B(n_161), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_12), .A2(n_401), .B1(n_402), .B2(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_12), .Y(n_401) );
AO22x2_ASAP7_75t_L g414 ( .A1(n_13), .A2(n_29), .B1(n_411), .B2(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g444 ( .A1(n_14), .A2(n_46), .B1(n_445), .B2(n_448), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_15), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_16), .A2(n_155), .B(n_206), .C(n_208), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_17), .B(n_114), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_18), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_19), .B(n_114), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_20), .Y(n_96) );
INVx1_ASAP7_75t_L g168 ( .A(n_21), .Y(n_168) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_22), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_23), .Y(n_183) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_24), .A2(n_54), .B1(n_454), .B2(n_458), .Y(n_453) );
INVx1_ASAP7_75t_L g137 ( .A(n_25), .Y(n_137) );
INVx2_ASAP7_75t_L g100 ( .A(n_26), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_28), .Y(n_189) );
OAI221xp5_ASAP7_75t_L g485 ( .A1(n_29), .A2(n_41), .B1(n_53), .B2(n_486), .C(n_487), .Y(n_485) );
INVxp67_ASAP7_75t_L g488 ( .A(n_29), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_30), .A2(n_155), .B(n_156), .C(n_158), .Y(n_154) );
INVxp67_ASAP7_75t_L g140 ( .A(n_31), .Y(n_140) );
CKINVDCx14_ASAP7_75t_R g153 ( .A(n_32), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g166 ( .A1(n_33), .A2(n_105), .B(n_167), .C(n_171), .Y(n_166) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_34), .A2(n_39), .B1(n_423), .B2(n_429), .Y(n_422) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_35), .A2(n_116), .B(n_196), .C(n_197), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_36), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_37), .Y(n_133) );
INVx1_ASAP7_75t_L g204 ( .A(n_38), .Y(n_204) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_40), .Y(n_396) );
AO22x2_ASAP7_75t_L g418 ( .A1(n_41), .A2(n_64), .B1(n_411), .B2(n_415), .Y(n_418) );
INVxp67_ASAP7_75t_L g489 ( .A(n_41), .Y(n_489) );
CKINVDCx14_ASAP7_75t_R g194 ( .A(n_42), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_42), .A2(n_194), .B1(n_394), .B2(n_398), .Y(n_393) );
INVx1_ASAP7_75t_L g103 ( .A(n_44), .Y(n_103) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_45), .Y(n_392) );
INVx1_ASAP7_75t_L g93 ( .A(n_47), .Y(n_93) );
INVx1_ASAP7_75t_SL g157 ( .A(n_48), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_49), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_50), .B(n_161), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_51), .A2(n_71), .B1(n_471), .B2(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
AO22x2_ASAP7_75t_L g420 ( .A1(n_53), .A2(n_70), .B1(n_411), .B2(n_412), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_55), .A2(n_131), .B(n_193), .Y(n_192) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_56), .A2(n_72), .B1(n_477), .B2(n_480), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_57), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_58), .A2(n_131), .B(n_217), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_59), .A2(n_130), .B(n_132), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_60), .Y(n_165) );
INVx1_ASAP7_75t_L g218 ( .A(n_61), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_62), .A2(n_131), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g221 ( .A(n_63), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_65), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g91 ( .A(n_66), .Y(n_91) );
INVx1_ASAP7_75t_L g186 ( .A(n_67), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_68), .A2(n_395), .B1(n_396), .B2(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_68), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g104 ( .A1(n_69), .A2(n_105), .B(n_108), .C(n_118), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_73), .B(n_89), .Y(n_199) );
INVx1_ASAP7_75t_L g411 ( .A(n_74), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_74), .Y(n_413) );
XOR2xp5_ASAP7_75t_L g508 ( .A(n_75), .B(n_402), .Y(n_508) );
INVx2_ASAP7_75t_L g207 ( .A(n_76), .Y(n_207) );
AOI221xp5_ASAP7_75t_SL g77 ( .A1(n_78), .A2(n_384), .B1(n_389), .B2(n_482), .C(n_494), .Y(n_77) );
OR2x2_ASAP7_75t_L g78 ( .A(n_79), .B(n_318), .Y(n_78) );
NAND5xp2_ASAP7_75t_L g79 ( .A(n_80), .B(n_247), .C(n_277), .D(n_298), .E(n_304), .Y(n_79) );
AOI221xp5_ASAP7_75t_SL g80 ( .A1(n_81), .A2(n_177), .B1(n_211), .B2(n_213), .C(n_224), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_174), .Y(n_82) );
NOR2xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_146), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
A2O1A1Ixp33_ASAP7_75t_SL g298 ( .A1(n_85), .A2(n_162), .B(n_299), .C(n_302), .Y(n_298) );
AND2x2_ASAP7_75t_L g368 ( .A(n_85), .B(n_163), .Y(n_368) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_124), .Y(n_85) );
AND2x2_ASAP7_75t_L g226 ( .A(n_86), .B(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g230 ( .A(n_86), .B(n_227), .Y(n_230) );
OR2x2_ASAP7_75t_L g256 ( .A(n_86), .B(n_163), .Y(n_256) );
AND2x2_ASAP7_75t_L g258 ( .A(n_86), .B(n_149), .Y(n_258) );
AND2x2_ASAP7_75t_L g276 ( .A(n_86), .B(n_148), .Y(n_276) );
INVx1_ASAP7_75t_L g309 ( .A(n_86), .Y(n_309) );
INVx2_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
BUFx2_ASAP7_75t_L g176 ( .A(n_87), .Y(n_176) );
AND2x2_ASAP7_75t_L g212 ( .A(n_87), .B(n_149), .Y(n_212) );
AND2x2_ASAP7_75t_L g365 ( .A(n_87), .B(n_163), .Y(n_365) );
AO21x2_ASAP7_75t_L g87 ( .A1(n_88), .A2(n_95), .B(n_120), .Y(n_87) );
INVx3_ASAP7_75t_L g161 ( .A(n_88), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_88), .B(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_88), .B(n_189), .Y(n_188) );
INVx4_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g127 ( .A(n_90), .Y(n_127) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_92), .Y(n_90) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_91), .B(n_92), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g92 ( .A(n_93), .B(n_94), .Y(n_92) );
OAI21xp5_ASAP7_75t_L g95 ( .A1(n_96), .A2(n_97), .B(n_104), .Y(n_95) );
O2A1O1Ixp33_ASAP7_75t_L g164 ( .A1(n_97), .A2(n_123), .B(n_165), .C(n_166), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_97), .A2(n_183), .B(n_184), .Y(n_182) );
NAND2x1p5_ASAP7_75t_L g97 ( .A(n_98), .B(n_102), .Y(n_97) );
AND2x4_ASAP7_75t_L g131 ( .A(n_98), .B(n_102), .Y(n_131) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_101), .Y(n_98) );
INVx1_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g106 ( .A(n_100), .Y(n_106) );
INVx1_ASAP7_75t_L g209 ( .A(n_100), .Y(n_209) );
INVx1_ASAP7_75t_L g107 ( .A(n_101), .Y(n_107) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_101), .Y(n_112) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_101), .Y(n_114) );
INVx3_ASAP7_75t_L g139 ( .A(n_101), .Y(n_139) );
INVx4_ASAP7_75t_SL g119 ( .A(n_102), .Y(n_119) );
BUFx3_ASAP7_75t_L g171 ( .A(n_102), .Y(n_171) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_103), .Y(n_491) );
INVx5_ASAP7_75t_L g134 ( .A(n_105), .Y(n_134) );
AND2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
BUFx3_ASAP7_75t_L g117 ( .A(n_106), .Y(n_117) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_106), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_110), .B(n_113), .C(n_115), .Y(n_108) );
O2A1O1Ixp5_ASAP7_75t_L g185 ( .A1(n_110), .A2(n_115), .B(n_186), .C(n_187), .Y(n_185) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_110), .Y(n_387) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx4_ASAP7_75t_L g141 ( .A(n_112), .Y(n_141) );
INVx4_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
INVx2_ASAP7_75t_L g196 ( .A(n_114), .Y(n_196) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g222 ( .A(n_117), .Y(n_222) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
O2A1O1Ixp33_ASAP7_75t_SL g132 ( .A1(n_119), .A2(n_133), .B(n_134), .C(n_135), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_119), .A2(n_134), .B(n_153), .C(n_154), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_SL g193 ( .A1(n_119), .A2(n_134), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_SL g203 ( .A1(n_119), .A2(n_134), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_SL g217 ( .A1(n_119), .A2(n_134), .B(n_218), .C(n_219), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_119), .B(n_170), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g145 ( .A(n_122), .Y(n_145) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g181 ( .A(n_123), .Y(n_181) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_123), .A2(n_192), .B(n_199), .Y(n_191) );
AND2x2_ASAP7_75t_L g246 ( .A(n_124), .B(n_147), .Y(n_246) );
OR2x2_ASAP7_75t_L g250 ( .A(n_124), .B(n_163), .Y(n_250) );
AND2x2_ASAP7_75t_L g275 ( .A(n_124), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_SL g322 ( .A(n_124), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_124), .B(n_284), .Y(n_370) );
AO21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_128), .B(n_143), .Y(n_124) );
INVx1_ASAP7_75t_L g228 ( .A(n_125), .Y(n_228) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_129), .A2(n_144), .B(n_228), .Y(n_227) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_136), .B(n_142), .Y(n_135) );
OAI22xp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B1(n_140), .B2(n_141), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_138), .A2(n_168), .B(n_169), .C(n_170), .Y(n_167) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_139), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_141), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_141), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI322xp33_ASAP7_75t_L g371 ( .A1(n_146), .A2(n_307), .A3(n_330), .B1(n_351), .B2(n_372), .C1(n_374), .C2(n_375), .Y(n_371) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_147), .B(n_227), .Y(n_374) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_162), .Y(n_147) );
AND2x2_ASAP7_75t_L g175 ( .A(n_148), .B(n_176), .Y(n_175) );
AND2x4_ASAP7_75t_L g243 ( .A(n_148), .B(n_163), .Y(n_243) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g284 ( .A(n_149), .B(n_163), .Y(n_284) );
AND2x2_ASAP7_75t_L g328 ( .A(n_149), .B(n_162), .Y(n_328) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_160), .Y(n_149) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_150), .A2(n_202), .B(n_210), .Y(n_201) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_150), .A2(n_216), .B(n_223), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_155), .B(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g211 ( .A(n_162), .B(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g229 ( .A(n_162), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_162), .B(n_258), .Y(n_382) );
INVx3_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g174 ( .A(n_163), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_163), .B(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g296 ( .A(n_163), .B(n_227), .Y(n_296) );
AND2x2_ASAP7_75t_L g323 ( .A(n_163), .B(n_258), .Y(n_323) );
OR2x2_ASAP7_75t_L g379 ( .A(n_163), .B(n_230), .Y(n_379) );
OR2x6_ASAP7_75t_L g163 ( .A(n_164), .B(n_172), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_170), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_SL g265 ( .A(n_174), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_175), .B(n_296), .Y(n_297) );
AND2x2_ASAP7_75t_L g331 ( .A(n_175), .B(n_321), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_175), .B(n_254), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_175), .B(n_376), .Y(n_375) );
OAI31xp33_ASAP7_75t_L g349 ( .A1(n_177), .A2(n_211), .A3(n_350), .B(n_352), .Y(n_349) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_190), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_178), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g332 ( .A(n_178), .B(n_267), .Y(n_332) );
OR2x2_ASAP7_75t_L g339 ( .A(n_178), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g351 ( .A(n_178), .B(n_240), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
OR2x2_ASAP7_75t_L g285 ( .A(n_179), .B(n_286), .Y(n_285) );
BUFx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g213 ( .A(n_180), .B(n_214), .Y(n_213) );
INVx4_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
AND2x2_ASAP7_75t_L g271 ( .A(n_180), .B(n_215), .Y(n_271) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_188), .Y(n_180) );
AND2x2_ASAP7_75t_L g270 ( .A(n_190), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g340 ( .A(n_190), .Y(n_340) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_200), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_191), .B(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g240 ( .A(n_191), .B(n_201), .Y(n_240) );
INVx2_ASAP7_75t_L g260 ( .A(n_191), .Y(n_260) );
AND2x2_ASAP7_75t_L g274 ( .A(n_191), .B(n_201), .Y(n_274) );
AND2x2_ASAP7_75t_L g281 ( .A(n_191), .B(n_237), .Y(n_281) );
BUFx3_ASAP7_75t_L g291 ( .A(n_191), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_191), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g236 ( .A(n_200), .Y(n_236) );
AND2x2_ASAP7_75t_L g244 ( .A(n_200), .B(n_234), .Y(n_244) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g214 ( .A(n_201), .B(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_SL g251 ( .A(n_212), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_212), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_212), .B(n_321), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_213), .B(n_291), .Y(n_344) );
INVx1_ASAP7_75t_SL g378 ( .A(n_213), .Y(n_378) );
INVx1_ASAP7_75t_SL g286 ( .A(n_214), .Y(n_286) );
INVx1_ASAP7_75t_SL g237 ( .A(n_215), .Y(n_237) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
OR2x2_ASAP7_75t_L g259 ( .A(n_215), .B(n_234), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_215), .B(n_234), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_215), .B(n_263), .Y(n_325) );
INVx1_ASAP7_75t_L g496 ( .A(n_218), .Y(n_496) );
OAI322xp33_ASAP7_75t_L g494 ( .A1(n_221), .A2(n_495), .A3(n_498), .B1(n_502), .B2(n_503), .C1(n_508), .C2(n_509), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_229), .B(n_231), .C(n_242), .Y(n_224) );
AOI31xp33_ASAP7_75t_L g341 ( .A1(n_225), .A2(n_342), .A3(n_343), .B(n_344), .Y(n_341) );
AND2x2_ASAP7_75t_L g314 ( .A(n_226), .B(n_243), .Y(n_314) );
BUFx3_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_227), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g290 ( .A(n_227), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_227), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g245 ( .A(n_230), .Y(n_245) );
OAI222xp33_ASAP7_75t_L g354 ( .A1(n_230), .A2(n_355), .B1(n_358), .B2(n_359), .C1(n_360), .C2(n_361), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
INVx1_ASAP7_75t_L g360 ( .A(n_232), .Y(n_360) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_234), .B(n_237), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_234), .B(n_260), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_234), .B(n_235), .Y(n_330) );
INVx1_ASAP7_75t_L g381 ( .A(n_234), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_235), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g383 ( .A(n_235), .Y(n_383) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_237), .Y(n_306) );
AOI32xp33_ASAP7_75t_L g242 ( .A1(n_238), .A2(n_243), .A3(n_244), .B1(n_245), .B2(n_246), .Y(n_242) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_240), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g317 ( .A(n_240), .Y(n_317) );
OR2x2_ASAP7_75t_L g358 ( .A(n_240), .B(n_259), .Y(n_358) );
INVx1_ASAP7_75t_L g294 ( .A(n_241), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_243), .B(n_254), .Y(n_279) );
INVx3_ASAP7_75t_L g288 ( .A(n_243), .Y(n_288) );
AOI322xp5_ASAP7_75t_L g304 ( .A1(n_243), .A2(n_288), .A3(n_305), .B1(n_307), .B2(n_310), .C1(n_314), .C2(n_315), .Y(n_304) );
AND2x2_ASAP7_75t_L g280 ( .A(n_244), .B(n_281), .Y(n_280) );
INVxp67_ASAP7_75t_L g357 ( .A(n_244), .Y(n_357) );
A2O1A1O1Ixp25_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_252), .C(n_260), .D(n_261), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_248), .B(n_291), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OAI221xp5_ASAP7_75t_L g261 ( .A1(n_250), .A2(n_262), .B1(n_265), .B2(n_266), .C(n_269), .Y(n_261) );
INVx1_ASAP7_75t_SL g376 ( .A(n_250), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .B(n_259), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_254), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI221xp5_ASAP7_75t_SL g346 ( .A1(n_256), .A2(n_340), .B1(n_347), .B2(n_348), .C(n_349), .Y(n_346) );
OAI222xp33_ASAP7_75t_L g377 ( .A1(n_257), .A2(n_378), .B1(n_379), .B2(n_380), .C1(n_382), .C2(n_383), .Y(n_377) );
AND2x2_ASAP7_75t_L g335 ( .A(n_258), .B(n_321), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_258), .A2(n_273), .B(n_320), .Y(n_347) );
INVx1_ASAP7_75t_L g361 ( .A(n_258), .Y(n_361) );
INVx2_ASAP7_75t_SL g264 ( .A(n_259), .Y(n_264) );
AND2x2_ASAP7_75t_L g267 ( .A(n_260), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_SL g301 ( .A(n_263), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_263), .B(n_273), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_264), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_264), .B(n_274), .Y(n_303) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OAI21xp5_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_272), .B(n_275), .Y(n_269) );
INVx1_ASAP7_75t_SL g287 ( .A(n_271), .Y(n_287) );
AND2x2_ASAP7_75t_L g334 ( .A(n_271), .B(n_317), .Y(n_334) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x2_ASAP7_75t_L g373 ( .A(n_273), .B(n_291), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_274), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g359 ( .A(n_275), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B1(n_282), .B2(n_289), .C(n_292), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B1(n_287), .B2(n_288), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_286), .A2(n_293), .B1(n_295), .B2(n_297), .Y(n_292) );
OR2x2_ASAP7_75t_L g363 ( .A(n_287), .B(n_291), .Y(n_363) );
OR2x2_ASAP7_75t_L g366 ( .A(n_287), .B(n_301), .Y(n_366) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_308), .A2(n_363), .B1(n_364), .B2(n_366), .C(n_367), .Y(n_362) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND3xp33_ASAP7_75t_SL g318 ( .A(n_319), .B(n_333), .C(n_345), .Y(n_318) );
AOI222xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_324), .B1(n_326), .B2(n_329), .C1(n_331), .C2(n_332), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_321), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g343 ( .A(n_323), .Y(n_343) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVxp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_336), .B2(n_338), .C(n_341), .Y(n_333) );
INVx1_ASAP7_75t_L g348 ( .A(n_334), .Y(n_348) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_338), .A2(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
NOR5xp2_ASAP7_75t_L g345 ( .A(n_346), .B(n_354), .C(n_362), .D(n_371), .E(n_377), .Y(n_345) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_385), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g506 ( .A(n_387), .Y(n_506) );
XOR2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_400), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_393), .B2(n_399), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_392), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_393), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_394), .Y(n_398) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_SL g495 ( .A1(n_402), .A2(n_403), .B1(n_496), .B2(n_497), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND3x1_ASAP7_75t_L g404 ( .A(n_405), .B(n_452), .C(n_469), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_431), .Y(n_405) );
OAI21xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_421), .B(n_422), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x6_ASAP7_75t_L g408 ( .A(n_409), .B(n_416), .Y(n_408) );
AND2x4_ASAP7_75t_L g449 ( .A(n_409), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_414), .Y(n_409) );
AND2x2_ASAP7_75t_L g428 ( .A(n_410), .B(n_418), .Y(n_428) );
INVx2_ASAP7_75t_L g436 ( .A(n_410), .Y(n_436) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_413), .Y(n_415) );
INVx2_ASAP7_75t_L g427 ( .A(n_414), .Y(n_427) );
AND2x2_ASAP7_75t_L g435 ( .A(n_414), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g443 ( .A(n_414), .B(n_436), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_414), .Y(n_447) );
AND2x2_ASAP7_75t_L g456 ( .A(n_416), .B(n_457), .Y(n_456) );
AND2x6_ASAP7_75t_L g479 ( .A(n_416), .B(n_442), .Y(n_479) );
AND2x4_ASAP7_75t_L g481 ( .A(n_416), .B(n_435), .Y(n_481) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
AND2x2_ASAP7_75t_L g437 ( .A(n_417), .B(n_420), .Y(n_437) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g464 ( .A(n_418), .B(n_451), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_418), .B(n_420), .Y(n_468) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g426 ( .A(n_420), .Y(n_426) );
INVx1_ASAP7_75t_L g451 ( .A(n_420), .Y(n_451) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_426), .Y(n_430) );
AND2x2_ASAP7_75t_L g457 ( .A(n_427), .B(n_436), .Y(n_457) );
AND2x4_ASAP7_75t_L g429 ( .A(n_428), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g445 ( .A(n_428), .B(n_446), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_438), .C(n_444), .Y(n_431) );
BUFx4f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x6_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
AND2x2_ASAP7_75t_L g463 ( .A(n_435), .B(n_464), .Y(n_463) );
AND2x4_ASAP7_75t_L g441 ( .A(n_437), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g459 ( .A(n_437), .B(n_457), .Y(n_459) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx4_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x6_ASAP7_75t_L g467 ( .A(n_447), .B(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_460), .Y(n_452) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g472 ( .A(n_457), .B(n_464), .Y(n_472) );
AND2x4_ASAP7_75t_L g474 ( .A(n_457), .B(n_475), .Y(n_474) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx8_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx6_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g475 ( .A(n_468), .Y(n_475) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .Y(n_469) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx11_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
AND3x1_ASAP7_75t_SL g484 ( .A(n_485), .B(n_490), .C(n_492), .Y(n_484) );
INVxp67_ASAP7_75t_L g501 ( .A(n_485), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_SL g502 ( .A(n_490), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_490), .A2(n_505), .B(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g512 ( .A(n_490), .Y(n_512) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_491), .B(n_493), .Y(n_507) );
OR2x2_ASAP7_75t_SL g511 ( .A(n_492), .B(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_496), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
endmodule