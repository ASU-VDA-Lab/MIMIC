module fake_netlist_6_3569_n_1690 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1690);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1690;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_108),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_37),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_86),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_58),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_43),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_84),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_80),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_8),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_81),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_30),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_144),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_52),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_119),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_55),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_129),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_73),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_52),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

CKINVDCx11_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_56),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_91),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_43),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_100),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_61),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_92),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_146),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_125),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_99),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_23),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_51),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_77),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_0),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_67),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_102),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_94),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_71),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_59),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_64),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_19),
.Y(n_214)
);

INVxp33_ASAP7_75t_R g215 ( 
.A(n_12),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_5),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_82),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_121),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_39),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_90),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_87),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_0),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_72),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_29),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_35),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_135),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_70),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_35),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_48),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_40),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_27),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_50),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_83),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_45),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_4),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_39),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_105),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_112),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_59),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_68),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_63),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_3),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_9),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_48),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_96),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_17),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_56),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_22),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_158),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_24),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_11),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_21),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_154),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_13),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_156),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_142),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_106),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_145),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_44),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_155),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_49),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_46),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_116),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_150),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_75),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_109),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_63),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_104),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_16),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_114),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_58),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_93),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_141),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_132),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_88),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_101),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_64),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_97),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_44),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_20),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_69),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_12),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_30),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_61),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_34),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_53),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_130),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_34),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_1),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_65),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_57),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_98),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_115),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_95),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_128),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_122),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_118),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_41),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_78),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_133),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_137),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_89),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_153),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_38),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_85),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_74),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_24),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_21),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_15),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_20),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_9),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_16),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_57),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_6),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_136),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_140),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_7),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_65),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_49),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_66),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_38),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_13),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_103),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_234),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_191),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_189),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_176),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_161),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_181),
.B(n_1),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_231),
.Y(n_341)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_234),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_162),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_163),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_232),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_166),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_167),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_268),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_181),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g352 ( 
.A(n_270),
.B(n_2),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_254),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_191),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_295),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_236),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_236),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_270),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_168),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_239),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_172),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_182),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_239),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_242),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_184),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_303),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_325),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_165),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_192),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_253),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_253),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_185),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_325),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_195),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_192),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_197),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_198),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_302),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_302),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_326),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_170),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_217),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_171),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_294),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_178),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_294),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_309),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_R g390 ( 
.A(n_199),
.B(n_110),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_202),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_180),
.B(n_2),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_194),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_194),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_207),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_241),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_196),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_196),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_217),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_208),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_210),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_190),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_225),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_204),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_204),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_180),
.B(n_5),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_228),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_238),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_201),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_246),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_206),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_206),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_213),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_164),
.B(n_6),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_262),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_241),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_263),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_271),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_213),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_219),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_219),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_272),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_227),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_274),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_334),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_366),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_334),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_276),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_247),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_339),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_344),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_346),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_366),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_366),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_205),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_392),
.B(n_278),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_345),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_336),
.B(n_355),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_282),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_357),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_338),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_357),
.B(n_242),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_393),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_393),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_352),
.B(n_221),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_348),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_404),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_371),
.B(n_377),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_352),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_349),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_353),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_383),
.B(n_209),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_362),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_341),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_362),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_347),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_221),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_365),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_361),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_411),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_350),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_363),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_368),
.Y(n_482)
);

NOR2x1_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_211),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_353),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_412),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_413),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_365),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_389),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_419),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_419),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_420),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_369),
.B(n_247),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_400),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_364),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_372),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_356),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_367),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_374),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_401),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_420),
.B(n_283),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_372),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_380),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_455),
.B(n_211),
.Y(n_504)
);

BUFx10_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_483),
.B(n_226),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_430),
.B(n_164),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_468),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_468),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_428),
.B(n_376),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_483),
.B(n_226),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_431),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_378),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_440),
.B(n_242),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_445),
.B(n_379),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_445),
.B(n_395),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_442),
.B(n_410),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_449),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_468),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_473),
.A2(n_375),
.B1(n_342),
.B2(n_335),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_452),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_453),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_454),
.Y(n_526)
);

OAI22xp33_ASAP7_75t_L g527 ( 
.A1(n_473),
.A2(n_416),
.B1(n_396),
.B2(n_267),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_430),
.B(n_373),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_454),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_438),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_457),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_455),
.B(n_169),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_455),
.B(n_415),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_455),
.B(n_417),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_475),
.Y(n_536)
);

BUFx8_ASAP7_75t_SL g537 ( 
.A(n_448),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_418),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_R g539 ( 
.A(n_503),
.B(n_337),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_432),
.B(n_422),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

INVx4_ASAP7_75t_SL g542 ( 
.A(n_449),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_460),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_433),
.B(n_373),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_462),
.B(n_169),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_433),
.B(n_424),
.Y(n_547)
);

BUFx4f_ASAP7_75t_L g548 ( 
.A(n_443),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_468),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_463),
.B(n_387),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_466),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_463),
.B(n_311),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_438),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_449),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_501),
.B(n_311),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_493),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_478),
.A2(n_381),
.B1(n_416),
.B2(n_396),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_496),
.Y(n_562)
);

CKINVDCx8_ASAP7_75t_R g563 ( 
.A(n_465),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_501),
.B(n_242),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_434),
.B(n_403),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_473),
.A2(n_493),
.B1(n_320),
.B2(n_249),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_496),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_475),
.B(n_394),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_443),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_496),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_473),
.B(n_402),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_471),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_476),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_443),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_476),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_496),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_479),
.B(n_480),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_484),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_435),
.B(n_407),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_480),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_443),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_473),
.B(n_409),
.Y(n_584)
);

AO21x2_ASAP7_75t_L g585 ( 
.A1(n_467),
.A2(n_177),
.B(n_174),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_456),
.B(n_408),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_496),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_478),
.B(n_356),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_485),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_464),
.B(n_242),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_485),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_481),
.B(n_174),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_465),
.B(n_497),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_496),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_494),
.Y(n_595)
);

BUFx4f_ASAP7_75t_L g596 ( 
.A(n_443),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_495),
.B(n_177),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_486),
.B(n_487),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_498),
.B(n_179),
.Y(n_600)
);

AND3x2_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_299),
.C(n_351),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_499),
.B(n_179),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_489),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_490),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_425),
.B(n_266),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_425),
.B(n_281),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_427),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_447),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_427),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_429),
.B(n_436),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_475),
.B(n_382),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_491),
.B(n_351),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_429),
.Y(n_615)
);

BUFx4f_ASAP7_75t_L g616 ( 
.A(n_447),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_491),
.B(n_360),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_492),
.B(n_360),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_447),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_SL g620 ( 
.A1(n_492),
.A2(n_260),
.B1(n_290),
.B2(n_186),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_461),
.B(n_394),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_436),
.B(n_441),
.Y(n_622)
);

AND3x2_ASAP7_75t_L g623 ( 
.A(n_450),
.B(n_398),
.C(n_188),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_441),
.B(n_284),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_444),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_444),
.B(n_186),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_446),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_447),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_459),
.B(n_386),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_446),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_426),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_459),
.B(n_386),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_459),
.B(n_388),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_474),
.A2(n_249),
.B1(n_320),
.B2(n_227),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_446),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_474),
.B(n_398),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_446),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_469),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_474),
.B(n_285),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_437),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_437),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_461),
.B(n_183),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_502),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_502),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_502),
.A2(n_240),
.B1(n_257),
.B2(n_332),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_502),
.Y(n_646)
);

AND2x6_ASAP7_75t_L g647 ( 
.A(n_437),
.B(n_193),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_449),
.B(n_200),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_598),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_578),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_598),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_559),
.B(n_552),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_514),
.B(n_200),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_516),
.B(n_203),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_517),
.B(n_510),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_578),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_559),
.B(n_175),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_607),
.Y(n_658)
);

BUFx5_ASAP7_75t_L g659 ( 
.A(n_504),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_636),
.B(n_218),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_518),
.B(n_218),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_585),
.A2(n_314),
.B1(n_317),
.B2(n_286),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_644),
.B(n_578),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_532),
.B(n_220),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_538),
.B(n_212),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_532),
.B(n_223),
.Y(n_666)
);

AND2x4_ASAP7_75t_SL g667 ( 
.A(n_513),
.B(n_472),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_571),
.A2(n_256),
.B1(n_312),
.B2(n_273),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_532),
.B(n_512),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_611),
.B(n_390),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_609),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_609),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_540),
.B(n_214),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_523),
.B(n_223),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_547),
.B(n_216),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_528),
.B(n_421),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_524),
.B(n_243),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_525),
.B(n_243),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_527),
.B(n_229),
.C(n_224),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_526),
.B(n_244),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_592),
.B(n_230),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_529),
.Y(n_682)
);

OAI21xp33_ASAP7_75t_L g683 ( 
.A1(n_545),
.A2(n_257),
.B(n_240),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_621),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_507),
.B(n_287),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_637),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_SL g687 ( 
.A(n_563),
.B(n_500),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_615),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_536),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_528),
.B(n_421),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_554),
.A2(n_258),
.B(n_259),
.C(n_280),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_585),
.A2(n_258),
.B1(n_259),
.B2(n_280),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_568),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_531),
.B(n_244),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_545),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_541),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_592),
.B(n_233),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_543),
.B(n_251),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_544),
.B(n_251),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_549),
.B(n_255),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_629),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_SL g702 ( 
.A(n_584),
.B(n_187),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_507),
.A2(n_506),
.B1(n_511),
.B2(n_534),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_553),
.B(n_255),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_572),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_629),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_568),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_L g708 ( 
.A(n_566),
.B(n_250),
.C(n_248),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_632),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_573),
.B(n_575),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_579),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_632),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_597),
.B(n_235),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_582),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_589),
.B(n_256),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_591),
.B(n_260),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_597),
.B(n_237),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_585),
.A2(n_286),
.B1(n_314),
.B2(n_317),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_L g719 ( 
.A(n_561),
.B(n_292),
.C(n_293),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_600),
.B(n_245),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_604),
.B(n_264),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_633),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_506),
.A2(n_511),
.B1(n_535),
.B2(n_600),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_633),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_602),
.B(n_261),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_640),
.Y(n_726)
);

AO221x1_ASAP7_75t_L g727 ( 
.A1(n_630),
.A2(n_322),
.B1(n_331),
.B2(n_332),
.C(n_265),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_602),
.B(n_505),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_625),
.B(n_637),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_599),
.B(n_291),
.C(n_297),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_639),
.B(n_558),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_640),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_630),
.B(n_296),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_504),
.B(n_304),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_505),
.B(n_305),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_505),
.B(n_269),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_546),
.B(n_423),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_558),
.B(n_265),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_641),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_568),
.B(n_277),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_568),
.A2(n_306),
.B1(n_333),
.B2(n_316),
.Y(n_741)
);

NAND2x1p5_ASAP7_75t_L g742 ( 
.A(n_536),
.B(n_273),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_588),
.A2(n_315),
.B1(n_333),
.B2(n_316),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_643),
.B(n_290),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_646),
.B(n_306),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_630),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_641),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_631),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_590),
.B(n_279),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_546),
.A2(n_315),
.B(n_312),
.C(n_313),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_614),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

NAND2x1p5_ASAP7_75t_L g753 ( 
.A(n_519),
.B(n_313),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_624),
.B(n_450),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_610),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_627),
.B(n_450),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_631),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_635),
.B(n_451),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_504),
.A2(n_590),
.B1(n_522),
.B2(n_554),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_519),
.B(n_307),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_546),
.B(n_423),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_580),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_515),
.A2(n_322),
.B1(n_331),
.B2(n_252),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_605),
.A2(n_310),
.B1(n_330),
.B2(n_289),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_638),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_564),
.B(n_451),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_622),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_593),
.Y(n_768)
);

AND2x6_ASAP7_75t_SL g769 ( 
.A(n_612),
.B(n_215),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_564),
.B(n_451),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_606),
.A2(n_323),
.B1(n_321),
.B2(n_298),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_515),
.B(n_458),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_588),
.B(n_300),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_574),
.B(n_458),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_574),
.B(n_628),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_603),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_519),
.B(n_557),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_574),
.B(n_470),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_626),
.B(n_449),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_617),
.B(n_301),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_618),
.B(n_241),
.Y(n_781)
);

OAI221xp5_ASAP7_75t_L g782 ( 
.A1(n_645),
.A2(n_324),
.B1(n_308),
.B2(n_318),
.C(n_319),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_626),
.A2(n_328),
.B1(n_327),
.B2(n_222),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_634),
.A2(n_488),
.B1(n_470),
.B2(n_388),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_593),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_623),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_620),
.A2(n_488),
.B(n_470),
.C(n_426),
.Y(n_787)
);

AND2x6_ASAP7_75t_SL g788 ( 
.A(n_565),
.B(n_329),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_508),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_638),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_521),
.B(n_488),
.Y(n_791)
);

AND3x1_ASAP7_75t_L g792 ( 
.A(n_581),
.B(n_329),
.C(n_275),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_513),
.B(n_329),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_533),
.B(n_426),
.Y(n_794)
);

O2A1O1Ixp5_ASAP7_75t_L g795 ( 
.A1(n_548),
.A2(n_596),
.B(n_616),
.C(n_556),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_661),
.A2(n_648),
.B(n_560),
.C(n_567),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_653),
.A2(n_586),
.B(n_648),
.C(n_570),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_751),
.B(n_513),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_652),
.B(n_563),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_695),
.B(n_595),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_723),
.A2(n_482),
.B1(n_477),
.B2(n_509),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_767),
.B(n_626),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_762),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_765),
.Y(n_804)
);

OAI321xp33_ASAP7_75t_L g805 ( 
.A1(n_763),
.A2(n_329),
.A3(n_275),
.B1(n_241),
.B2(n_601),
.C(n_173),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_767),
.B(n_626),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_795),
.A2(n_616),
.B(n_520),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_684),
.B(n_520),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_755),
.B(n_626),
.Y(n_809)
);

OAI321xp33_ASAP7_75t_L g810 ( 
.A1(n_763),
.A2(n_275),
.A3(n_173),
.B1(n_539),
.B2(n_550),
.C(n_560),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_654),
.B(n_626),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_652),
.B(n_533),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_775),
.A2(n_569),
.B(n_619),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_701),
.B(n_555),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_701),
.B(n_555),
.Y(n_815)
);

AOI22x1_ASAP7_75t_L g816 ( 
.A1(n_706),
.A2(n_567),
.B1(n_570),
.B2(n_576),
.Y(n_816)
);

AOI21x1_ASAP7_75t_L g817 ( 
.A1(n_766),
.A2(n_562),
.B(n_576),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_706),
.B(n_555),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_781),
.B(n_642),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_709),
.B(n_556),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_728),
.B(n_556),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_703),
.A2(n_587),
.B1(n_594),
.B2(n_530),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_658),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_712),
.B(n_594),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_689),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_746),
.A2(n_583),
.B(n_613),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_768),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_770),
.A2(n_587),
.B(n_613),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_728),
.B(n_583),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_669),
.A2(n_551),
.B(n_530),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_712),
.B(n_551),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_729),
.A2(n_557),
.B(n_608),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_649),
.A2(n_647),
.B(n_173),
.C(n_275),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_785),
.B(n_608),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_734),
.A2(n_777),
.B(n_710),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_658),
.Y(n_836)
);

AND2x4_ASAP7_75t_SL g837 ( 
.A(n_650),
.B(n_173),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_759),
.A2(n_608),
.B1(n_577),
.B2(n_557),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_777),
.A2(n_557),
.B(n_577),
.Y(n_839)
);

AO22x1_ASAP7_75t_L g840 ( 
.A1(n_681),
.A2(n_647),
.B1(n_449),
.B2(n_14),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_681),
.A2(n_8),
.B(n_10),
.C(n_14),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_791),
.A2(n_542),
.B(n_647),
.Y(n_842)
);

O2A1O1Ixp5_ASAP7_75t_SL g843 ( 
.A1(n_660),
.A2(n_647),
.B(n_15),
.C(n_18),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_774),
.A2(n_542),
.B(n_647),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_657),
.B(n_542),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_776),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_778),
.A2(n_686),
.B(n_772),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_776),
.B(n_537),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_659),
.B(n_107),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_780),
.B(n_10),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_657),
.B(n_537),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_651),
.A2(n_18),
.B(n_19),
.C(n_22),
.Y(n_852)
);

NAND3xp33_ASAP7_75t_L g853 ( 
.A(n_697),
.B(n_23),
.C(n_25),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_671),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_697),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_722),
.B(n_26),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_650),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_724),
.B(n_28),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_794),
.A2(n_134),
.B(n_131),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_790),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_672),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_667),
.Y(n_862)
);

BUFx8_ASAP7_75t_L g863 ( 
.A(n_793),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_665),
.B(n_29),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_665),
.B(n_673),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_756),
.A2(n_31),
.B(n_32),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_693),
.Y(n_867)
);

OAI21xp33_ASAP7_75t_L g868 ( 
.A1(n_713),
.A2(n_31),
.B(n_32),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_673),
.B(n_33),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_738),
.A2(n_33),
.B(n_36),
.C(n_37),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_773),
.B(n_36),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_656),
.A2(n_62),
.B1(n_41),
.B2(n_42),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_748),
.A2(n_40),
.B(n_42),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_675),
.B(n_45),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_713),
.A2(n_46),
.B(n_47),
.C(n_50),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_773),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_689),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_659),
.B(n_47),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_758),
.A2(n_51),
.B(n_53),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_688),
.Y(n_880)
);

OAI321xp33_ASAP7_75t_L g881 ( 
.A1(n_717),
.A2(n_720),
.A3(n_725),
.B1(n_743),
.B2(n_668),
.C(n_741),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_676),
.B(n_54),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_675),
.B(n_54),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_667),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_717),
.A2(n_60),
.B(n_62),
.C(n_720),
.Y(n_885)
);

AOI21xp33_ASAP7_75t_L g886 ( 
.A1(n_725),
.A2(n_749),
.B(n_736),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_702),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_687),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_707),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_752),
.B(n_757),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_749),
.A2(n_733),
.B1(n_682),
.B2(n_696),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_752),
.A2(n_757),
.B(n_733),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_662),
.A2(n_718),
.B1(n_692),
.B2(n_711),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_662),
.A2(n_692),
.B(n_718),
.C(n_683),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_664),
.A2(n_666),
.B(n_789),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_726),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_769),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_736),
.B(n_783),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_726),
.A2(n_732),
.B(n_739),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_676),
.A2(n_690),
.B(n_691),
.C(n_740),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_690),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_705),
.B(n_714),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_739),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_760),
.A2(n_685),
.B(n_779),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_747),
.A2(n_745),
.B(n_744),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_737),
.B(n_761),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_737),
.B(n_761),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_787),
.A2(n_716),
.B(n_721),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_674),
.B(n_715),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_677),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_788),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_678),
.B(n_698),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_742),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_680),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_740),
.A2(n_679),
.B(n_708),
.C(n_782),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_694),
.A2(n_699),
.B(n_700),
.Y(n_916)
);

BUFx4f_ASAP7_75t_L g917 ( 
.A(n_786),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_704),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_735),
.A2(n_750),
.B1(n_792),
.B2(n_753),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_730),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_764),
.B(n_771),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_784),
.B(n_727),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_719),
.B(n_655),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_655),
.B(n_767),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_658),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_754),
.A2(n_731),
.B(n_663),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_655),
.B(n_767),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_762),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_655),
.A2(n_723),
.B1(n_703),
.B2(n_653),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_754),
.A2(n_731),
.B(n_663),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_L g932 ( 
.A1(n_780),
.A2(n_697),
.B(n_681),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_658),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_655),
.A2(n_723),
.B1(n_703),
.B2(n_653),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_785),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_655),
.A2(n_723),
.B1(n_703),
.B2(n_653),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_655),
.B(n_767),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_751),
.B(n_655),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_662),
.A2(n_718),
.B1(n_692),
.B2(n_706),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_658),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_L g941 ( 
.A(n_684),
.B(n_670),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_754),
.A2(n_731),
.B(n_663),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_655),
.B(n_767),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_762),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_689),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_892),
.A2(n_847),
.B(n_813),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_896),
.Y(n_947)
);

INVx4_ASAP7_75t_L g948 ( 
.A(n_825),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_925),
.B(n_928),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_896),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_937),
.A2(n_943),
.B(n_934),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_930),
.A2(n_936),
.B(n_931),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_861),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_927),
.A2(n_942),
.B(n_932),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_899),
.A2(n_807),
.B(n_895),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_845),
.B(n_809),
.Y(n_956)
);

OAI22x1_ASAP7_75t_L g957 ( 
.A1(n_898),
.A2(n_871),
.B1(n_938),
.B2(n_799),
.Y(n_957)
);

AND2x6_ASAP7_75t_SL g958 ( 
.A(n_848),
.B(n_798),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_825),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_938),
.B(n_865),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_835),
.A2(n_916),
.B(n_904),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_918),
.B(n_910),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_797),
.A2(n_886),
.B(n_908),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_825),
.B(n_945),
.Y(n_964)
);

OAI22x1_ASAP7_75t_L g965 ( 
.A1(n_898),
.A2(n_871),
.B1(n_799),
.B2(n_876),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_918),
.B(n_914),
.Y(n_966)
);

AOI21xp33_ASAP7_75t_L g967 ( 
.A1(n_881),
.A2(n_883),
.B(n_874),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_924),
.A2(n_921),
.B(n_894),
.C(n_891),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_939),
.B(n_909),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_830),
.A2(n_890),
.B(n_822),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_804),
.B(n_819),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_811),
.A2(n_802),
.B(n_806),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_890),
.A2(n_905),
.B(n_826),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_939),
.B(n_912),
.Y(n_974)
);

NAND3xp33_ASAP7_75t_L g975 ( 
.A(n_798),
.B(n_885),
.C(n_915),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_894),
.A2(n_915),
.B(n_900),
.C(n_893),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_821),
.B(n_829),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_884),
.Y(n_978)
);

OAI21xp33_ASAP7_75t_L g979 ( 
.A1(n_868),
.A2(n_902),
.B(n_929),
.Y(n_979)
);

INVx5_ASAP7_75t_L g980 ( 
.A(n_825),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_821),
.B(n_829),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_857),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_812),
.B(n_823),
.Y(n_983)
);

AO31x2_ASAP7_75t_L g984 ( 
.A1(n_797),
.A2(n_885),
.A3(n_900),
.B(n_838),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_823),
.B(n_836),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_824),
.A2(n_844),
.B(n_842),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_814),
.A2(n_820),
.B(n_818),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_810),
.A2(n_856),
.B(n_858),
.C(n_805),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_922),
.A2(n_907),
.B(n_853),
.C(n_913),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_843),
.A2(n_815),
.B(n_796),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_800),
.B(n_801),
.C(n_888),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_878),
.A2(n_831),
.B(n_849),
.Y(n_992)
);

AO31x2_ASAP7_75t_L g993 ( 
.A1(n_919),
.A2(n_855),
.A3(n_841),
.B(n_875),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_832),
.A2(n_854),
.B(n_880),
.Y(n_994)
);

AO31x2_ASAP7_75t_L g995 ( 
.A1(n_841),
.A2(n_875),
.A3(n_855),
.B(n_873),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_906),
.B(n_851),
.Y(n_996)
);

OA21x2_ASAP7_75t_L g997 ( 
.A1(n_878),
.A2(n_940),
.B(n_926),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_923),
.A2(n_839),
.B(n_857),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_901),
.B(n_944),
.Y(n_999)
);

BUFx5_ASAP7_75t_L g1000 ( 
.A(n_903),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_917),
.A2(n_901),
.B1(n_913),
.B2(n_887),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_933),
.B(n_834),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_935),
.B(n_882),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_834),
.A2(n_808),
.B(n_840),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_945),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_859),
.A2(n_866),
.B(n_879),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_945),
.B(n_877),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_833),
.A2(n_870),
.B(n_852),
.Y(n_1008)
);

AO31x2_ASAP7_75t_L g1009 ( 
.A1(n_872),
.A2(n_867),
.A3(n_837),
.B(n_860),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_945),
.B(n_941),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_846),
.B(n_803),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_827),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_889),
.B(n_884),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_837),
.B(n_920),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_889),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_917),
.Y(n_1016)
);

INVx3_ASAP7_75t_SL g1017 ( 
.A(n_848),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_862),
.A2(n_863),
.B(n_848),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_897),
.A2(n_863),
.B(n_911),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_930),
.A2(n_936),
.B(n_934),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_925),
.B(n_928),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_848),
.B(n_884),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_SL g1023 ( 
.A1(n_930),
.A2(n_936),
.B(n_934),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_925),
.B(n_928),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_817),
.A2(n_816),
.B(n_828),
.Y(n_1025)
);

OR2x6_ASAP7_75t_L g1026 ( 
.A(n_848),
.B(n_884),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_925),
.B(n_928),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_817),
.A2(n_816),
.B(n_828),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_861),
.Y(n_1029)
);

BUFx4_ASAP7_75t_SL g1030 ( 
.A(n_848),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_SL g1031 ( 
.A1(n_930),
.A2(n_936),
.B(n_934),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1032)
);

AOI221x1_ASAP7_75t_L g1033 ( 
.A1(n_932),
.A2(n_886),
.B1(n_871),
.B2(n_865),
.C(n_898),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_932),
.A2(n_865),
.B(n_886),
.C(n_898),
.Y(n_1034)
);

NOR2x1_ASAP7_75t_L g1035 ( 
.A(n_925),
.B(n_928),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_817),
.A2(n_816),
.B(n_828),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_SL g1038 ( 
.A(n_932),
.B(n_886),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_860),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_930),
.A2(n_936),
.B(n_934),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_861),
.Y(n_1041)
);

AND3x4_ASAP7_75t_L g1042 ( 
.A(n_941),
.B(n_730),
.C(n_776),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_925),
.B(n_928),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_886),
.B(n_932),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_938),
.B(n_819),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_L g1046 ( 
.A(n_932),
.B(n_865),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_SL g1047 ( 
.A1(n_930),
.A2(n_936),
.B(n_934),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_925),
.B(n_928),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_804),
.B(n_621),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_896),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_896),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_817),
.A2(n_816),
.B(n_828),
.Y(n_1054)
);

NAND2x1p5_ASAP7_75t_L g1055 ( 
.A(n_825),
.B(n_650),
.Y(n_1055)
);

AOI21xp33_ASAP7_75t_L g1056 ( 
.A1(n_932),
.A2(n_865),
.B(n_898),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_938),
.B(n_865),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_850),
.A2(n_869),
.B(n_864),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1059)
);

INVx3_ASAP7_75t_SL g1060 ( 
.A(n_848),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_938),
.B(n_819),
.Y(n_1061)
);

NOR2x1_ASAP7_75t_L g1062 ( 
.A(n_925),
.B(n_928),
.Y(n_1062)
);

AOI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_932),
.A2(n_865),
.B(n_898),
.Y(n_1063)
);

INVxp67_ASAP7_75t_SL g1064 ( 
.A(n_925),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_925),
.B(n_928),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_804),
.B(n_621),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_930),
.A2(n_936),
.A3(n_934),
.B(n_797),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_925),
.B(n_928),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_SL g1071 ( 
.A1(n_850),
.A2(n_869),
.B(n_864),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_930),
.A2(n_936),
.B(n_934),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_SL g1074 ( 
.A1(n_925),
.A2(n_937),
.B(n_928),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_865),
.A2(n_886),
.B(n_661),
.C(n_654),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_925),
.B(n_928),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_846),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_930),
.A2(n_936),
.B(n_934),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1057),
.A2(n_960),
.B1(n_1034),
.B2(n_1064),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_978),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_1039),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_1051),
.B(n_1067),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_1077),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_960),
.A2(n_1048),
.B1(n_1076),
.B2(n_1027),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_980),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_953),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_949),
.B(n_1021),
.Y(n_1087)
);

OAI33xp33_ASAP7_75t_L g1088 ( 
.A1(n_962),
.A2(n_966),
.A3(n_1076),
.B1(n_1024),
.B2(n_1021),
.B3(n_949),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_999),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1024),
.B(n_1027),
.Y(n_1090)
);

INVx3_ASAP7_75t_SL g1091 ( 
.A(n_1017),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1043),
.B(n_1048),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_950),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_1020),
.A2(n_1073),
.B(n_1040),
.C(n_1078),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1023),
.A2(n_1047),
.B(n_1031),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_980),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1045),
.B(n_1061),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1043),
.B(n_1065),
.Y(n_1098)
);

AOI222xp33_ASAP7_75t_L g1099 ( 
.A1(n_957),
.A2(n_965),
.B1(n_1078),
.B2(n_1020),
.C1(n_1040),
.C2(n_1073),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_1011),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_952),
.A2(n_961),
.B(n_954),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_952),
.A2(n_954),
.B(n_951),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1038),
.A2(n_996),
.B1(n_991),
.B2(n_1042),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1069),
.A2(n_981),
.B1(n_977),
.B2(n_975),
.Y(n_1104)
);

OR2x6_ASAP7_75t_L g1105 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1105)
);

AOI221x1_ASAP7_75t_L g1106 ( 
.A1(n_967),
.A2(n_1056),
.B1(n_1063),
.B2(n_963),
.C(n_976),
.Y(n_1106)
);

OA21x2_ASAP7_75t_L g1107 ( 
.A1(n_963),
.A2(n_990),
.B(n_955),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1003),
.B(n_1014),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_1013),
.B(n_1016),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_971),
.B(n_1056),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_962),
.B(n_966),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_1022),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_SL g1113 ( 
.A1(n_968),
.A2(n_974),
.B(n_969),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_959),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1035),
.B(n_1062),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1063),
.B(n_1012),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_1038),
.B(n_969),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_951),
.A2(n_1037),
.B(n_1050),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1030),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1007),
.B(n_1016),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1032),
.B(n_1049),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1044),
.B(n_977),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_980),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_958),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1046),
.A2(n_1001),
.B1(n_979),
.B2(n_1010),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_1007),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1059),
.A2(n_1066),
.B(n_1070),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1010),
.B(n_1001),
.Y(n_1129)
);

INVx5_ASAP7_75t_L g1130 ( 
.A(n_959),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1013),
.B(n_1026),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_967),
.A2(n_974),
.B1(n_956),
.B2(n_981),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1072),
.B(n_1033),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1074),
.B(n_989),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1008),
.A2(n_1029),
.B1(n_1041),
.B2(n_956),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1005),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_972),
.A2(n_1075),
.B(n_946),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1015),
.B(n_1009),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1018),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1009),
.B(n_964),
.Y(n_1140)
);

OAI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_988),
.A2(n_1002),
.B(n_992),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_983),
.B(n_1002),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_964),
.B(n_948),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_983),
.B(n_1068),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_948),
.B(n_1005),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_980),
.B(n_1005),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1060),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1068),
.B(n_993),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1068),
.B(n_993),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1055),
.Y(n_1151)
);

AOI21xp33_ASAP7_75t_L g1152 ( 
.A1(n_985),
.A2(n_1053),
.B(n_1052),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_982),
.Y(n_1153)
);

AND2x6_ASAP7_75t_L g1154 ( 
.A(n_993),
.B(n_984),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_995),
.B(n_984),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_956),
.A2(n_997),
.B1(n_1000),
.B2(n_998),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_995),
.B(n_984),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_995),
.B(n_956),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1000),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1019),
.B(n_1006),
.Y(n_1160)
);

AND2x6_ASAP7_75t_L g1161 ( 
.A(n_1000),
.B(n_1071),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_1000),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_987),
.B(n_970),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_R g1164 ( 
.A(n_1058),
.B(n_986),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_994),
.B(n_973),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1025),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1028),
.B(n_1036),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1054),
.B(n_1013),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_SL g1169 ( 
.A1(n_968),
.A2(n_1034),
.B(n_976),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1011),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_959),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1057),
.B(n_960),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_980),
.Y(n_1173)
);

OA21x2_ASAP7_75t_L g1174 ( 
.A1(n_963),
.A2(n_990),
.B(n_952),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1077),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_SL g1176 ( 
.A(n_980),
.B(n_962),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1057),
.A2(n_932),
.B1(n_898),
.B2(n_871),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1023),
.A2(n_1047),
.B(n_1031),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1057),
.B(n_932),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1013),
.B(n_1016),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1057),
.B(n_960),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1057),
.B(n_960),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1077),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1077),
.Y(n_1184)
);

OAI21xp33_ASAP7_75t_L g1185 ( 
.A1(n_1057),
.A2(n_932),
.B(n_938),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1011),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1057),
.B(n_960),
.Y(n_1187)
);

INVx3_ASAP7_75t_SL g1188 ( 
.A(n_1039),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_SL g1189 ( 
.A1(n_1020),
.A2(n_871),
.B(n_886),
.C(n_1040),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1051),
.B(n_1067),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1057),
.B(n_960),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1034),
.A2(n_932),
.B(n_886),
.C(n_865),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1051),
.B(n_1067),
.Y(n_1193)
);

OR2x6_ASAP7_75t_L g1194 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1057),
.B(n_932),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1077),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1011),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_978),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1051),
.B(n_1067),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1045),
.B(n_1061),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1057),
.B(n_932),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1045),
.A2(n_932),
.B1(n_898),
.B2(n_865),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1045),
.B(n_1061),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1077),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_953),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1077),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_947),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1057),
.B(n_960),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_991),
.B(n_803),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_980),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1023),
.A2(n_1047),
.B(n_1031),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_953),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1086),
.Y(n_1213)
);

OA21x2_ASAP7_75t_L g1214 ( 
.A1(n_1137),
.A2(n_1119),
.B(n_1128),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1179),
.A2(n_1201),
.B1(n_1195),
.B2(n_1177),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1179),
.A2(n_1201),
.B1(n_1195),
.B2(n_1103),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1079),
.A2(n_1191),
.B1(n_1172),
.B2(n_1181),
.Y(n_1217)
);

BUFx5_ASAP7_75t_L g1218 ( 
.A(n_1161),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1081),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1177),
.A2(n_1185),
.B1(n_1099),
.B2(n_1202),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1082),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1123),
.A2(n_1110),
.B1(n_1118),
.B2(n_1104),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1123),
.A2(n_1118),
.B1(n_1208),
.B2(n_1182),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1093),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_1081),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1089),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_1188),
.Y(n_1227)
);

BUFx8_ASAP7_75t_L g1228 ( 
.A(n_1183),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1097),
.A2(n_1200),
.B1(n_1203),
.B2(n_1209),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1083),
.Y(n_1230)
);

AOI22x1_ASAP7_75t_SL g1231 ( 
.A1(n_1125),
.A2(n_1162),
.B1(n_1206),
.B2(n_1100),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1205),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1212),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1187),
.A2(n_1092),
.B1(n_1098),
.B2(n_1090),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1154),
.A2(n_1211),
.B1(n_1095),
.B2(n_1178),
.Y(n_1235)
);

INVx11_ASAP7_75t_L g1236 ( 
.A(n_1112),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1108),
.B(n_1089),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1141),
.A2(n_1084),
.B1(n_1174),
.B2(n_1087),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1117),
.B(n_1127),
.Y(n_1239)
);

CKINVDCx11_ASAP7_75t_R g1240 ( 
.A(n_1188),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1121),
.B(n_1170),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1175),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1174),
.A2(n_1088),
.B1(n_1102),
.B2(n_1129),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_1096),
.B(n_1124),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1192),
.A2(n_1106),
.B(n_1126),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1207),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1105),
.B(n_1114),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1164),
.A2(n_1189),
.B(n_1102),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1130),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1154),
.A2(n_1162),
.B1(n_1174),
.B2(n_1169),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1153),
.Y(n_1251)
);

INVx5_ASAP7_75t_L g1252 ( 
.A(n_1173),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1186),
.B(n_1197),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1111),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1116),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1155),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1173),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1138),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1190),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1080),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1080),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1088),
.A2(n_1154),
.B1(n_1193),
.B2(n_1199),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1154),
.A2(n_1132),
.B1(n_1101),
.B2(n_1134),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1196),
.B(n_1204),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1173),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1154),
.A2(n_1101),
.B1(n_1114),
.B2(n_1105),
.Y(n_1266)
);

CKINVDCx11_ASAP7_75t_R g1267 ( 
.A(n_1091),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1083),
.A2(n_1105),
.B1(n_1194),
.B2(n_1114),
.Y(n_1268)
);

CKINVDCx14_ASAP7_75t_R g1269 ( 
.A(n_1131),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1115),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1157),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1194),
.A2(n_1189),
.B1(n_1094),
.B2(n_1148),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_SL g1273 ( 
.A1(n_1192),
.A2(n_1135),
.B(n_1160),
.Y(n_1273)
);

INVxp67_ASAP7_75t_L g1274 ( 
.A(n_1184),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_SL g1275 ( 
.A1(n_1194),
.A2(n_1094),
.B1(n_1148),
.B2(n_1122),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1107),
.A2(n_1139),
.B1(n_1142),
.B2(n_1133),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1136),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1107),
.A2(n_1144),
.B1(n_1150),
.B2(n_1149),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1109),
.B(n_1180),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1198),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1180),
.B(n_1146),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1113),
.B(n_1198),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1158),
.A2(n_1176),
.B1(n_1107),
.B2(n_1161),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1091),
.A2(n_1140),
.B1(n_1168),
.B2(n_1161),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1168),
.A2(n_1161),
.B1(n_1145),
.B2(n_1143),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1210),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1171),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1159),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1130),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1163),
.A2(n_1166),
.B(n_1167),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1210),
.Y(n_1291)
);

INVx3_ASAP7_75t_SL g1292 ( 
.A(n_1147),
.Y(n_1292)
);

NAND2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1096),
.B(n_1124),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1161),
.A2(n_1210),
.B1(n_1130),
.B2(n_1151),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1147),
.Y(n_1295)
);

CKINVDCx11_ASAP7_75t_R g1296 ( 
.A(n_1151),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1135),
.A2(n_1156),
.B1(n_1152),
.B2(n_1167),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1165),
.A2(n_932),
.B1(n_1195),
.B2(n_1179),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1120),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1086),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1086),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1177),
.A2(n_1057),
.B1(n_865),
.B2(n_1179),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1179),
.B(n_932),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1081),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1177),
.A2(n_561),
.B1(n_642),
.B2(n_792),
.Y(n_1305)
);

INVx4_ASAP7_75t_L g1306 ( 
.A(n_1085),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1131),
.B(n_1109),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1202),
.A2(n_865),
.B1(n_960),
.B2(n_1057),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1081),
.Y(n_1309)
);

AO21x1_ASAP7_75t_L g1310 ( 
.A1(n_1192),
.A2(n_886),
.B(n_865),
.Y(n_1310)
);

BUFx4f_ASAP7_75t_SL g1311 ( 
.A(n_1081),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1179),
.A2(n_898),
.B1(n_932),
.B2(n_865),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1202),
.A2(n_865),
.B1(n_960),
.B2(n_1057),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1089),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1271),
.B(n_1278),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_SL g1316 ( 
.A1(n_1266),
.A2(n_1310),
.B(n_1282),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1226),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1256),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1258),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1213),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1290),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1290),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1222),
.B(n_1250),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1226),
.B(n_1314),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1314),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1247),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1222),
.B(n_1248),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1232),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1223),
.B(n_1254),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1247),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1285),
.B(n_1266),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1260),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1233),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1300),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1301),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1234),
.A2(n_1302),
.B(n_1312),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1223),
.B(n_1303),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1251),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1245),
.B(n_1243),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1273),
.B(n_1297),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1250),
.B(n_1298),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1242),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1218),
.Y(n_1343)
);

NOR2xp67_ASAP7_75t_SL g1344 ( 
.A(n_1252),
.B(n_1249),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1288),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1214),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1261),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1298),
.B(n_1239),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1243),
.B(n_1263),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1263),
.A2(n_1276),
.B(n_1238),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1218),
.Y(n_1351)
);

CKINVDCx6p67_ASAP7_75t_R g1352 ( 
.A(n_1240),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1276),
.A2(n_1238),
.B(n_1220),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1296),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1218),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1218),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1284),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1259),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1305),
.A2(n_1303),
.B1(n_1216),
.B2(n_1215),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1283),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_SL g1361 ( 
.A1(n_1308),
.A2(n_1313),
.B(n_1289),
.C(n_1255),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1224),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1221),
.B(n_1215),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1246),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1275),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1262),
.B(n_1220),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1275),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1237),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1235),
.A2(n_1217),
.B(n_1229),
.C(n_1272),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1217),
.A2(n_1313),
.B(n_1308),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1235),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1230),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1272),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1268),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1280),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1294),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1294),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1241),
.B(n_1262),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1264),
.B(n_1274),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1274),
.B(n_1281),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1270),
.A2(n_1277),
.B(n_1253),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1228),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1292),
.B(n_1307),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1228),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1370),
.A2(n_1267),
.B1(n_1269),
.B2(n_1311),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1360),
.B(n_1279),
.Y(n_1386)
);

INVx3_ASAP7_75t_SL g1387 ( 
.A(n_1352),
.Y(n_1387)
);

AOI221xp5_ASAP7_75t_L g1388 ( 
.A1(n_1336),
.A2(n_1269),
.B1(n_1309),
.B2(n_1304),
.C(n_1227),
.Y(n_1388)
);

INVxp67_ASAP7_75t_SL g1389 ( 
.A(n_1321),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1371),
.B(n_1265),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1330),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_L g1392 ( 
.A(n_1359),
.B(n_1231),
.C(n_1286),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1350),
.B(n_1257),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1315),
.B(n_1292),
.Y(n_1394)
);

AOI211xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1336),
.A2(n_1311),
.B(n_1225),
.C(n_1219),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1318),
.B(n_1329),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1350),
.B(n_1287),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1321),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1337),
.B(n_1306),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1346),
.Y(n_1400)
);

INVxp67_ASAP7_75t_L g1401 ( 
.A(n_1381),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1327),
.B(n_1291),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1369),
.A2(n_1244),
.B(n_1293),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1327),
.B(n_1295),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1322),
.B(n_1236),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1343),
.B(n_1351),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1359),
.A2(n_1299),
.B1(n_1340),
.B2(n_1341),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1340),
.B(n_1351),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1340),
.B(n_1355),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1317),
.B(n_1325),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1381),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1324),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1340),
.A2(n_1361),
.B(n_1366),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1340),
.B(n_1356),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1396),
.B(n_1358),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1388),
.A2(n_1341),
.B1(n_1323),
.B2(n_1357),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1408),
.B(n_1331),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1410),
.B(n_1345),
.Y(n_1418)
);

AOI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1413),
.A2(n_1365),
.B1(n_1367),
.B2(n_1373),
.C(n_1323),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1392),
.A2(n_1366),
.B1(n_1367),
.B2(n_1365),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1395),
.A2(n_1357),
.B(n_1331),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_SL g1422 ( 
.A(n_1387),
.B(n_1352),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1395),
.B(n_1339),
.C(n_1378),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1392),
.A2(n_1373),
.B1(n_1363),
.B2(n_1339),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1388),
.A2(n_1384),
.B(n_1382),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1412),
.B(n_1342),
.Y(n_1426)
);

AND2x6_ASAP7_75t_L g1427 ( 
.A(n_1409),
.B(n_1326),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1412),
.B(n_1368),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1413),
.A2(n_1316),
.B1(n_1348),
.B2(n_1372),
.C(n_1377),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1407),
.A2(n_1374),
.B1(n_1349),
.B2(n_1354),
.Y(n_1430)
);

NAND3xp33_ASAP7_75t_L g1431 ( 
.A(n_1403),
.B(n_1348),
.C(n_1326),
.Y(n_1431)
);

OAI221xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1385),
.A2(n_1349),
.B1(n_1377),
.B2(n_1376),
.C(n_1374),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1404),
.B(n_1338),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1403),
.B(n_1326),
.Y(n_1434)
);

NAND3xp33_ASAP7_75t_L g1435 ( 
.A(n_1397),
.B(n_1326),
.C(n_1353),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1404),
.B(n_1399),
.Y(n_1436)
);

NAND4xp25_ASAP7_75t_L g1437 ( 
.A(n_1399),
.B(n_1379),
.C(n_1372),
.D(n_1380),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1402),
.B(n_1324),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1397),
.B(n_1326),
.C(n_1353),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1387),
.A2(n_1354),
.B1(n_1380),
.B2(n_1379),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1414),
.A2(n_1382),
.B(n_1384),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1394),
.B(n_1316),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1387),
.A2(n_1354),
.B1(n_1405),
.B2(n_1383),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1390),
.B(n_1320),
.Y(n_1444)
);

OAI21xp33_ASAP7_75t_L g1445 ( 
.A1(n_1386),
.A2(n_1333),
.B(n_1335),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1397),
.B(n_1362),
.C(n_1364),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1393),
.B(n_1319),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1400),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1402),
.B(n_1391),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1402),
.B(n_1319),
.Y(n_1450)
);

OAI21xp33_ASAP7_75t_L g1451 ( 
.A1(n_1386),
.A2(n_1334),
.B(n_1328),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1427),
.B(n_1406),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1450),
.B(n_1398),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1448),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1448),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1438),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1436),
.B(n_1437),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1447),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1442),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1438),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1444),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1427),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1449),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1427),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1435),
.B(n_1401),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1427),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1442),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1427),
.B(n_1406),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1439),
.B(n_1401),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1434),
.B(n_1344),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1426),
.B(n_1411),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1446),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1418),
.B(n_1411),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1456),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1465),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1454),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1464),
.B(n_1452),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1470),
.B(n_1422),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1472),
.B(n_1445),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1456),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1460),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1454),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1472),
.B(n_1445),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1460),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1459),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1459),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1455),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1462),
.B(n_1434),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1465),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1455),
.Y(n_1490)
);

OA21x2_ASAP7_75t_L g1491 ( 
.A1(n_1465),
.A2(n_1431),
.B(n_1389),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1473),
.B(n_1428),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1463),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1463),
.Y(n_1494)
);

NOR2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1462),
.B(n_1354),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1455),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1454),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1454),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1453),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1464),
.B(n_1449),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1462),
.B(n_1417),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1464),
.B(n_1452),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1453),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1467),
.B(n_1451),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1467),
.B(n_1451),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1457),
.B(n_1354),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1452),
.B(n_1468),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1458),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1473),
.B(n_1415),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1462),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1462),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1473),
.B(n_1433),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1476),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1474),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1474),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1477),
.B(n_1502),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1479),
.B(n_1457),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1479),
.B(n_1461),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1476),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1480),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1480),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1476),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1477),
.B(n_1466),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1481),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1481),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1482),
.Y(n_1526)
);

NAND2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_1466),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1482),
.Y(n_1528)
);

AOI21xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1478),
.A2(n_1506),
.B(n_1425),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1475),
.B(n_1499),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1484),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1485),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1502),
.B(n_1466),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1483),
.B(n_1485),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1495),
.B(n_1466),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1475),
.B(n_1471),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1491),
.B(n_1466),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1484),
.Y(n_1538)
);

AOI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1489),
.A2(n_1469),
.B(n_1440),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1487),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1487),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1490),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1486),
.B(n_1461),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1499),
.B(n_1471),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1504),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1490),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1486),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1503),
.B(n_1471),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1507),
.B(n_1501),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1496),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1482),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1496),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1504),
.B(n_1505),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1510),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1535),
.B(n_1495),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1534),
.B(n_1532),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1514),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1545),
.B(n_1505),
.Y(n_1558)
);

CKINVDCx16_ASAP7_75t_R g1559 ( 
.A(n_1547),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1516),
.B(n_1488),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1554),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1536),
.B(n_1509),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1517),
.A2(n_1529),
.B(n_1553),
.Y(n_1564)
);

NOR2x1_ASAP7_75t_L g1565 ( 
.A(n_1554),
.B(n_1510),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1554),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1516),
.B(n_1488),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1519),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1549),
.B(n_1488),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1530),
.B(n_1509),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1529),
.A2(n_1491),
.B(n_1421),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1549),
.B(n_1488),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1518),
.B(n_1503),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1514),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1515),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1515),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1535),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1492),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1535),
.B(n_1523),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1535),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_SL g1581 ( 
.A(n_1539),
.B(n_1443),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1520),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1544),
.B(n_1492),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1520),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1521),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1523),
.Y(n_1586)
);

NOR2x1_ASAP7_75t_L g1587 ( 
.A(n_1543),
.B(n_1491),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1533),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1533),
.Y(n_1589)
);

NAND3xp33_ASAP7_75t_L g1590 ( 
.A(n_1544),
.B(n_1491),
.C(n_1424),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1559),
.B(n_1512),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1557),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1564),
.B(n_1548),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1556),
.B(n_1512),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1574),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1556),
.B(n_1548),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1581),
.B(n_1501),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1558),
.B(n_1501),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1571),
.A2(n_1537),
.B(n_1527),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1555),
.B(n_1501),
.Y(n_1600)
);

OAI211xp5_ASAP7_75t_L g1601 ( 
.A1(n_1565),
.A2(n_1590),
.B(n_1587),
.C(n_1580),
.Y(n_1601)
);

OAI222xp33_ASAP7_75t_L g1602 ( 
.A1(n_1577),
.A2(n_1537),
.B1(n_1527),
.B2(n_1469),
.C1(n_1432),
.C2(n_1470),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1575),
.Y(n_1603)
);

INVxp67_ASAP7_75t_SL g1604 ( 
.A(n_1562),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1576),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1566),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1582),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1573),
.A2(n_1537),
.B(n_1527),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1584),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1579),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1578),
.B(n_1521),
.Y(n_1611)
);

AOI21xp33_ASAP7_75t_L g1612 ( 
.A1(n_1561),
.A2(n_1525),
.B(n_1524),
.Y(n_1612)
);

AOI211xp5_ASAP7_75t_L g1613 ( 
.A1(n_1561),
.A2(n_1420),
.B(n_1441),
.C(n_1429),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1570),
.A2(n_1416),
.B1(n_1511),
.B2(n_1470),
.C(n_1419),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1585),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1511),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1591),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1604),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1604),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1610),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1611),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1600),
.B(n_1555),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1591),
.B(n_1555),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1593),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_SL g1625 ( 
.A(n_1602),
.B(n_1586),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1592),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1596),
.B(n_1570),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1595),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1616),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1606),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1603),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1605),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1607),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1597),
.B(n_1579),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1609),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_1579),
.Y(n_1636)
);

AOI21xp33_ASAP7_75t_L g1637 ( 
.A1(n_1617),
.A2(n_1601),
.B(n_1599),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1624),
.B(n_1594),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1620),
.B(n_1613),
.Y(n_1639)
);

NOR2xp67_ASAP7_75t_L g1640 ( 
.A(n_1629),
.B(n_1598),
.Y(n_1640)
);

OAI222xp33_ASAP7_75t_L g1641 ( 
.A1(n_1618),
.A2(n_1614),
.B1(n_1608),
.B2(n_1589),
.C1(n_1588),
.C2(n_1578),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1620),
.B(n_1594),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1629),
.B(n_1615),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1627),
.B(n_1616),
.Y(n_1644)
);

AOI221x1_ASAP7_75t_L g1645 ( 
.A1(n_1619),
.A2(n_1612),
.B1(n_1568),
.B2(n_1531),
.C(n_1525),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1625),
.A2(n_1563),
.B1(n_1583),
.B2(n_1569),
.C(n_1572),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1619),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1623),
.B(n_1563),
.C(n_1583),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1640),
.B(n_1622),
.Y(n_1649)
);

AOI322xp5_ASAP7_75t_L g1650 ( 
.A1(n_1638),
.A2(n_1630),
.A3(n_1626),
.B1(n_1633),
.B2(n_1632),
.C1(n_1628),
.C2(n_1621),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1648),
.B(n_1621),
.Y(n_1651)
);

NAND4xp75_ASAP7_75t_L g1652 ( 
.A(n_1645),
.B(n_1634),
.C(n_1636),
.D(n_1622),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1637),
.B(n_1635),
.C(n_1631),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_L g1654 ( 
.A(n_1642),
.B(n_1634),
.C(n_1631),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_SL g1655 ( 
.A(n_1641),
.B(n_1636),
.Y(n_1655)
);

NOR2x1_ASAP7_75t_L g1656 ( 
.A(n_1647),
.B(n_1635),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1646),
.A2(n_1572),
.B(n_1569),
.Y(n_1657)
);

OAI211xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1639),
.A2(n_1644),
.B(n_1643),
.C(n_1568),
.Y(n_1658)
);

NOR3x1_ASAP7_75t_L g1659 ( 
.A(n_1639),
.B(n_1511),
.C(n_1524),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1653),
.A2(n_1567),
.B1(n_1560),
.B2(n_1519),
.C(n_1522),
.Y(n_1660)
);

AOI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1651),
.A2(n_1655),
.B(n_1649),
.C(n_1658),
.Y(n_1661)
);

AOI211xp5_ASAP7_75t_L g1662 ( 
.A1(n_1654),
.A2(n_1567),
.B(n_1560),
.C(n_1430),
.Y(n_1662)
);

NAND3xp33_ASAP7_75t_L g1663 ( 
.A(n_1650),
.B(n_1522),
.C(n_1519),
.Y(n_1663)
);

NOR4xp25_ASAP7_75t_SL g1664 ( 
.A(n_1652),
.B(n_1531),
.C(n_1538),
.D(n_1550),
.Y(n_1664)
);

AO22x1_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1656),
.B1(n_1659),
.B2(n_1657),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1663),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1661),
.A2(n_1538),
.B1(n_1546),
.B2(n_1552),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1660),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1662),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1660),
.A2(n_1522),
.B1(n_1528),
.B2(n_1423),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1665),
.B(n_1540),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_L g1672 ( 
.A(n_1666),
.B(n_1332),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1668),
.B(n_1540),
.Y(n_1673)
);

NOR3xp33_ASAP7_75t_L g1674 ( 
.A(n_1669),
.B(n_1375),
.C(n_1347),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1667),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1671),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1672),
.Y(n_1677)
);

XNOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1675),
.B(n_1347),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1670),
.B1(n_1673),
.B2(n_1674),
.Y(n_1679)
);

NAND4xp25_ASAP7_75t_SL g1680 ( 
.A(n_1679),
.B(n_1676),
.C(n_1677),
.D(n_1528),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1680),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1680),
.A2(n_1551),
.B1(n_1526),
.B2(n_1513),
.Y(n_1682)
);

A2O1A1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1681),
.A2(n_1528),
.B(n_1551),
.C(n_1526),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1682),
.A2(n_1513),
.B1(n_1550),
.B2(n_1552),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1684),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1683),
.A2(n_1542),
.B(n_1541),
.Y(n_1686)
);

OAI222xp33_ASAP7_75t_L g1687 ( 
.A1(n_1685),
.A2(n_1546),
.B1(n_1542),
.B2(n_1541),
.C1(n_1375),
.C2(n_1470),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1686),
.B1(n_1494),
.B2(n_1493),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1498),
.B1(n_1497),
.B2(n_1500),
.C(n_1508),
.Y(n_1689)
);

AOI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1689),
.A2(n_1344),
.B(n_1469),
.C(n_1498),
.Y(n_1690)
);


endmodule