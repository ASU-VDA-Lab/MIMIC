module real_aes_10149_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
HB1xp67_ASAP7_75t_L g655 ( .A(n_0), .Y(n_655) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_1), .Y(n_557) );
INVx1_ASAP7_75t_L g577 ( .A(n_1), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_2), .A2(n_73), .B1(n_589), .B2(n_600), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_2), .A2(n_73), .B1(n_628), .B2(n_632), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_3), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_4), .B(n_119), .Y(n_191) );
INVx2_ASAP7_75t_L g481 ( .A(n_5), .Y(n_481) );
BUFx2_ASAP7_75t_L g528 ( .A(n_6), .Y(n_528) );
INVx1_ASAP7_75t_L g573 ( .A(n_6), .Y(n_573) );
BUFx2_ASAP7_75t_L g593 ( .A(n_6), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_7), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_8), .B(n_125), .Y(n_188) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_8), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_9), .B(n_111), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_10), .B(n_111), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_11), .B(n_187), .Y(n_265) );
AND2x2_ASAP7_75t_L g161 ( .A(n_12), .B(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_13), .A2(n_24), .B1(n_477), .B2(n_487), .Y(n_476) );
INVx1_ASAP7_75t_L g566 ( .A(n_13), .Y(n_566) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_15), .A2(n_70), .B1(n_515), .B2(n_518), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_15), .A2(n_70), .B1(n_560), .B2(n_562), .C(n_565), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_16), .B(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_17), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_18), .B(n_170), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_19), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_19), .Y(n_472) );
NAND2xp33_ASAP7_75t_L g232 ( .A(n_20), .B(n_118), .Y(n_232) );
NAND2xp33_ASAP7_75t_L g126 ( .A(n_21), .B(n_118), .Y(n_126) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_22), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_23), .Y(n_137) );
INVx1_ASAP7_75t_L g619 ( .A(n_24), .Y(n_619) );
INVx1_ASAP7_75t_L g526 ( .A(n_25), .Y(n_526) );
INVx1_ASAP7_75t_L g684 ( .A(n_25), .Y(n_684) );
INVx1_ASAP7_75t_L g543 ( .A(n_26), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_27), .B(n_209), .Y(n_235) );
OAI21x1_ASAP7_75t_L g113 ( .A1(n_28), .A2(n_47), .B(n_114), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_29), .A2(n_143), .B(n_166), .C(n_167), .Y(n_165) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_29), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_30), .B(n_141), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_31), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g268 ( .A(n_32), .B(n_147), .Y(n_268) );
AND2x6_ASAP7_75t_L g83 ( .A(n_33), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_33), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_33), .B(n_643), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_34), .B(n_140), .Y(n_223) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_35), .A2(n_57), .B1(n_531), .B2(n_538), .C(n_542), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_35), .A2(n_57), .B1(n_589), .B2(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g513 ( .A(n_36), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_37), .B(n_124), .Y(n_123) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_38), .B(n_147), .Y(n_192) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_38), .Y(n_686) );
INVx1_ASAP7_75t_L g84 ( .A(n_39), .Y(n_84) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_39), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_40), .Y(n_151) );
INVx1_ASAP7_75t_L g510 ( .A(n_41), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_42), .B(n_147), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_43), .Y(n_201) );
AND2x2_ASAP7_75t_L g169 ( .A(n_44), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_45), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g537 ( .A(n_46), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_48), .Y(n_234) );
NAND2xp33_ASAP7_75t_L g219 ( .A(n_49), .B(n_90), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_50), .B(n_231), .Y(n_267) );
BUFx10_ASAP7_75t_L g678 ( .A(n_51), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_52), .B(n_89), .Y(n_120) );
INVx1_ASAP7_75t_L g597 ( .A(n_53), .Y(n_597) );
INVx1_ASAP7_75t_L g558 ( .A(n_54), .Y(n_558) );
INVx2_ASAP7_75t_L g576 ( .A(n_54), .Y(n_576) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_55), .A2(n_497), .B(n_502), .C(n_505), .Y(n_496) );
INVx1_ASAP7_75t_L g569 ( .A(n_55), .Y(n_569) );
NAND2xp33_ASAP7_75t_L g224 ( .A(n_56), .B(n_125), .Y(n_224) );
INVx1_ASAP7_75t_L g547 ( .A(n_58), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_59), .B(n_118), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_60), .Y(n_168) );
INVx2_ASAP7_75t_L g114 ( .A(n_61), .Y(n_114) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_62), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_63), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_64), .B(n_211), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_65), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_66), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g160 ( .A(n_67), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_68), .Y(n_139) );
AND2x2_ASAP7_75t_L g152 ( .A(n_69), .B(n_111), .Y(n_152) );
INVx2_ASAP7_75t_L g534 ( .A(n_71), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_72), .B(n_170), .Y(n_225) );
INVx1_ASAP7_75t_L g484 ( .A(n_74), .Y(n_484) );
BUFx3_ASAP7_75t_L g493 ( .A(n_74), .Y(n_493) );
INVx1_ASAP7_75t_L g486 ( .A(n_75), .Y(n_486) );
BUFx3_ASAP7_75t_L g495 ( .A(n_75), .Y(n_495) );
INVx1_ASAP7_75t_L g598 ( .A(n_76), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_95), .B(n_470), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx8_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_82), .A2(n_135), .B(n_144), .Y(n_134) );
NOR2xp67_ASAP7_75t_L g155 ( .A(n_82), .B(n_156), .Y(n_155) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
BUFx2_ASAP7_75t_L g269 ( .A(n_83), .Y(n_269) );
INVxp67_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g696 ( .A1(n_86), .A2(n_697), .B(n_698), .Y(n_696) );
NAND2xp33_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g202 ( .A(n_89), .Y(n_202) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g187 ( .A(n_90), .Y(n_187) );
INVx2_ASAP7_75t_L g221 ( .A(n_90), .Y(n_221) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g119 ( .A(n_91), .Y(n_119) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_91), .Y(n_125) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_91), .Y(n_150) );
INVx1_ASAP7_75t_L g164 ( .A(n_91), .Y(n_164) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_92), .A2(n_159), .B(n_161), .Y(n_158) );
BUFx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_93), .Y(n_121) );
INVx3_ASAP7_75t_L g189 ( .A(n_93), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_93), .A2(n_267), .B(n_268), .Y(n_266) );
BUFx12f_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx5_ASAP7_75t_L g128 ( .A(n_94), .Y(n_128) );
INVx5_ASAP7_75t_L g143 ( .A(n_94), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_94), .A2(n_201), .B(n_202), .C(n_203), .Y(n_200) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_381), .Y(n_98) );
NOR3xp33_ASAP7_75t_L g99 ( .A(n_100), .B(n_302), .C(n_346), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g100 ( .A(n_101), .B(n_276), .Y(n_100) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_195), .B(n_237), .Y(n_101) );
NAND2x1_ASAP7_75t_SL g102 ( .A(n_103), .B(n_172), .Y(n_102) );
OAI221xp5_ASAP7_75t_L g237 ( .A1(n_103), .A2(n_238), .B1(n_246), .B2(n_253), .C(n_258), .Y(n_237) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_131), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_107), .B(n_176), .Y(n_393) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g179 ( .A(n_108), .Y(n_179) );
INVx1_ASAP7_75t_L g252 ( .A(n_108), .Y(n_252) );
AND2x2_ASAP7_75t_L g293 ( .A(n_108), .B(n_180), .Y(n_293) );
AND2x2_ASAP7_75t_L g322 ( .A(n_108), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g341 ( .A(n_108), .B(n_132), .Y(n_341) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_108), .Y(n_358) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_115), .B(n_130), .Y(n_108) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_109), .A2(n_262), .B(n_270), .Y(n_261) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_109), .A2(n_262), .B(n_270), .Y(n_280) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx4_ASAP7_75t_L g133 ( .A(n_111), .Y(n_133) );
BUFx4f_ASAP7_75t_L g182 ( .A(n_111), .Y(n_182) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_111), .A2(n_217), .B(n_225), .Y(n_216) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_111), .A2(n_217), .B(n_225), .Y(n_240) );
OA21x2_ASAP7_75t_L g271 ( .A1(n_111), .A2(n_217), .B(n_225), .Y(n_271) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g212 ( .A(n_112), .Y(n_212) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g171 ( .A(n_113), .Y(n_171) );
OAI21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_122), .B(n_129), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_120), .B(n_121), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_118), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g147 ( .A(n_119), .Y(n_147) );
INVx1_ASAP7_75t_L g209 ( .A(n_119), .Y(n_209) );
OAI21xp33_ASAP7_75t_L g144 ( .A1(n_121), .A2(n_145), .B(n_148), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B(n_127), .Y(n_122) );
INVx2_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
INVx2_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_125), .B(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g207 ( .A(n_125), .Y(n_207) );
INVx2_ASAP7_75t_L g231 ( .A(n_125), .Y(n_231) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_128), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21x1_ASAP7_75t_L g263 ( .A1(n_128), .A2(n_264), .B(n_265), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_129), .A2(n_184), .B(n_190), .Y(n_183) );
OAI21x1_ASAP7_75t_L g199 ( .A1(n_129), .A2(n_200), .B(n_204), .Y(n_199) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_129), .A2(n_218), .B(n_222), .Y(n_217) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_129), .A2(n_229), .B(n_233), .Y(n_228) );
AND2x2_ASAP7_75t_L g309 ( .A(n_131), .B(n_289), .Y(n_309) );
INVx2_ASAP7_75t_L g356 ( .A(n_131), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_131), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g427 ( .A(n_131), .B(n_293), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_131), .B(n_312), .Y(n_443) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_153), .Y(n_131) );
AND2x2_ASAP7_75t_L g330 ( .A(n_132), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g432 ( .A(n_132), .B(n_181), .Y(n_432) );
AO21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B(n_152), .Y(n_132) );
INVx3_ASAP7_75t_L g156 ( .A(n_133), .Y(n_156) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_133), .A2(n_134), .B(n_152), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_138), .B(n_142), .Y(n_135) );
NOR2xp67_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
CKINVDCx6p67_ASAP7_75t_R g193 ( .A(n_143), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
NOR2xp33_ASAP7_75t_SL g148 ( .A(n_149), .B(n_151), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_149), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g174 ( .A(n_153), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g323 ( .A(n_153), .Y(n_323) );
INVx1_ASAP7_75t_L g331 ( .A(n_153), .Y(n_331) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g249 ( .A(n_154), .Y(n_249) );
AOI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_169), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_165), .Y(n_157) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx5_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_177), .Y(n_173) );
AND2x4_ASAP7_75t_L g300 ( .A(n_174), .B(n_293), .Y(n_300) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_175), .Y(n_377) );
INVx2_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_176), .B(n_180), .Y(n_274) );
INVx1_ASAP7_75t_L g321 ( .A(n_176), .Y(n_321) );
INVx1_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g289 ( .A(n_178), .Y(n_289) );
OR2x2_ASAP7_75t_L g301 ( .A(n_178), .B(n_247), .Y(n_301) );
OR2x2_ASAP7_75t_L g374 ( .A(n_178), .B(n_344), .Y(n_374) );
OR2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
BUFx3_ASAP7_75t_L g405 ( .A(n_180), .Y(n_405) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g251 ( .A(n_181), .Y(n_251) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_194), .Y(n_181) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_182), .A2(n_199), .B(n_210), .Y(n_198) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_182), .A2(n_228), .B(n_236), .Y(n_227) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_182), .A2(n_228), .B(n_236), .Y(n_245) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_182), .A2(n_199), .B(n_210), .Y(n_257) );
O2A1O1Ixp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .C(n_189), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_189), .A2(n_205), .B(n_206), .C(n_208), .Y(n_204) );
O2A1O1Ixp5_ASAP7_75t_L g233 ( .A1(n_189), .A2(n_206), .B(n_234), .C(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_193), .A2(n_219), .B(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_193), .A2(n_230), .B(n_232), .Y(n_229) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_213), .Y(n_195) );
INVx1_ASAP7_75t_L g364 ( .A(n_196), .Y(n_364) );
OAI32xp33_ASAP7_75t_L g373 ( .A1(n_196), .A2(n_374), .A3(n_375), .B1(n_378), .B2(n_379), .Y(n_373) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2x1_ASAP7_75t_L g241 ( .A(n_197), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_197), .B(n_226), .Y(n_308) );
AND2x4_ASAP7_75t_SL g397 ( .A(n_197), .B(n_388), .Y(n_397) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g316 ( .A(n_198), .Y(n_316) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_198), .Y(n_380) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_214), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_215), .B(n_226), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_216), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g284 ( .A(n_216), .B(n_243), .Y(n_284) );
INVx1_ASAP7_75t_L g440 ( .A(n_226), .Y(n_440) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g335 ( .A(n_227), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
OR2x2_ASAP7_75t_L g295 ( .A(n_239), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g333 ( .A(n_239), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_SL g306 ( .A(n_240), .Y(n_306) );
INVx2_ASAP7_75t_SL g345 ( .A(n_240), .Y(n_345) );
BUFx2_ASAP7_75t_L g360 ( .A(n_240), .Y(n_360) );
INVx1_ASAP7_75t_L g412 ( .A(n_241), .Y(n_412) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_243), .B(n_336), .Y(n_348) );
OR2x2_ASAP7_75t_L g353 ( .A(n_243), .B(n_345), .Y(n_353) );
AND2x2_ASAP7_75t_L g389 ( .A(n_243), .B(n_257), .Y(n_389) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g297 ( .A(n_244), .B(n_279), .Y(n_297) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g361 ( .A(n_245), .B(n_279), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
OR2x2_ASAP7_75t_L g454 ( .A(n_247), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g372 ( .A(n_248), .B(n_341), .Y(n_372) );
AND2x2_ASAP7_75t_L g435 ( .A(n_248), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g275 ( .A(n_249), .Y(n_275) );
INVxp67_ASAP7_75t_SL g288 ( .A(n_249), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_249), .B(n_251), .Y(n_409) );
INVx1_ASAP7_75t_L g425 ( .A(n_250), .Y(n_425) );
INVx1_ASAP7_75t_L g455 ( .A(n_250), .Y(n_455) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g319 ( .A(n_251), .Y(n_319) );
OR2x2_ASAP7_75t_L g357 ( .A(n_251), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_251), .B(n_275), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_251), .B(n_321), .Y(n_418) );
INVx1_ASAP7_75t_L g312 ( .A(n_252), .Y(n_312) );
INVxp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g368 ( .A(n_254), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx2_ASAP7_75t_L g452 ( .A(n_256), .Y(n_452) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g278 ( .A(n_257), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g326 ( .A(n_257), .B(n_261), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_272), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_271), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_260), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_260), .B(n_345), .Y(n_416) );
BUFx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B(n_269), .Y(n_262) );
NOR3xp33_ASAP7_75t_L g313 ( .A(n_271), .B(n_309), .C(n_314), .Y(n_313) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_271), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g402 ( .A(n_271), .Y(n_402) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_271), .Y(n_423) );
AND2x2_ASAP7_75t_L g428 ( .A(n_271), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g311 ( .A(n_273), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B1(n_294), .B2(n_298), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_277), .A2(n_407), .B1(n_410), .B2(n_412), .C(n_413), .Y(n_406) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g343 ( .A(n_278), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g336 ( .A(n_279), .Y(n_336) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .B1(n_290), .B2(n_292), .Y(n_281) );
NOR2xp67_ASAP7_75t_SL g437 ( .A(n_282), .B(n_351), .Y(n_437) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g396 ( .A(n_284), .Y(n_396) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_286), .A2(n_350), .B1(n_354), .B2(n_359), .Y(n_349) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
OR2x2_ASAP7_75t_L g420 ( .A(n_287), .B(n_357), .Y(n_420) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp67_ASAP7_75t_L g329 ( .A(n_293), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g365 ( .A(n_293), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g430 ( .A(n_293), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g314 ( .A(n_297), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g363 ( .A(n_297), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g459 ( .A(n_297), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_300), .A2(n_447), .B1(n_449), .B2(n_451), .C(n_453), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_313), .B1(n_317), .B2(n_324), .C(n_327), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .B(n_309), .C(n_310), .Y(n_303) );
AND2x2_ASAP7_75t_L g462 ( .A(n_305), .B(n_351), .Y(n_462) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_SL g414 ( .A(n_307), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI211xp5_ASAP7_75t_L g346 ( .A1(n_311), .A2(n_347), .B(n_349), .C(n_362), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_312), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g424 ( .A(n_315), .B(n_361), .Y(n_424) );
AND2x4_ASAP7_75t_L g467 ( .A(n_315), .B(n_388), .Y(n_467) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x4_ASAP7_75t_L g339 ( .A(n_319), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g456 ( .A(n_319), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
BUFx2_ASAP7_75t_SL g400 ( .A(n_321), .Y(n_400) );
INVx1_ASAP7_75t_L g419 ( .A(n_322), .Y(n_419) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g352 ( .A(n_326), .Y(n_352) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_332), .B1(n_337), .B2(n_342), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g441 ( .A(n_330), .B(n_404), .Y(n_441) );
INVx1_ASAP7_75t_L g457 ( .A(n_330), .Y(n_457) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_333), .A2(n_414), .B1(n_417), .B2(n_420), .Y(n_413) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g388 ( .A(n_336), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_337), .A2(n_462), .B1(n_463), .B2(n_464), .C(n_468), .Y(n_461) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g463 ( .A(n_339), .B(n_367), .Y(n_463) );
AND2x2_ASAP7_75t_L g410 ( .A(n_340), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g378 ( .A(n_341), .B(n_367), .Y(n_378) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g466 ( .A(n_344), .Y(n_466) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g379 ( .A(n_348), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g429 ( .A(n_348), .Y(n_429) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2x1_ASAP7_75t_SL g445 ( .A(n_352), .B(n_353), .Y(n_445) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g460 ( .A(n_360), .Y(n_460) );
INVx1_ASAP7_75t_L g370 ( .A(n_361), .Y(n_370) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_361), .B(n_452), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B1(n_368), .B2(n_371), .C(n_373), .Y(n_362) );
AOI222xp33_ASAP7_75t_L g426 ( .A1(n_363), .A2(n_386), .B1(n_427), .B2(n_428), .C1(n_430), .C2(n_432), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_366), .B(n_422), .C(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g450 ( .A(n_366), .Y(n_450) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_369), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_369), .B(n_410), .Y(n_469) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI21xp33_ASAP7_75t_L g449 ( .A1(n_374), .A2(n_391), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g431 ( .A(n_376), .Y(n_431) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_378), .A2(n_443), .B(n_444), .Y(n_442) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_380), .Y(n_448) );
NOR2xp33_ASAP7_75t_SL g381 ( .A(n_382), .B(n_433), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_406), .C(n_421), .D(n_426), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_390), .B(n_394), .Y(n_383) );
INVxp33_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
OR2x2_ASAP7_75t_L g408 ( .A(n_393), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g436 ( .A(n_393), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_398), .B1(n_401), .B2(n_403), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
AND2x4_ASAP7_75t_L g447 ( .A(n_396), .B(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_409), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g439 ( .A(n_416), .B(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_446), .C(n_461), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_438), .B2(n_441), .C(n_442), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI21xp33_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_456), .B(n_458), .Y(n_453) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVxp33_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B1(n_639), .B2(n_646), .C(n_689), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_473), .A2(n_690), .B1(n_694), .B2(n_695), .Y(n_689) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND3x1_ASAP7_75t_SL g474 ( .A(n_475), .B(n_529), .C(n_601), .Y(n_474) );
OAI31xp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_496), .A3(n_514), .B(n_524), .Y(n_475) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g498 ( .A(n_479), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g504 ( .A(n_479), .Y(n_504) );
AND2x6_ASAP7_75t_L g516 ( .A(n_479), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x6_ASAP7_75t_L g511 ( .A(n_480), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_481), .Y(n_490) );
INVx1_ASAP7_75t_L g521 ( .A(n_481), .Y(n_521) );
AND2x2_ASAP7_75t_L g581 ( .A(n_481), .B(n_526), .Y(n_581) );
INVx2_ASAP7_75t_L g595 ( .A(n_481), .Y(n_595) );
INVx2_ASAP7_75t_L g584 ( .A(n_482), .Y(n_584) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
AND2x2_ASAP7_75t_L g587 ( .A(n_483), .B(n_485), .Y(n_587) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g523 ( .A(n_484), .B(n_495), .Y(n_523) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_L g517 ( .A(n_486), .B(n_493), .Y(n_517) );
INVx4_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
AND2x4_ASAP7_75t_L g506 ( .A(n_489), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g512 ( .A(n_492), .Y(n_512) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g501 ( .A(n_493), .B(n_495), .Y(n_501) );
INVx1_ASAP7_75t_L g509 ( .A(n_494), .Y(n_509) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g503 ( .A(n_500), .B(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
CKINVDCx8_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_510), .B1(n_511), .B2(n_513), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g676 ( .A(n_509), .Y(n_676) );
AOI222xp33_ASAP7_75t_L g603 ( .A1(n_510), .A2(n_513), .B1(n_598), .B2(n_604), .C1(n_608), .C2(n_611), .Y(n_603) );
CKINVDCx6p67_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g589 ( .A(n_517), .Y(n_589) );
INVx4_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_522), .Y(n_590) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_523), .Y(n_600) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g594 ( .A(n_526), .B(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g554 ( .A(n_528), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_552), .B1(n_559), .B2(n_570), .C(n_578), .Y(n_529) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_532), .Y(n_564) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_533), .B(n_537), .Y(n_631) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g540 ( .A(n_534), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_534), .B(n_537), .Y(n_546) );
INVx1_ASAP7_75t_L g551 ( .A(n_534), .Y(n_551) );
INVx1_ASAP7_75t_L g607 ( .A(n_534), .Y(n_607) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g541 ( .A(n_537), .Y(n_541) );
INVx1_ASAP7_75t_L g550 ( .A(n_537), .Y(n_550) );
INVx1_ASAP7_75t_L g610 ( .A(n_537), .Y(n_610) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_SL g561 ( .A(n_539), .Y(n_561) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g635 ( .A(n_540), .Y(n_635) );
AND2x4_ASAP7_75t_L g606 ( .A(n_541), .B(n_607), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_547), .B2(n_548), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g582 ( .A1(n_543), .A2(n_547), .B1(n_583), .B2(n_585), .C(n_588), .Y(n_582) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g568 ( .A(n_545), .Y(n_568) );
OR2x6_ASAP7_75t_L g618 ( .A(n_545), .B(n_609), .Y(n_618) );
OR2x6_ASAP7_75t_L g621 ( .A(n_545), .B(n_622), .Y(n_621) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp33_ASAP7_75t_SL g565 ( .A1(n_548), .A2(n_566), .B1(n_567), .B2(n_569), .Y(n_565) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
BUFx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
OR2x2_ASAP7_75t_L g579 ( .A(n_554), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_556), .Y(n_638) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g609 ( .A(n_558), .Y(n_609) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx6_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x6_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g615 ( .A(n_575), .Y(n_615) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g623 ( .A(n_576), .Y(n_623) );
OAI22xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_582), .B1(n_591), .B2(n_596), .Y(n_578) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_SL g672 ( .A(n_581), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_583), .A2(n_585), .B1(n_597), .B2(n_598), .C(n_599), .Y(n_596) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x6_ASAP7_75t_L g637 ( .A(n_593), .B(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g682 ( .A(n_595), .B(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_597), .A2(n_617), .B1(n_619), .B2(n_620), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_627), .B(n_636), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_616), .C(n_624), .Y(n_602) );
BUFx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g625 ( .A(n_606), .B(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AND2x4_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g626 ( .A(n_615), .Y(n_626) );
INVx8_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx4_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g629 ( .A(n_622), .Y(n_629) );
AND2x4_ASAP7_75t_L g633 ( .A(n_622), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
CKINVDCx11_ASAP7_75t_R g624 ( .A(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
BUFx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx5_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
CKINVDCx16_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
BUFx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_643), .B(n_645), .Y(n_668) );
INVx1_ASAP7_75t_SL g697 ( .A(n_643), .Y(n_697) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_664), .B1(n_686), .B2(n_687), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_647), .A2(n_686), .B1(n_691), .B2(n_692), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_653), .B1(n_662), .B2(n_663), .Y(n_647) );
INVx1_ASAP7_75t_L g662 ( .A(n_648), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_648) );
CKINVDCx16_ASAP7_75t_R g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_651), .Y(n_652) );
INVx1_ASAP7_75t_L g663 ( .A(n_653), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_660), .B2(n_661), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx8_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx8_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
CKINVDCx20_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_667), .Y(n_691) );
OR2x6_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
OR2x4_ASAP7_75t_L g688 ( .A(n_668), .B(n_670), .Y(n_688) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI31xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .A3(n_677), .B(n_679), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g685 ( .A(n_676), .Y(n_685) );
INVx6_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVxp67_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx8_ASAP7_75t_L g693 ( .A(n_688), .Y(n_693) );
INVx8_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
endmodule