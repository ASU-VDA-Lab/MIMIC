module fake_netlist_5_976_n_1964 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1964);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1964;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_1058;
wire n_586;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_980;
wire n_698;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_SL g199 ( 
.A(n_72),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_113),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_57),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_14),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_73),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_97),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_172),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_108),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_60),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_104),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_32),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_47),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_75),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_155),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_118),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_70),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_141),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_38),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_42),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_76),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_10),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_112),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_45),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_22),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_109),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_71),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_106),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_196),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_142),
.Y(n_238)
);

INVxp33_ASAP7_75t_R g239 ( 
.A(n_9),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_63),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_61),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_77),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_115),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_138),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_105),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_42),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_13),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_86),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_23),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_80),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_156),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_88),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_177),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_82),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_191),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_102),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_48),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_146),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_14),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_79),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_10),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_46),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_190),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_69),
.Y(n_267)
);

BUFx2_ASAP7_75t_SL g268 ( 
.A(n_2),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_160),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_84),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_83),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_182),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_68),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_145),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_44),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_56),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_3),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_148),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_157),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_62),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_192),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_12),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_60),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_135),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_67),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_147),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_64),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_92),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_59),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_161),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_95),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_144),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_51),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_26),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_37),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_91),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_178),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_40),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_27),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_53),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_51),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_128),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_131),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_185),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_126),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_54),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_64),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_85),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_151),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_100),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_169),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_24),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_28),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_165),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_15),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_16),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_29),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_0),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_43),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_96),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_99),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_54),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_197),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_67),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_25),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_111),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_13),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_49),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_44),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_98),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_170),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_87),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_21),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_124),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_59),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_35),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_120),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_194),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_183),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_81),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_19),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_195),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_123),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_34),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_89),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_116),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_184),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_78),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_53),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_137),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_43),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_133),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_187),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_121),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_18),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_164),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_122),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_46),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_62),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_57),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_25),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_7),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_32),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_134),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_140),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_93),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_38),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_36),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_139),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_37),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_20),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_176),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_74),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_41),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_174),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_129),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_167),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_90),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_119),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_1),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_1),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_130),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_26),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_16),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_6),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_136),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_63),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_55),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_94),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_153),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_179),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_110),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_27),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_2),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_0),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_302),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_301),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_207),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_235),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_302),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_302),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_206),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_337),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_248),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_264),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_332),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_211),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_301),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_243),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_210),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_301),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_251),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_301),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_301),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_304),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_304),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_253),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_277),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_259),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_265),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_294),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_276),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_300),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_342),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_352),
.Y(n_429)
);

BUFx10_ASAP7_75t_L g430 ( 
.A(n_304),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_279),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_304),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_304),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_383),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_315),
.Y(n_435)
);

INVxp33_ASAP7_75t_SL g436 ( 
.A(n_215),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_283),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_315),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_280),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_285),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_390),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_286),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_280),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_288),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_303),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_303),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_315),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_315),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_315),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_229),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_215),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_388),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_290),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_305),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_377),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_388),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_247),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_298),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_310),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_201),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_202),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_232),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_241),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_217),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_249),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_260),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_296),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_274),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_278),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_252),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_254),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_296),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_295),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_292),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_322),
.Y(n_478)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_296),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_217),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_322),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_255),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_345),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_220),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_345),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_348),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_220),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_316),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_257),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_295),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_348),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_226),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_297),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_318),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_311),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_397),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_309),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_214),
.Y(n_499)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_329),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_319),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_333),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_364),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_321),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_499),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_457),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_438),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_476),
.B(n_200),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_438),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_473),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_200),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_499),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_447),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_401),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_447),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_499),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_214),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_423),
.B(n_204),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_496),
.B(n_311),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_499),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_313),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_439),
.B(n_340),
.Y(n_525)
);

BUFx12f_ASAP7_75t_L g526 ( 
.A(n_408),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_448),
.B(n_205),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_443),
.B(n_340),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_415),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_406),
.B(n_313),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_417),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_418),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_414),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_419),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_420),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_411),
.B(n_199),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_420),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_432),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_400),
.B(n_334),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_432),
.B(n_214),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_433),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_445),
.B(n_334),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_433),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_449),
.B(n_205),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_456),
.B(n_208),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_450),
.B(n_219),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_435),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_454),
.B(n_455),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_446),
.B(n_458),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_435),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_452),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_430),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_452),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_459),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_462),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_408),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_421),
.B(n_320),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_404),
.B(n_208),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_502),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_405),
.A2(n_368),
.B(n_231),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_430),
.B(n_209),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_430),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_502),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_474),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_478),
.B(n_231),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_436),
.B(n_245),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_467),
.B(n_338),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_478),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_481),
.B(n_214),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_482),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_463),
.B(n_204),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_494),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_481),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_483),
.B(n_214),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_416),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_498),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_498),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_464),
.B(n_209),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_416),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_409),
.A2(n_359),
.B1(n_353),
.B2(n_387),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_483),
.Y(n_586)
);

NOR2x1p5_ASAP7_75t_L g587 ( 
.A(n_526),
.B(n_226),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_509),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_566),
.B(n_424),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_507),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_509),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_507),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_508),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_537),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_507),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_515),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_513),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_515),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_540),
.A2(n_385),
.B1(n_410),
.B2(n_407),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_R g600 ( 
.A(n_506),
.B(n_511),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_546),
.B(n_485),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_530),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_517),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_519),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_510),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_517),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_556),
.Y(n_608)
);

BUFx4f_ASAP7_75t_L g609 ( 
.A(n_564),
.Y(n_609)
);

BUFx4f_ASAP7_75t_L g610 ( 
.A(n_564),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_510),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_523),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_513),
.Y(n_614)
);

INVx8_ASAP7_75t_L g615 ( 
.A(n_519),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_550),
.A2(n_230),
.B1(n_233),
.B2(n_227),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_566),
.B(n_424),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_523),
.Y(n_618)
);

AOI22x1_ASAP7_75t_L g619 ( 
.A1(n_525),
.A2(n_480),
.B1(n_484),
.B2(n_451),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_513),
.Y(n_620)
);

BUFx4f_ASAP7_75t_L g621 ( 
.A(n_564),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_510),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_570),
.B(n_493),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_514),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_514),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_513),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_514),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_516),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_516),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_513),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_516),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_536),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_565),
.B(n_426),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_527),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_546),
.B(n_485),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_571),
.B(n_426),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_508),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_512),
.B(n_431),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_522),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_532),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_562),
.B(n_466),
.C(n_465),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_512),
.B(n_431),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_L g643 ( 
.A1(n_531),
.A2(n_323),
.B1(n_328),
.B2(n_326),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_536),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_532),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_556),
.B(n_437),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_556),
.B(n_437),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_533),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_552),
.B(n_204),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_536),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_L g651 ( 
.A(n_578),
.B(n_258),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_565),
.B(n_440),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_533),
.Y(n_653)
);

INVx8_ASAP7_75t_L g654 ( 
.A(n_519),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_520),
.B(n_490),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_534),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_528),
.B(n_440),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_530),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_526),
.B(n_268),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_584),
.B(n_442),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_534),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_538),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_576),
.B(n_444),
.Y(n_663)
);

AND2x2_ASAP7_75t_SL g664 ( 
.A(n_564),
.B(n_368),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_561),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_541),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_541),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_541),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_576),
.B(n_444),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_530),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_530),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_538),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_539),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_521),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_522),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_547),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_R g677 ( 
.A(n_568),
.B(n_402),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_547),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_543),
.A2(n_366),
.B1(n_389),
.B2(n_372),
.Y(n_679)
);

BUFx4f_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_547),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_575),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_526),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_543),
.B(n_486),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_561),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_583),
.B(n_453),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_543),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_555),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_585),
.A2(n_479),
.B1(n_475),
.B2(n_403),
.Y(n_689)
);

AND2x2_ASAP7_75t_SL g690 ( 
.A(n_560),
.B(n_379),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_543),
.B(n_486),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_555),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_539),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_583),
.A2(n_375),
.B1(n_384),
.B2(n_378),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_522),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_528),
.B(n_548),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_530),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_569),
.B(n_379),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_548),
.B(n_549),
.Y(n_700)
);

AND2x6_ASAP7_75t_L g701 ( 
.A(n_525),
.B(n_269),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_557),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_557),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_524),
.B(n_453),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_562),
.B(n_469),
.C(n_468),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_580),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_549),
.B(n_460),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_505),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_529),
.B(n_460),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_557),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_522),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_542),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_542),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_505),
.B(n_461),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_553),
.B(n_461),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_522),
.Y(n_716)
);

INVxp33_ASAP7_75t_L g717 ( 
.A(n_585),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_551),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_529),
.B(n_488),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_551),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_554),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_505),
.B(n_488),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_554),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_530),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_559),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_559),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_505),
.B(n_495),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_569),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_573),
.B(n_472),
.C(n_471),
.Y(n_729)
);

BUFx6f_ASAP7_75t_SL g730 ( 
.A(n_569),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_559),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_569),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_535),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_559),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_535),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_573),
.B(n_495),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_518),
.B(n_501),
.Y(n_737)
);

AND2x4_ASAP7_75t_SL g738 ( 
.A(n_659),
.B(n_413),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_697),
.A2(n_577),
.B(n_582),
.C(n_581),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_609),
.A2(n_522),
.B(n_518),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_594),
.Y(n_741)
);

NAND2x1_ASAP7_75t_L g742 ( 
.A(n_597),
.B(n_519),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_649),
.A2(n_500),
.B1(n_398),
.B2(n_262),
.Y(n_743)
);

NAND2x1_ASAP7_75t_L g744 ( 
.A(n_597),
.B(n_519),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_594),
.B(n_501),
.Y(n_745)
);

INVxp33_ASAP7_75t_L g746 ( 
.A(n_613),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_590),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_590),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_593),
.B(n_567),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_593),
.B(n_567),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_637),
.B(n_567),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_690),
.B(n_269),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_637),
.B(n_567),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_687),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_592),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_623),
.B(n_504),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_592),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_687),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_700),
.B(n_567),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_674),
.B(n_504),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_613),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_719),
.B(n_487),
.Y(n_762)
);

INVxp33_ASAP7_75t_L g763 ( 
.A(n_677),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_690),
.B(n_269),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_602),
.B(n_577),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_674),
.B(n_578),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_690),
.B(n_269),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_736),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_638),
.B(n_642),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_728),
.B(n_578),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_684),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_728),
.B(n_578),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_732),
.B(n_535),
.Y(n_773)
);

INVx8_ASAP7_75t_L g774 ( 
.A(n_730),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_649),
.B(n_470),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_732),
.A2(n_422),
.B1(n_425),
.B2(n_427),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_706),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_657),
.B(n_704),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_664),
.B(n_535),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_715),
.B(n_589),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_665),
.B(n_489),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_602),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_684),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_609),
.A2(n_336),
.B(n_213),
.C(n_216),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_691),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_664),
.B(n_535),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_707),
.A2(n_582),
.B(n_581),
.C(n_477),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_595),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_609),
.B(n_610),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_664),
.B(n_535),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_636),
.B(n_497),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_686),
.B(n_212),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_709),
.B(n_212),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_617),
.B(n_218),
.Y(n_794)
);

NAND3xp33_ASAP7_75t_L g795 ( 
.A(n_633),
.B(n_221),
.C(n_218),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_635),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_588),
.B(n_545),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_635),
.B(n_428),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_610),
.B(n_269),
.Y(n_799)
);

NAND2x1p5_ASAP7_75t_L g800 ( 
.A(n_605),
.B(n_608),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_691),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_588),
.B(n_545),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_606),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_706),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_591),
.B(n_545),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_591),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_596),
.B(n_545),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_606),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_652),
.A2(n_429),
.B1(n_434),
.B2(n_441),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_596),
.B(n_545),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_663),
.B(n_221),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_611),
.Y(n_812)
);

OAI22xp33_ASAP7_75t_L g813 ( 
.A1(n_717),
.A2(n_233),
.B1(n_230),
.B2(n_331),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_598),
.B(n_545),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_610),
.B(n_203),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_598),
.B(n_518),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_L g817 ( 
.A(n_701),
.B(n_261),
.Y(n_817)
);

OA22x2_ASAP7_75t_L g818 ( 
.A1(n_616),
.A2(n_227),
.B1(n_240),
.B2(n_374),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_604),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_611),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_615),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_665),
.B(n_503),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_622),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_604),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_607),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_622),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_607),
.B(n_558),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_669),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_612),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_612),
.B(n_558),
.Y(n_830)
);

AO22x2_ASAP7_75t_L g831 ( 
.A1(n_660),
.A2(n_242),
.B1(n_244),
.B2(n_396),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_618),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_621),
.B(n_222),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_726),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_621),
.B(n_223),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_737),
.B(n_225),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_621),
.A2(n_327),
.B1(n_267),
.B2(n_395),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_608),
.B(n_503),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_695),
.B(n_224),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_714),
.Y(n_840)
);

OAI22xp33_ASAP7_75t_L g841 ( 
.A1(n_616),
.A2(n_355),
.B1(n_339),
.B2(n_240),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_730),
.A2(n_271),
.B1(n_263),
.B2(n_266),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_624),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_634),
.B(n_640),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_634),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_655),
.B(n_563),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_624),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_625),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_682),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_722),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_727),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_625),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_646),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_627),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_640),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_627),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_645),
.B(n_558),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_641),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_641),
.Y(n_859)
);

AND2x6_ASAP7_75t_L g860 ( 
.A(n_699),
.B(n_228),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_628),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_648),
.B(n_558),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_699),
.B(n_246),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_685),
.B(n_331),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_685),
.B(n_339),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_647),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_699),
.B(n_250),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_599),
.B(n_225),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_648),
.B(n_558),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_730),
.A2(n_275),
.B1(n_270),
.B2(n_272),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_628),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_699),
.B(n_605),
.Y(n_872)
);

NOR2x1p5_ASAP7_75t_L g873 ( 
.A(n_683),
.B(n_355),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_643),
.B(n_234),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_653),
.B(n_558),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_656),
.B(n_256),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_619),
.Y(n_877)
);

BUFx5_ASAP7_75t_L g878 ( 
.A(n_726),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_605),
.B(n_306),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_661),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_661),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_701),
.A2(n_386),
.B1(n_370),
.B2(n_346),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_662),
.B(n_234),
.Y(n_883)
);

AND2x6_ASAP7_75t_SL g884 ( 
.A(n_659),
.B(n_239),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_629),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_672),
.B(n_344),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_672),
.B(n_376),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_673),
.B(n_381),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_629),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_705),
.B(n_563),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_694),
.B(n_382),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_631),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_694),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_712),
.B(n_236),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_619),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_631),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_605),
.B(n_394),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_701),
.A2(n_365),
.B1(n_367),
.B2(n_363),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_712),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_713),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_899),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_762),
.B(n_745),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_769),
.B(n_713),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_741),
.Y(n_904)
);

AOI22x1_ASAP7_75t_L g905 ( 
.A1(n_806),
.A2(n_824),
.B1(n_825),
.B2(n_819),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_769),
.B(n_689),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_747),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_899),
.Y(n_908)
);

BUFx12f_ASAP7_75t_L g909 ( 
.A(n_884),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_829),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_759),
.B(n_720),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_832),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_796),
.B(n_659),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_849),
.Y(n_914)
);

OR2x6_ASAP7_75t_L g915 ( 
.A(n_774),
.B(n_777),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_840),
.B(n_720),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_840),
.B(n_718),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_850),
.B(n_718),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_851),
.B(n_721),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_752),
.A2(n_701),
.B1(n_721),
.B2(n_723),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_782),
.B(n_659),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_768),
.B(n_844),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_768),
.B(n_723),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_858),
.B(n_725),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_771),
.B(n_659),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_779),
.A2(n_680),
.B(n_654),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_748),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_783),
.B(n_587),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_853),
.B(n_866),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_778),
.B(n_651),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_821),
.B(n_605),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_785),
.B(n_587),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_822),
.B(n_682),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_758),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_845),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_756),
.B(n_708),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_846),
.B(n_600),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_752),
.A2(n_701),
.B1(n_708),
.B2(n_731),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_756),
.B(n_708),
.Y(n_939)
);

O2A1O1Ixp5_ASAP7_75t_L g940 ( 
.A1(n_764),
.A2(n_680),
.B(n_735),
.C(n_734),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_864),
.B(n_683),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_755),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_855),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_780),
.B(n_605),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_801),
.B(n_729),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_757),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_764),
.A2(n_701),
.B1(n_734),
.B2(n_731),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_836),
.B(n_679),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_821),
.B(n_733),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_836),
.B(n_733),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_860),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_798),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_789),
.A2(n_725),
.B(n_680),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_788),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_760),
.B(n_236),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_L g956 ( 
.A(n_741),
.B(n_729),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_761),
.B(n_397),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_761),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_858),
.B(n_735),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_746),
.B(n_237),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_880),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_758),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_881),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_781),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_758),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_838),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_786),
.A2(n_654),
.B(n_615),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_775),
.B(n_237),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_804),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_775),
.B(n_238),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_793),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_791),
.B(n_238),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_803),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_860),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_859),
.B(n_330),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_765),
.B(n_492),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_L g977 ( 
.A(n_758),
.B(n_615),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_893),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_900),
.B(n_601),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_804),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_766),
.B(n_754),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_774),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_808),
.Y(n_983)
);

INVx4_ASAP7_75t_SL g984 ( 
.A(n_860),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_789),
.A2(n_644),
.B(n_632),
.Y(n_985)
);

INVx8_ASAP7_75t_L g986 ( 
.A(n_774),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_790),
.B(n_632),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_776),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_816),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_812),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_754),
.B(n_890),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_820),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_823),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_809),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_791),
.B(n_335),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_799),
.A2(n_654),
.B(n_615),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_SL g997 ( 
.A(n_841),
.B(n_363),
.C(n_362),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_826),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_828),
.B(n_492),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_883),
.B(n_601),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_860),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_843),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_SL g1003 ( 
.A1(n_799),
.A2(n_666),
.B(n_650),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_767),
.A2(n_678),
.B1(n_666),
.B2(n_710),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_865),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_860),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_847),
.Y(n_1007)
);

AND2x2_ASAP7_75t_SL g1008 ( 
.A(n_738),
.B(n_289),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_828),
.B(n_335),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_868),
.B(n_362),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_877),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_868),
.B(n_365),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_895),
.B(n_341),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_848),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_SL g1015 ( 
.A1(n_792),
.A2(n_371),
.B1(n_367),
.B2(n_374),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_898),
.A2(n_391),
.B1(n_392),
.B2(n_399),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_831),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_872),
.B(n_603),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_852),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_742),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_883),
.B(n_601),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_854),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_856),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_749),
.B(n_650),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_873),
.B(n_615),
.Y(n_1025)
);

NOR2xp67_ASAP7_75t_L g1026 ( 
.A(n_795),
.B(n_792),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_750),
.B(n_667),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_898),
.A2(n_371),
.B1(n_391),
.B2(n_392),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_763),
.B(n_341),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_751),
.B(n_667),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_872),
.B(n_603),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_861),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_876),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_871),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_744),
.Y(n_1035)
);

NOR2x1p5_ASAP7_75t_L g1036 ( 
.A(n_753),
.B(n_399),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_885),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_811),
.B(n_343),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_889),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_874),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_831),
.A2(n_361),
.B1(n_343),
.B2(n_347),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_793),
.B(n_811),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_874),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_743),
.A2(n_360),
.B(n_347),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_794),
.B(n_614),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_743),
.B(n_349),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_894),
.B(n_620),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_892),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_896),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_R g1050 ( 
.A(n_817),
.B(n_349),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_815),
.A2(n_692),
.B(n_676),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_797),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_839),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_739),
.B(n_350),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_802),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_831),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_839),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_813),
.B(n_350),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_805),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_834),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_834),
.B(n_668),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_834),
.B(n_668),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_800),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_863),
.A2(n_675),
.B1(n_716),
.B2(n_626),
.Y(n_1064)
);

OAI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_886),
.A2(n_373),
.B1(n_351),
.B2(n_354),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_807),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_834),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_815),
.B(n_603),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_800),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_810),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_818),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_SL g1072 ( 
.A(n_841),
.B(n_393),
.C(n_373),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_863),
.A2(n_675),
.B1(n_716),
.B2(n_626),
.Y(n_1073)
);

AO21x2_ASAP7_75t_L g1074 ( 
.A1(n_833),
.A2(n_835),
.B(n_740),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_818),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_887),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_888),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_867),
.A2(n_675),
.B1(n_626),
.B2(n_620),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1042),
.B(n_842),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_987),
.A2(n_911),
.B(n_903),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_922),
.B(n_891),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_1038),
.A2(n_995),
.B(n_972),
.C(n_968),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_914),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_982),
.Y(n_1084)
);

OAI22x1_ASAP7_75t_L g1085 ( 
.A1(n_1043),
.A2(n_813),
.B1(n_870),
.B2(n_835),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_R g1086 ( 
.A(n_994),
.B(n_814),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_907),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_903),
.A2(n_833),
.B1(n_770),
.B2(n_772),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_987),
.A2(n_837),
.B(n_784),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_969),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_922),
.B(n_787),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_902),
.B(n_867),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_971),
.B(n_878),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_911),
.A2(n_773),
.B(n_875),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_948),
.A2(n_862),
.B(n_830),
.C(n_857),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_910),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_912),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_950),
.A2(n_1074),
.B(n_977),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_923),
.B(n_878),
.Y(n_1099)
);

AND2x2_ASAP7_75t_SL g1100 ( 
.A(n_1040),
.B(n_882),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_982),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_906),
.A2(n_827),
.B(n_869),
.C(n_879),
.Y(n_1102)
);

NOR2xp67_ASAP7_75t_L g1103 ( 
.A(n_933),
.B(n_879),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1076),
.B(n_878),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_927),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1077),
.B(n_917),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1074),
.A2(n_939),
.B(n_936),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1011),
.A2(n_688),
.B(n_678),
.C(n_703),
.Y(n_1108)
);

OA22x2_ASAP7_75t_L g1109 ( 
.A1(n_1071),
.A2(n_351),
.B1(n_393),
.B2(n_354),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_917),
.B(n_882),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_926),
.A2(n_981),
.B(n_1000),
.Y(n_1111)
);

O2A1O1Ixp5_ASAP7_75t_L g1112 ( 
.A1(n_1054),
.A2(n_897),
.B(n_692),
.C(n_688),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1026),
.A2(n_897),
.B1(n_273),
.B2(n_281),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_916),
.B(n_681),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_964),
.B(n_356),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1053),
.A2(n_282),
.B1(n_284),
.B2(n_287),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1033),
.B(n_356),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_982),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1021),
.A2(n_654),
.B(n_671),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_980),
.B(n_357),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1046),
.A2(n_360),
.B(n_369),
.C(n_361),
.Y(n_1121)
);

BUFx2_ASAP7_75t_R g1122 ( 
.A(n_952),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_985),
.A2(n_703),
.B(n_702),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_SL g1124 ( 
.A(n_986),
.B(n_289),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_916),
.B(n_681),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_SL g1126 ( 
.A(n_986),
.B(n_289),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_904),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_L g1128 ( 
.A(n_1058),
.B(n_369),
.C(n_357),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1047),
.A2(n_724),
.B(n_603),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_958),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_962),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_901),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_930),
.A2(n_693),
.B(n_702),
.C(n_724),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_908),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_967),
.A2(n_724),
.B(n_658),
.Y(n_1135)
);

OA22x2_ASAP7_75t_L g1136 ( 
.A1(n_1075),
.A2(n_291),
.B1(n_293),
.B2(n_299),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_970),
.A2(n_693),
.B(n_698),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_962),
.Y(n_1138)
);

NAND2x1_ASAP7_75t_L g1139 ( 
.A(n_1060),
.B(n_630),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_959),
.A2(n_572),
.B(n_586),
.C(n_358),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1061),
.A2(n_724),
.B(n_658),
.Y(n_1141)
);

NOR3xp33_ASAP7_75t_SL g1142 ( 
.A(n_1016),
.B(n_307),
.C(n_308),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1053),
.A2(n_312),
.B1(n_325),
.B2(n_314),
.Y(n_1143)
);

NOR2x1_ASAP7_75t_R g1144 ( 
.A(n_909),
.B(n_317),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1057),
.B(n_956),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1005),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1057),
.A2(n_988),
.B1(n_991),
.B2(n_1036),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_918),
.B(n_572),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_918),
.B(n_572),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_942),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_941),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_962),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_935),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1029),
.B(n_324),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_919),
.B(n_586),
.Y(n_1155)
);

INVx3_ASAP7_75t_SL g1156 ( 
.A(n_915),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1061),
.A2(n_586),
.B(n_698),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_919),
.B(n_380),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_946),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_966),
.B(n_658),
.Y(n_1160)
);

AOI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1062),
.A2(n_1027),
.B(n_1024),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_SL g1162 ( 
.A(n_986),
.B(n_358),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_959),
.A2(n_358),
.B(n_4),
.C(n_5),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_945),
.A2(n_696),
.B(n_639),
.C(n_630),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1010),
.B(n_658),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1062),
.A2(n_670),
.B(n_698),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1024),
.A2(n_670),
.B(n_698),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_915),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_954),
.Y(n_1169)
);

OA21x2_ASAP7_75t_L g1170 ( 
.A1(n_940),
.A2(n_670),
.B(n_671),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1017),
.A2(n_711),
.B(n_696),
.C(n_639),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1012),
.B(n_671),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_929),
.B(n_937),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_991),
.A2(n_671),
.B1(n_696),
.B2(n_711),
.Y(n_1174)
);

NOR3xp33_ASAP7_75t_SL g1175 ( 
.A(n_1016),
.B(n_1028),
.C(n_1044),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_L g1176 ( 
.A(n_934),
.B(n_630),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_989),
.B(n_711),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_924),
.B(n_711),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_924),
.B(n_639),
.Y(n_1179)
);

OR2x6_ASAP7_75t_SL g1180 ( 
.A(n_1028),
.B(n_3),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1027),
.A2(n_519),
.B(n_574),
.Y(n_1181)
);

AOI22x1_ASAP7_75t_L g1182 ( 
.A1(n_1052),
.A2(n_579),
.B1(n_574),
.B2(n_544),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1030),
.A2(n_519),
.B(n_574),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1056),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1068),
.A2(n_198),
.B1(n_193),
.B2(n_189),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_921),
.B(n_159),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_943),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_973),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1030),
.A2(n_996),
.B(n_953),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1013),
.A2(n_8),
.B(n_11),
.C(n_12),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_SL g1191 ( 
.A(n_1008),
.B(n_519),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_L g1192 ( 
.A(n_915),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_985),
.A2(n_544),
.B(n_579),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_961),
.B(n_15),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1068),
.A2(n_158),
.B1(n_152),
.B2(n_150),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_976),
.A2(n_579),
.B1(n_574),
.B2(n_544),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_913),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_928),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_963),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_976),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_978),
.A2(n_579),
.B1(n_574),
.B2(n_544),
.Y(n_1201)
);

AO21x1_ASAP7_75t_L g1202 ( 
.A1(n_1041),
.A2(n_17),
.B(n_21),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_983),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1022),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_999),
.B(n_22),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_925),
.B(n_149),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_960),
.B(n_23),
.Y(n_1207)
);

CKINVDCx16_ASAP7_75t_R g1208 ( 
.A(n_928),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_990),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1063),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1037),
.Y(n_1211)
);

AND3x2_ASAP7_75t_L g1212 ( 
.A(n_925),
.B(n_24),
.C(n_28),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_955),
.A2(n_932),
.B1(n_975),
.B2(n_1045),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1009),
.B(n_30),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_932),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1003),
.A2(n_544),
.B(n_579),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1049),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_953),
.A2(n_579),
.B(n_574),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1045),
.A2(n_544),
.B1(n_574),
.B2(n_579),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1055),
.B(n_30),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_951),
.B(n_143),
.Y(n_1221)
);

AO22x1_ASAP7_75t_L g1222 ( 
.A1(n_1041),
.A2(n_957),
.B1(n_965),
.B2(n_934),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1051),
.A2(n_544),
.B(n_132),
.Y(n_1223)
);

AOI221xp5_ASAP7_75t_L g1224 ( 
.A1(n_997),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.C(n_36),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1065),
.A2(n_117),
.B1(n_114),
.B2(n_107),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1059),
.B(n_31),
.Y(n_1226)
);

OR2x6_ASAP7_75t_L g1227 ( 
.A(n_1025),
.B(n_103),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1123),
.A2(n_1051),
.B(n_905),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1082),
.A2(n_1015),
.B(n_1072),
.C(n_1066),
.Y(n_1229)
);

BUFx8_ASAP7_75t_L g1230 ( 
.A(n_1083),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1080),
.A2(n_1001),
.B(n_951),
.Y(n_1231)
);

INVx3_ASAP7_75t_SL g1232 ( 
.A(n_1084),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1080),
.A2(n_1001),
.B(n_951),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1207),
.A2(n_1070),
.B(n_1002),
.C(n_1048),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1096),
.Y(n_1235)
);

NOR2xp67_ASAP7_75t_L g1236 ( 
.A(n_1173),
.B(n_965),
.Y(n_1236)
);

NAND3x1_ASAP7_75t_L g1237 ( 
.A(n_1147),
.B(n_1019),
.C(n_992),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1135),
.A2(n_1157),
.B(n_1141),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1146),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1222),
.A2(n_944),
.B(n_979),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1107),
.A2(n_1189),
.B(n_1098),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1106),
.B(n_1014),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1141),
.A2(n_949),
.B(n_1067),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_1132),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1154),
.B(n_1023),
.C(n_993),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1098),
.A2(n_1006),
.B(n_974),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1089),
.A2(n_1189),
.B(n_1111),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1210),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1197),
.B(n_1025),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1094),
.A2(n_1004),
.B(n_920),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1094),
.A2(n_947),
.B(n_938),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1081),
.B(n_1039),
.Y(n_1252)
);

BUFx4f_ASAP7_75t_L g1253 ( 
.A(n_1156),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1092),
.B(n_1025),
.Y(n_1254)
);

AOI21xp33_ASAP7_75t_L g1255 ( 
.A1(n_1140),
.A2(n_1032),
.B(n_998),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1111),
.A2(n_951),
.B(n_974),
.Y(n_1256)
);

BUFx8_ASAP7_75t_L g1257 ( 
.A(n_1198),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1127),
.Y(n_1258)
);

NOR2x1_ASAP7_75t_L g1259 ( 
.A(n_1210),
.B(n_1007),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_SL g1260 ( 
.A1(n_1202),
.A2(n_1078),
.B(n_1073),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1145),
.B(n_1034),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1131),
.Y(n_1262)
);

AND2x2_ASAP7_75t_SL g1263 ( 
.A(n_1100),
.B(n_1069),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1208),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1079),
.B(n_1069),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1131),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1091),
.B(n_1050),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1088),
.A2(n_974),
.B(n_1001),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1090),
.B(n_1069),
.Y(n_1269)
);

BUFx2_ASAP7_75t_R g1270 ( 
.A(n_1101),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1166),
.A2(n_1018),
.B(n_1031),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1151),
.B(n_1031),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1119),
.A2(n_974),
.B(n_1001),
.Y(n_1273)
);

OAI21xp33_ASAP7_75t_L g1274 ( 
.A1(n_1175),
.A2(n_1214),
.B(n_1224),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1165),
.B(n_1063),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1119),
.A2(n_1006),
.B(n_931),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1097),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1137),
.A2(n_1018),
.A3(n_1064),
.B(n_984),
.Y(n_1278)
);

OAI22x1_ASAP7_75t_L g1279 ( 
.A1(n_1213),
.A2(n_1006),
.B1(n_39),
.B2(n_40),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1130),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1172),
.A2(n_1006),
.B(n_1063),
.C(n_1020),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1086),
.B(n_984),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1110),
.A2(n_1035),
.B1(n_1020),
.B2(n_931),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1121),
.A2(n_33),
.B(n_39),
.C(n_41),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1131),
.Y(n_1285)
);

NAND3xp33_ASAP7_75t_SL g1286 ( 
.A(n_1124),
.B(n_45),
.C(n_47),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1095),
.A2(n_1035),
.B(n_101),
.Y(n_1287)
);

AOI221x1_ASAP7_75t_L g1288 ( 
.A1(n_1085),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.C(n_52),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1153),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1167),
.A2(n_55),
.B(n_56),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1114),
.B(n_58),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1223),
.A2(n_58),
.B(n_61),
.Y(n_1292)
);

AOI221xp5_ASAP7_75t_L g1293 ( 
.A1(n_1190),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.C(n_1163),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1118),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_SL g1295 ( 
.A(n_1122),
.B(n_65),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_1128),
.B(n_66),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1168),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1138),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1223),
.A2(n_1102),
.B(n_1133),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1138),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1167),
.A2(n_1129),
.B(n_1161),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1158),
.B(n_1125),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1180),
.A2(n_1099),
.B1(n_1093),
.B2(n_1226),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1142),
.A2(n_1103),
.B(n_1220),
.C(n_1190),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_SL g1306 ( 
.A1(n_1171),
.A2(n_1164),
.B(n_1104),
.C(n_1221),
.Y(n_1306)
);

AND2x6_ASAP7_75t_L g1307 ( 
.A(n_1138),
.B(n_1152),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1112),
.A2(n_1129),
.B(n_1178),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1152),
.Y(n_1309)
);

AND2x2_ASAP7_75t_SL g1310 ( 
.A(n_1192),
.B(n_1126),
.Y(n_1310)
);

AO22x2_ASAP7_75t_L g1311 ( 
.A1(n_1194),
.A2(n_1195),
.B1(n_1185),
.B2(n_1186),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1139),
.A2(n_1108),
.B(n_1183),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1209),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1155),
.B(n_1200),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1218),
.A2(n_1183),
.A3(n_1181),
.B(n_1179),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1087),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1177),
.B(n_1169),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1206),
.A2(n_1184),
.B(n_1187),
.C(n_1199),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1134),
.Y(n_1319)
);

BUFx4f_ASAP7_75t_L g1320 ( 
.A(n_1197),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1192),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1227),
.A2(n_1225),
.B1(n_1174),
.B2(n_1205),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1108),
.A2(n_1181),
.B(n_1218),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1140),
.A2(n_1216),
.B(n_1193),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1163),
.A2(n_1115),
.B(n_1113),
.C(n_1191),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1105),
.B(n_1188),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1117),
.A2(n_1120),
.B(n_1211),
.C(n_1204),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1109),
.A2(n_1136),
.B1(n_1217),
.B2(n_1203),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1109),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1150),
.A2(n_1159),
.B(n_1162),
.C(n_1143),
.Y(n_1330)
);

OAI22x1_ASAP7_75t_L g1331 ( 
.A1(n_1116),
.A2(n_1136),
.B1(n_1212),
.B2(n_1176),
.Y(n_1331)
);

AOI211x1_ASAP7_75t_L g1332 ( 
.A1(n_1227),
.A2(n_1152),
.B(n_1144),
.C(n_1160),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1160),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1227),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1170),
.A2(n_1219),
.B(n_1182),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1196),
.Y(n_1336)
);

OA22x2_ASAP7_75t_L g1337 ( 
.A1(n_1201),
.A2(n_1043),
.B1(n_613),
.B2(n_594),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1127),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1081),
.B(n_903),
.Y(n_1339)
);

AO221x2_ASAP7_75t_L g1340 ( 
.A1(n_1085),
.A2(n_841),
.B1(n_743),
.B2(n_599),
.C(n_1041),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1080),
.A2(n_1082),
.B(n_977),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1123),
.A2(n_1135),
.B(n_1157),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1210),
.Y(n_1343)
);

NOR2x1_ASAP7_75t_SL g1344 ( 
.A(n_1227),
.B(n_951),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1080),
.A2(n_1082),
.B(n_977),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1080),
.A2(n_1082),
.B(n_977),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1131),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1131),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1092),
.B(n_902),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1098),
.A2(n_1107),
.A3(n_1137),
.B(n_1189),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1123),
.A2(n_1135),
.B(n_1157),
.Y(n_1351)
);

O2A1O1Ixp5_ASAP7_75t_L g1352 ( 
.A1(n_1082),
.A2(n_1038),
.B(n_968),
.C(n_906),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1146),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1082),
.A2(n_821),
.B(n_789),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1098),
.A2(n_1107),
.A3(n_1137),
.B(n_1189),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1210),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1197),
.B(n_1215),
.Y(n_1357)
);

AOI221xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1082),
.A2(n_906),
.B1(n_743),
.B2(n_1224),
.C(n_1071),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1098),
.A2(n_1107),
.A3(n_1137),
.B(n_1189),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1146),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1082),
.A2(n_1042),
.B1(n_903),
.B2(n_1043),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_SL g1362 ( 
.A(n_1082),
.B(n_1043),
.C(n_756),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1123),
.A2(n_1135),
.B(n_1157),
.Y(n_1363)
);

O2A1O1Ixp5_ASAP7_75t_L g1364 ( 
.A1(n_1082),
.A2(n_1038),
.B(n_968),
.C(n_906),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1081),
.B(n_903),
.Y(n_1365)
);

AOI221x1_ASAP7_75t_L g1366 ( 
.A1(n_1082),
.A2(n_1038),
.B1(n_1207),
.B2(n_968),
.C(n_1098),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1081),
.B(n_903),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1107),
.A2(n_1189),
.B(n_1098),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1106),
.B(n_769),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1096),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1080),
.A2(n_1082),
.B(n_977),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1107),
.A2(n_1189),
.B(n_1098),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1131),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1082),
.A2(n_1042),
.B1(n_903),
.B2(n_1043),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1096),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1082),
.B(n_594),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1277),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1349),
.B(n_1319),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1352),
.B(n_1364),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1289),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1320),
.B(n_1249),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1249),
.B(n_1254),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1274),
.A2(n_1292),
.B(n_1287),
.C(n_1361),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1263),
.B(n_1369),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1333),
.B(n_1357),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1299),
.A2(n_1301),
.B(n_1247),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1274),
.A2(n_1292),
.B(n_1287),
.C(n_1374),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1264),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1366),
.A2(n_1267),
.B(n_1362),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1245),
.A2(n_1325),
.B(n_1304),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1243),
.A2(n_1271),
.B(n_1256),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1257),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1295),
.A2(n_1288),
.B1(n_1374),
.B2(n_1361),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1239),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1340),
.A2(n_1293),
.B1(n_1376),
.B2(n_1286),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1299),
.A2(n_1324),
.B(n_1323),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1358),
.A2(n_1339),
.B(n_1365),
.C(n_1367),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1294),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1303),
.B(n_1339),
.Y(n_1399)
);

AOI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1246),
.A2(n_1233),
.B(n_1231),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1324),
.A2(n_1228),
.B(n_1346),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1253),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1303),
.B(n_1365),
.Y(n_1403)
);

AND2x4_ASAP7_75t_SL g1404 ( 
.A(n_1258),
.B(n_1338),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1370),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1235),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1315),
.Y(n_1407)
);

AO21x2_ASAP7_75t_L g1408 ( 
.A1(n_1341),
.A2(n_1345),
.B(n_1371),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1367),
.B(n_1319),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1332),
.B(n_1354),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1344),
.A2(n_1260),
.B(n_1291),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1273),
.A2(n_1276),
.B(n_1312),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1252),
.B(n_1242),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1272),
.B(n_1229),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1329),
.B(n_1340),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1270),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1358),
.A2(n_1251),
.B(n_1284),
.C(n_1250),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1315),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1253),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1314),
.B(n_1302),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1244),
.B(n_1265),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1268),
.A2(n_1281),
.B(n_1251),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1375),
.B(n_1291),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1313),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1335),
.A2(n_1290),
.B(n_1240),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1326),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1316),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1241),
.A2(n_1368),
.B(n_1372),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1317),
.Y(n_1429)
);

NAND2xp33_ASAP7_75t_SL g1430 ( 
.A(n_1279),
.B(n_1282),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1296),
.A2(n_1322),
.B1(n_1311),
.B2(n_1295),
.Y(n_1431)
);

AO32x2_ASAP7_75t_L g1432 ( 
.A1(n_1322),
.A2(n_1283),
.A3(n_1350),
.B1(n_1355),
.B2(n_1359),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1357),
.B(n_1321),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1311),
.A2(n_1310),
.B1(n_1337),
.B2(n_1245),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1261),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1255),
.A2(n_1234),
.B(n_1306),
.Y(n_1436)
);

INVx6_ASAP7_75t_L g1437 ( 
.A(n_1257),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1308),
.A2(n_1241),
.B(n_1305),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1350),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1237),
.A2(n_1275),
.B1(n_1334),
.B2(n_1328),
.Y(n_1440)
);

AOI22x1_ASAP7_75t_L g1441 ( 
.A1(n_1331),
.A2(n_1336),
.B1(n_1356),
.B2(n_1248),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1360),
.B(n_1353),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1236),
.B(n_1259),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1280),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1350),
.Y(n_1445)
);

CKINVDCx6p67_ASAP7_75t_R g1446 ( 
.A(n_1232),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1320),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1343),
.A2(n_1356),
.B(n_1262),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1330),
.B(n_1327),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1269),
.B(n_1318),
.Y(n_1450)
);

INVxp67_ASAP7_75t_SL g1451 ( 
.A(n_1343),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1355),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1262),
.A2(n_1285),
.B(n_1300),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1230),
.Y(n_1454)
);

AOI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1355),
.A2(n_1359),
.B(n_1278),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1230),
.A2(n_1297),
.B1(n_1300),
.B2(n_1285),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1266),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1307),
.A2(n_1266),
.B(n_1298),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1307),
.A2(n_1298),
.B(n_1309),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1309),
.A2(n_1347),
.B(n_1348),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1309),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1347),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1347),
.A2(n_1348),
.B(n_1373),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1348),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1373),
.A2(n_1351),
.B(n_1342),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1373),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1239),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1277),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1332),
.B(n_1227),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1340),
.A2(n_1274),
.B1(n_1362),
.B2(n_1042),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1366),
.A2(n_1247),
.A3(n_1107),
.B(n_1082),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1352),
.B(n_1082),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1253),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1249),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1349),
.B(n_902),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1277),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1274),
.A2(n_775),
.B1(n_756),
.B2(n_743),
.C(n_599),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1340),
.A2(n_1040),
.B1(n_1043),
.B2(n_649),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1342),
.A2(n_1363),
.B(n_1351),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1349),
.B(n_902),
.Y(n_1480)
);

XOR2xp5_ASAP7_75t_L g1481 ( 
.A(n_1297),
.B(n_506),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1362),
.A2(n_1082),
.B(n_906),
.C(n_756),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1277),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1315),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1249),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1277),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1320),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1342),
.A2(n_1363),
.B(n_1351),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1239),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1299),
.A2(n_1301),
.B(n_1238),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1249),
.B(n_1254),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1249),
.B(n_1254),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_SL g1493 ( 
.A1(n_1344),
.A2(n_1292),
.B(n_1287),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1277),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1342),
.A2(n_1363),
.B(n_1351),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1274),
.A2(n_775),
.B1(n_756),
.B2(n_743),
.C(n_599),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1264),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1362),
.B(n_1082),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1315),
.Y(n_1499)
);

NAND2x1p5_ASAP7_75t_L g1500 ( 
.A(n_1320),
.B(n_1192),
.Y(n_1500)
);

BUFx2_ASAP7_75t_SL g1501 ( 
.A(n_1353),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1362),
.B(n_1082),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1362),
.B(n_1082),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1257),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1277),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1277),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1249),
.B(n_1254),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1299),
.A2(n_1301),
.B(n_1238),
.Y(n_1508)
);

AO21x1_ASAP7_75t_L g1509 ( 
.A1(n_1292),
.A2(n_1374),
.B(n_1361),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1247),
.A2(n_1082),
.B(n_1341),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1349),
.B(n_902),
.Y(n_1511)
);

AO21x2_ASAP7_75t_L g1512 ( 
.A1(n_1299),
.A2(n_1247),
.B(n_1324),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1320),
.B(n_1192),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1342),
.A2(n_1363),
.B(n_1351),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1299),
.A2(n_1301),
.B(n_1238),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1253),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1349),
.B(n_902),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1369),
.B(n_769),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1315),
.Y(n_1519)
);

O2A1O1Ixp5_ASAP7_75t_L g1520 ( 
.A1(n_1509),
.A2(n_1472),
.B(n_1387),
.C(n_1383),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1477),
.B(n_1496),
.Y(n_1521)
);

CKINVDCx11_ASAP7_75t_R g1522 ( 
.A(n_1388),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1447),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1420),
.B(n_1413),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1385),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1482),
.A2(n_1387),
.B(n_1383),
.C(n_1498),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1510),
.A2(n_1472),
.B(n_1512),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1399),
.A2(n_1403),
.B1(n_1503),
.B2(n_1498),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_R g1529 ( 
.A(n_1416),
.B(n_1398),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1502),
.A2(n_1503),
.B(n_1390),
.C(n_1403),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1478),
.A2(n_1431),
.B1(n_1395),
.B2(n_1470),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1384),
.B(n_1415),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1475),
.B(n_1480),
.Y(n_1533)
);

O2A1O1Ixp5_ASAP7_75t_L g1534 ( 
.A1(n_1379),
.A2(n_1502),
.B(n_1393),
.C(n_1389),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1511),
.B(n_1517),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1378),
.B(n_1423),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1512),
.A2(n_1408),
.B(n_1379),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1399),
.A2(n_1431),
.B(n_1395),
.C(n_1450),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1408),
.A2(n_1417),
.B(n_1422),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1406),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1470),
.A2(n_1393),
.B1(n_1434),
.B2(n_1518),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1397),
.A2(n_1450),
.B(n_1419),
.Y(n_1542)
);

AOI21x1_ASAP7_75t_SL g1543 ( 
.A1(n_1439),
.A2(n_1418),
.B(n_1407),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1409),
.B(n_1435),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1434),
.A2(n_1421),
.B1(n_1414),
.B2(n_1456),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1407),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1398),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1447),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1409),
.B(n_1426),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1397),
.A2(n_1402),
.B(n_1516),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1436),
.A2(n_1449),
.B(n_1386),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1421),
.A2(n_1414),
.B1(n_1456),
.B2(n_1469),
.Y(n_1552)
);

AOI21x1_ASAP7_75t_SL g1553 ( 
.A1(n_1484),
.A2(n_1519),
.B(n_1499),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1430),
.A2(n_1440),
.B(n_1474),
.C(n_1485),
.Y(n_1554)
);

OA21x2_ASAP7_75t_L g1555 ( 
.A1(n_1425),
.A2(n_1428),
.B(n_1438),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1473),
.A2(n_1449),
.B(n_1469),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_SL g1557 ( 
.A(n_1410),
.B(n_1449),
.Y(n_1557)
);

AND2x6_ASAP7_75t_L g1558 ( 
.A(n_1429),
.B(n_1474),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1484),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1469),
.A2(n_1500),
.B(n_1513),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_1388),
.Y(n_1561)
);

AND2x2_ASAP7_75t_SL g1562 ( 
.A(n_1396),
.B(n_1386),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1493),
.A2(n_1411),
.B(n_1500),
.C(n_1513),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1447),
.A2(n_1487),
.B(n_1416),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1442),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1424),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1487),
.A2(n_1443),
.B(n_1410),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1394),
.Y(n_1568)
);

CKINVDCx16_ASAP7_75t_R g1569 ( 
.A(n_1497),
.Y(n_1569)
);

AOI21x1_ASAP7_75t_SL g1570 ( 
.A1(n_1499),
.A2(n_1519),
.B(n_1385),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1382),
.B(n_1491),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1429),
.B(n_1380),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1405),
.B(n_1468),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1394),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1492),
.B(n_1507),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1485),
.B(n_1385),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1441),
.A2(n_1410),
.B1(n_1444),
.B2(n_1467),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1467),
.Y(n_1578)
);

NOR2xp67_ASAP7_75t_L g1579 ( 
.A(n_1427),
.B(n_1454),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1381),
.A2(n_1489),
.B1(n_1501),
.B2(n_1404),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1433),
.B(n_1468),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1483),
.B(n_1486),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1433),
.B(n_1483),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1486),
.B(n_1506),
.Y(n_1584)
);

O2A1O1Ixp5_ASAP7_75t_L g1585 ( 
.A1(n_1455),
.A2(n_1400),
.B(n_1445),
.C(n_1452),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1479),
.A2(n_1495),
.B(n_1488),
.Y(n_1586)
);

AOI21x1_ASAP7_75t_SL g1587 ( 
.A1(n_1433),
.A2(n_1471),
.B(n_1432),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1381),
.A2(n_1404),
.B1(n_1481),
.B2(n_1504),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1377),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_R g1590 ( 
.A(n_1457),
.B(n_1497),
.Y(n_1590)
);

AOI21x1_ASAP7_75t_SL g1591 ( 
.A1(n_1471),
.A2(n_1432),
.B(n_1401),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1476),
.A2(n_1505),
.B(n_1494),
.C(n_1463),
.Y(n_1592)
);

AOI21x1_ASAP7_75t_SL g1593 ( 
.A1(n_1471),
.A2(n_1432),
.B(n_1401),
.Y(n_1593)
);

AND2x2_ASAP7_75t_SL g1594 ( 
.A(n_1396),
.B(n_1401),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1471),
.Y(n_1595)
);

AOI21x1_ASAP7_75t_SL g1596 ( 
.A1(n_1432),
.A2(n_1396),
.B(n_1459),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1451),
.Y(n_1597)
);

A2O1A1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1487),
.A2(n_1464),
.B(n_1466),
.C(n_1458),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1448),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1465),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1453),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1392),
.A2(n_1504),
.B1(n_1437),
.B2(n_1457),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1392),
.A2(n_1504),
.B1(n_1437),
.B2(n_1443),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1443),
.A2(n_1462),
.B(n_1461),
.C(n_1515),
.Y(n_1604)
);

O2A1O1Ixp5_ASAP7_75t_L g1605 ( 
.A1(n_1490),
.A2(n_1508),
.B(n_1412),
.C(n_1391),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1446),
.B(n_1460),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1508),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1392),
.B(n_1437),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1514),
.B(n_1384),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1478),
.A2(n_1043),
.B1(n_1040),
.B2(n_1082),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1378),
.B(n_1423),
.Y(n_1611)
);

CKINVDCx11_ASAP7_75t_R g1612 ( 
.A(n_1388),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1384),
.B(n_1415),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1478),
.A2(n_1043),
.B1(n_1040),
.B2(n_1082),
.Y(n_1614)
);

O2A1O1Ixp5_ASAP7_75t_L g1615 ( 
.A1(n_1509),
.A2(n_1082),
.B(n_1364),
.C(n_1352),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1382),
.B(n_1491),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1407),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1378),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1384),
.B(n_1415),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1420),
.B(n_1413),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1384),
.B(n_1415),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1384),
.B(n_1415),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1384),
.B(n_1415),
.Y(n_1623)
);

NOR2xp67_ASAP7_75t_L g1624 ( 
.A(n_1402),
.B(n_1419),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1420),
.B(n_1413),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1407),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1478),
.A2(n_1043),
.B1(n_1040),
.B2(n_1082),
.Y(n_1627)
);

CKINVDCx16_ASAP7_75t_R g1628 ( 
.A(n_1388),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1384),
.B(n_1415),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1510),
.A2(n_1082),
.B(n_1247),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1420),
.B(n_1413),
.Y(n_1631)
);

NAND4xp25_ASAP7_75t_L g1632 ( 
.A(n_1477),
.B(n_1496),
.C(n_868),
.D(n_775),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1609),
.B(n_1601),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1607),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1586),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1605),
.A2(n_1585),
.B(n_1551),
.Y(n_1636)
);

AO21x2_ASAP7_75t_L g1637 ( 
.A1(n_1539),
.A2(n_1537),
.B(n_1527),
.Y(n_1637)
);

BUFx4f_ASAP7_75t_L g1638 ( 
.A(n_1558),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1528),
.B(n_1530),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1528),
.B(n_1544),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1546),
.B(n_1559),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1526),
.A2(n_1615),
.B(n_1534),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1521),
.A2(n_1632),
.B1(n_1531),
.B2(n_1545),
.Y(n_1643)
);

BUFx5_ASAP7_75t_L g1644 ( 
.A(n_1562),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1532),
.B(n_1613),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1619),
.B(n_1621),
.Y(n_1646)
);

AO21x1_ASAP7_75t_L g1647 ( 
.A1(n_1541),
.A2(n_1630),
.B(n_1614),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1559),
.B(n_1626),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1599),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1549),
.B(n_1524),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1617),
.Y(n_1651)
);

BUFx2_ASAP7_75t_SL g1652 ( 
.A(n_1579),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1540),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1623),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1555),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1595),
.B(n_1617),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1629),
.B(n_1566),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1597),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1538),
.A2(n_1627),
.B1(n_1610),
.B2(n_1625),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1589),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1594),
.Y(n_1661)
);

BUFx2_ASAP7_75t_SL g1662 ( 
.A(n_1578),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1594),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1600),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1596),
.A2(n_1591),
.B(n_1593),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1562),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1558),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_SL g1668 ( 
.A(n_1602),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1536),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1611),
.B(n_1618),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1581),
.B(n_1583),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1573),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1620),
.B(n_1631),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1582),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1558),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1553),
.A2(n_1543),
.B(n_1570),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1584),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1572),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1557),
.B(n_1525),
.Y(n_1679)
);

AO22x1_ASAP7_75t_L g1680 ( 
.A1(n_1642),
.A2(n_1552),
.B1(n_1603),
.B2(n_1577),
.Y(n_1680)
);

NOR2x1_ASAP7_75t_L g1681 ( 
.A(n_1642),
.B(n_1604),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1634),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1661),
.B(n_1520),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1664),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1643),
.A2(n_1588),
.B1(n_1554),
.B2(n_1533),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1661),
.B(n_1534),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1641),
.B(n_1565),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1653),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1651),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1635),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1535),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1666),
.B(n_1587),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1633),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1633),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1641),
.B(n_1568),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1647),
.A2(n_1571),
.B1(n_1575),
.B2(n_1616),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1678),
.B(n_1542),
.Y(n_1697)
);

OAI33xp33_ASAP7_75t_L g1698 ( 
.A1(n_1659),
.A2(n_1639),
.A3(n_1640),
.B1(n_1673),
.B2(n_1650),
.B3(n_1660),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1670),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1660),
.B(n_1574),
.Y(n_1700)
);

INVx6_ASAP7_75t_L g1701 ( 
.A(n_1679),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1639),
.A2(n_1659),
.B1(n_1647),
.B2(n_1640),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1669),
.B(n_1592),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1637),
.A2(n_1556),
.B(n_1567),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1668),
.A2(n_1569),
.B1(n_1628),
.B2(n_1560),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1644),
.B(n_1665),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1672),
.B(n_1598),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1671),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1648),
.B(n_1606),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1694),
.B(n_1644),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1682),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1690),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1702),
.B(n_1673),
.C(n_1650),
.Y(n_1713)
);

NAND2xp33_ASAP7_75t_R g1714 ( 
.A(n_1703),
.B(n_1529),
.Y(n_1714)
);

INVxp67_ASAP7_75t_SL g1715 ( 
.A(n_1707),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1682),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1695),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1702),
.A2(n_1654),
.B1(n_1645),
.B2(n_1646),
.C(n_1657),
.Y(n_1718)
);

AOI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1680),
.A2(n_1550),
.B(n_1580),
.C(n_1563),
.Y(n_1719)
);

OAI211xp5_ASAP7_75t_L g1720 ( 
.A1(n_1681),
.A2(n_1590),
.B(n_1658),
.C(n_1670),
.Y(n_1720)
);

NAND2xp33_ASAP7_75t_R g1721 ( 
.A(n_1703),
.B(n_1529),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1684),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1684),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1693),
.B(n_1644),
.Y(n_1724)
);

NAND4xp25_ASAP7_75t_L g1725 ( 
.A(n_1681),
.B(n_1624),
.C(n_1657),
.D(n_1654),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1698),
.A2(n_1645),
.B1(n_1646),
.B2(n_1677),
.C(n_1674),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1695),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_L g1728 ( 
.A(n_1705),
.B(n_1590),
.Y(n_1728)
);

NAND3xp33_ASAP7_75t_L g1729 ( 
.A(n_1697),
.B(n_1680),
.C(n_1685),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1693),
.B(n_1644),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1698),
.A2(n_1679),
.B1(n_1571),
.B2(n_1644),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1685),
.A2(n_1668),
.B1(n_1576),
.B2(n_1652),
.Y(n_1732)
);

OAI31xp33_ASAP7_75t_L g1733 ( 
.A1(n_1705),
.A2(n_1679),
.A3(n_1675),
.B(n_1667),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

OAI31xp33_ASAP7_75t_SL g1735 ( 
.A1(n_1686),
.A2(n_1679),
.A3(n_1608),
.B(n_1676),
.Y(n_1735)
);

AO21x1_ASAP7_75t_SL g1736 ( 
.A1(n_1697),
.A2(n_1648),
.B(n_1656),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1688),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1696),
.A2(n_1652),
.B1(n_1576),
.B2(n_1638),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1700),
.Y(n_1739)
);

OAI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1704),
.A2(n_1699),
.B1(n_1707),
.B2(n_1700),
.C(n_1687),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1699),
.A2(n_1638),
.B1(n_1637),
.B2(n_1662),
.Y(n_1741)
);

NAND4xp25_ASAP7_75t_SL g1742 ( 
.A(n_1686),
.B(n_1564),
.C(n_1561),
.D(n_1522),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_SL g1743 ( 
.A(n_1708),
.B(n_1547),
.C(n_1675),
.Y(n_1743)
);

AOI31xp33_ASAP7_75t_SL g1744 ( 
.A1(n_1709),
.A2(n_1656),
.A3(n_1649),
.B(n_1655),
.Y(n_1744)
);

OR2x6_ASAP7_75t_L g1745 ( 
.A(n_1701),
.B(n_1667),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1689),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1734),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1734),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1737),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_SL g1751 ( 
.A(n_1729),
.B(n_1686),
.C(n_1687),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1723),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1723),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1722),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1712),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1737),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1745),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1715),
.B(n_1683),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1711),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1711),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1716),
.Y(n_1761)
);

INVx4_ASAP7_75t_L g1762 ( 
.A(n_1745),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1745),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1720),
.B(n_1638),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1717),
.B(n_1683),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1745),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1745),
.B(n_1706),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1741),
.A2(n_1636),
.B(n_1665),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1724),
.B(n_1692),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1724),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1750),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1759),
.Y(n_1772)
);

NAND2x1p5_ASAP7_75t_L g1773 ( 
.A(n_1764),
.B(n_1741),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1753),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1757),
.B(n_1736),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1759),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1751),
.B(n_1612),
.Y(n_1777)
);

NOR2x1_ASAP7_75t_L g1778 ( 
.A(n_1751),
.B(n_1725),
.Y(n_1778)
);

CKINVDCx16_ASAP7_75t_R g1779 ( 
.A(n_1762),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1762),
.B(n_1730),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1757),
.B(n_1763),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1757),
.B(n_1736),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1758),
.B(n_1726),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1762),
.B(n_1730),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1758),
.B(n_1739),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1763),
.B(n_1735),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1762),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1750),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1754),
.B(n_1739),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1763),
.B(n_1710),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1766),
.B(n_1762),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1766),
.B(n_1710),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1761),
.Y(n_1793)
);

INVx4_ASAP7_75t_L g1794 ( 
.A(n_1766),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1761),
.Y(n_1795)
);

XOR2xp5_ASAP7_75t_L g1796 ( 
.A(n_1764),
.B(n_1742),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1747),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1753),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1754),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1747),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1765),
.B(n_1713),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1767),
.A2(n_1728),
.B1(n_1743),
.B2(n_1740),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1748),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1748),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1765),
.B(n_1727),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1752),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1769),
.B(n_1746),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1749),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1752),
.B(n_1718),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1749),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1756),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1767),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1756),
.B(n_1691),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_SL g1814 ( 
.A(n_1767),
.B(n_1733),
.Y(n_1814)
);

AND2x4_ASAP7_75t_SL g1815 ( 
.A(n_1767),
.B(n_1732),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1797),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1778),
.A2(n_1719),
.B1(n_1714),
.B2(n_1721),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1778),
.A2(n_1732),
.B1(n_1637),
.B2(n_1768),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1799),
.B(n_1687),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1797),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1779),
.B(n_1767),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1800),
.Y(n_1822)
);

AOI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1796),
.A2(n_1719),
.B1(n_1738),
.B2(n_1731),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1800),
.Y(n_1824)
);

INVx2_ASAP7_75t_SL g1825 ( 
.A(n_1774),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1796),
.A2(n_1802),
.B1(n_1777),
.B2(n_1773),
.Y(n_1826)
);

INVx5_ASAP7_75t_L g1827 ( 
.A(n_1794),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1773),
.A2(n_1768),
.B1(n_1637),
.B2(n_1683),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1803),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1803),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1804),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1799),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1806),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1804),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1809),
.B(n_1709),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1781),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1808),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1794),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1779),
.B(n_1770),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1808),
.Y(n_1840)
);

INVxp67_ASAP7_75t_SL g1841 ( 
.A(n_1798),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1810),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1815),
.B(n_1770),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1810),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1783),
.B(n_1691),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1811),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1772),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1772),
.Y(n_1848)
);

INVx2_ASAP7_75t_SL g1849 ( 
.A(n_1807),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1776),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1776),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1801),
.B(n_1709),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1833),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1846),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1846),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1828),
.B(n_1786),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1828),
.B(n_1786),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1832),
.B(n_1805),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1827),
.Y(n_1859)
);

INVx1_ASAP7_75t_SL g1860 ( 
.A(n_1827),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1827),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1816),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1820),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1821),
.B(n_1775),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1832),
.B(n_1805),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1822),
.Y(n_1866)
);

BUFx3_ASAP7_75t_L g1867 ( 
.A(n_1827),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1826),
.A2(n_1773),
.B1(n_1814),
.B2(n_1815),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1849),
.Y(n_1869)
);

INVx1_ASAP7_75t_SL g1870 ( 
.A(n_1825),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1849),
.Y(n_1871)
);

AO21x2_ASAP7_75t_L g1872 ( 
.A1(n_1841),
.A2(n_1795),
.B(n_1793),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1843),
.B(n_1781),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1825),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1838),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1841),
.B(n_1793),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1817),
.A2(n_1823),
.B1(n_1818),
.B2(n_1836),
.Y(n_1877)
);

INVx3_ASAP7_75t_SL g1878 ( 
.A(n_1838),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1839),
.B(n_1775),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1824),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1868),
.A2(n_1818),
.B1(n_1836),
.B2(n_1789),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1853),
.B(n_1814),
.Y(n_1882)
);

NOR3xp33_ASAP7_75t_L g1883 ( 
.A(n_1877),
.B(n_1848),
.C(n_1847),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1877),
.A2(n_1815),
.B1(n_1782),
.B2(n_1791),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1854),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1858),
.B(n_1845),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1854),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1867),
.Y(n_1888)
);

AOI221xp5_ASAP7_75t_L g1889 ( 
.A1(n_1853),
.A2(n_1851),
.B1(n_1850),
.B2(n_1794),
.C(n_1844),
.Y(n_1889)
);

OAI211xp5_ASAP7_75t_L g1890 ( 
.A1(n_1856),
.A2(n_1794),
.B(n_1787),
.C(n_1791),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1856),
.A2(n_1857),
.B(n_1876),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1855),
.Y(n_1892)
);

AND2x4_ASAP7_75t_SL g1893 ( 
.A(n_1873),
.B(n_1782),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1874),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1864),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1855),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1856),
.A2(n_1857),
.B1(n_1870),
.B2(n_1874),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1872),
.Y(n_1898)
);

OAI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1857),
.A2(n_1819),
.B1(n_1812),
.B2(n_1835),
.Y(n_1899)
);

AOI222xp33_ASAP7_75t_L g1900 ( 
.A1(n_1870),
.A2(n_1876),
.B1(n_1860),
.B2(n_1859),
.C1(n_1864),
.C2(n_1880),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1872),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1894),
.B(n_1891),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1893),
.B(n_1864),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1882),
.A2(n_1879),
.B1(n_1873),
.B2(n_1787),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1900),
.B(n_1895),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1897),
.B(n_1879),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1897),
.B(n_1858),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1888),
.Y(n_1908)
);

INVx1_ASAP7_75t_SL g1909 ( 
.A(n_1886),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1883),
.A2(n_1879),
.B1(n_1860),
.B2(n_1859),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1884),
.B(n_1865),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1889),
.B(n_1869),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1881),
.B(n_1865),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1885),
.B(n_1869),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1887),
.B(n_1869),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1902),
.A2(n_1881),
.B(n_1898),
.Y(n_1916)
);

AOI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1913),
.A2(n_1907),
.B(n_1905),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1906),
.A2(n_1901),
.B(n_1899),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1911),
.A2(n_1890),
.B1(n_1892),
.B2(n_1896),
.C(n_1880),
.Y(n_1919)
);

AOI21xp33_ASAP7_75t_SL g1920 ( 
.A1(n_1910),
.A2(n_1878),
.B(n_1871),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1914),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1914),
.Y(n_1922)
);

NOR3xp33_ASAP7_75t_L g1923 ( 
.A(n_1912),
.B(n_1861),
.C(n_1867),
.Y(n_1923)
);

O2A1O1Ixp33_ASAP7_75t_L g1924 ( 
.A1(n_1915),
.A2(n_1909),
.B(n_1908),
.C(n_1867),
.Y(n_1924)
);

AOI21xp33_ASAP7_75t_SL g1925 ( 
.A1(n_1903),
.A2(n_1878),
.B(n_1871),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1904),
.B(n_1871),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_SL g1927 ( 
.A(n_1913),
.B(n_1861),
.C(n_1875),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1917),
.A2(n_1872),
.B1(n_1787),
.B2(n_1861),
.Y(n_1928)
);

A2O1A1Ixp33_ASAP7_75t_L g1929 ( 
.A1(n_1916),
.A2(n_1862),
.B(n_1866),
.C(n_1863),
.Y(n_1929)
);

NAND4xp25_ASAP7_75t_L g1930 ( 
.A(n_1919),
.B(n_1875),
.C(n_1866),
.D(n_1863),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_SL g1931 ( 
.A1(n_1918),
.A2(n_1787),
.B(n_1862),
.Y(n_1931)
);

A2O1A1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1920),
.A2(n_1875),
.B(n_1830),
.C(n_1829),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1925),
.B(n_1878),
.Y(n_1933)
);

AOI221xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1924),
.A2(n_1837),
.B1(n_1831),
.B2(n_1842),
.C(n_1840),
.Y(n_1934)
);

XNOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1931),
.B(n_1921),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1933),
.B(n_1923),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1929),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1934),
.Y(n_1938)
);

INVxp67_ASAP7_75t_L g1939 ( 
.A(n_1930),
.Y(n_1939)
);

XNOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1928),
.B(n_1922),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1932),
.Y(n_1941)
);

O2A1O1Ixp33_ASAP7_75t_L g1942 ( 
.A1(n_1937),
.A2(n_1927),
.B(n_1926),
.C(n_1872),
.Y(n_1942)
);

AOI211xp5_ASAP7_75t_L g1943 ( 
.A1(n_1936),
.A2(n_1834),
.B(n_1780),
.C(n_1784),
.Y(n_1943)
);

OA22x2_ASAP7_75t_L g1944 ( 
.A1(n_1939),
.A2(n_1795),
.B1(n_1812),
.B2(n_1811),
.Y(n_1944)
);

INVx4_ASAP7_75t_SL g1945 ( 
.A(n_1941),
.Y(n_1945)
);

AO221x1_ASAP7_75t_L g1946 ( 
.A1(n_1939),
.A2(n_1812),
.B1(n_1788),
.B2(n_1771),
.C(n_1548),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1935),
.Y(n_1947)
);

AOI211xp5_ASAP7_75t_L g1948 ( 
.A1(n_1942),
.A2(n_1947),
.B(n_1938),
.C(n_1943),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1945),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1944),
.A2(n_1940),
.B(n_1785),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1949),
.Y(n_1951)
);

NAND3xp33_ASAP7_75t_L g1952 ( 
.A(n_1951),
.B(n_1948),
.C(n_1950),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1952),
.B(n_1780),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1952),
.Y(n_1954)
);

AOI22x1_ASAP7_75t_L g1955 ( 
.A1(n_1954),
.A2(n_1946),
.B1(n_1771),
.B2(n_1788),
.Y(n_1955)
);

AOI21xp33_ASAP7_75t_L g1956 ( 
.A1(n_1953),
.A2(n_1852),
.B(n_1784),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_SL g1957 ( 
.A1(n_1955),
.A2(n_1812),
.B1(n_1662),
.B2(n_1780),
.Y(n_1957)
);

AOI22x1_ASAP7_75t_L g1958 ( 
.A1(n_1956),
.A2(n_1771),
.B1(n_1788),
.B2(n_1780),
.Y(n_1958)
);

XNOR2xp5_ASAP7_75t_L g1959 ( 
.A(n_1958),
.B(n_1784),
.Y(n_1959)
);

AO221x2_ASAP7_75t_L g1960 ( 
.A1(n_1959),
.A2(n_1957),
.B1(n_1813),
.B2(n_1750),
.C(n_1755),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1960),
.A2(n_1784),
.B(n_1790),
.Y(n_1961)
);

NAND3xp33_ASAP7_75t_L g1962 ( 
.A(n_1961),
.B(n_1792),
.C(n_1790),
.Y(n_1962)
);

AOI221xp5_ASAP7_75t_L g1963 ( 
.A1(n_1962),
.A2(n_1792),
.B1(n_1807),
.B2(n_1770),
.C(n_1760),
.Y(n_1963)
);

AOI211xp5_ASAP7_75t_L g1964 ( 
.A1(n_1963),
.A2(n_1523),
.B(n_1548),
.C(n_1744),
.Y(n_1964)
);


endmodule