module fake_jpeg_15659_n_215 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_18),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_26),
.B1(n_30),
.B2(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_23),
.B1(n_29),
.B2(n_28),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_24),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx2_ASAP7_75t_SL g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_57),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_23),
.B1(n_29),
.B2(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_35),
.B1(n_16),
.B2(n_24),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_52),
.B1(n_44),
.B2(n_53),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_39),
.B1(n_21),
.B2(n_20),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_77),
.Y(n_86)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_73),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_74),
.B1(n_66),
.B2(n_75),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_16),
.B(n_26),
.C(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_27),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_34),
.C(n_33),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_33),
.C(n_34),
.Y(n_94)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_44),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_55),
.C(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_99),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_42),
.B(n_58),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_71),
.B(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_92),
.B1(n_98),
.B2(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_42),
.B1(n_39),
.B2(n_47),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_54),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_96),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_80),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_34),
.C(n_33),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_64),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_25),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_72),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_34),
.B1(n_19),
.B2(n_2),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_72),
.B1(n_73),
.B2(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_113),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_76),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_117),
.B(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_115),
.Y(n_126)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_81),
.B(n_62),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_125),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_30),
.B(n_22),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_87),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_64),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_133),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_103),
.B1(n_84),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_143),
.B1(n_82),
.B2(n_77),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_84),
.B(n_98),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_109),
.B(n_120),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_90),
.B(n_83),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_112),
.B(n_101),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_137),
.B(n_25),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_107),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_139),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

AOI22x1_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_94),
.B1(n_100),
.B2(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_150),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_123),
.C(n_114),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_153),
.C(n_161),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_118),
.B(n_105),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_152),
.B1(n_157),
.B2(n_126),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_105),
.B(n_115),
.C(n_124),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_154),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_136),
.B(n_143),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_101),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_124),
.B(n_82),
.C(n_25),
.D(n_30),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_132),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_106),
.C(n_113),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_134),
.C(n_129),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_166),
.C(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_144),
.C(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_156),
.A2(n_127),
.B1(n_138),
.B2(n_77),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_169),
.A2(n_160),
.B1(n_154),
.B2(n_146),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_138),
.C(n_131),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_169),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_145),
.B1(n_157),
.B2(n_152),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_175),
.A2(n_185),
.B1(n_166),
.B2(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_173),
.A2(n_148),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_150),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_151),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_162),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_89),
.B1(n_1),
.B2(n_3),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_176),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_190),
.C(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_165),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_4),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_176),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_0),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.C(n_201),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_178),
.A3(n_182),
.B1(n_180),
.B2(n_185),
.C1(n_181),
.C2(n_67),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_200),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_182),
.C(n_5),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_67),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_193),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_189),
.C(n_193),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_5),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_12),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_5),
.B(n_6),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_12),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_206),
.B(n_4),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_208),
.B(n_209),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_6),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_9),
.B(n_10),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

AOI211xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_11),
.B(n_205),
.C(n_188),
.Y(n_214)
);


endmodule