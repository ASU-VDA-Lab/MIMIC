module fake_jpeg_13144_n_388 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_388);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_388;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_50),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_60),
.Y(n_102)
);

INVx8_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_82),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_0),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_24),
.B(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_74),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_83),
.B(n_28),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_32),
.B1(n_17),
.B2(n_42),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_104),
.B1(n_108),
.B2(n_75),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_32),
.B1(n_38),
.B2(n_15),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_87),
.A2(n_103),
.B(n_8),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

OA22x2_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_38),
.B1(n_28),
.B2(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_45),
.A2(n_15),
.B1(n_26),
.B2(n_18),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_25),
.B1(n_12),
.B2(n_11),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_47),
.A2(n_14),
.B1(n_13),
.B2(n_18),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_1),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_43),
.A2(n_28),
.B1(n_26),
.B2(n_18),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_110),
.A2(n_115),
.B(n_127),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_46),
.A2(n_64),
.B1(n_58),
.B2(n_77),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_13),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_122),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_46),
.A2(n_16),
.B1(n_80),
.B2(n_63),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_72),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_70),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_0),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_132),
.B(n_1),
.Y(n_135)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_135),
.B(n_147),
.Y(n_186)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_136),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_53),
.B1(n_52),
.B2(n_44),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_137),
.A2(n_138),
.B1(n_144),
.B2(n_160),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_48),
.B1(n_62),
.B2(n_67),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx6_ASAP7_75t_SL g198 ( 
.A(n_140),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_141),
.B(n_142),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_105),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_84),
.B(n_73),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_150),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_50),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_95),
.A2(n_68),
.B1(n_51),
.B2(n_71),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_155),
.Y(n_211)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_96),
.A2(n_121),
.B1(n_99),
.B2(n_88),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_159),
.B1(n_168),
.B2(n_131),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_164),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_49),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_98),
.A2(n_57),
.B(n_78),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_156),
.A2(n_167),
.B(n_173),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_1),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_169),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_99),
.A2(n_57),
.B1(n_4),
.B2(n_5),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_110),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_165),
.B1(n_171),
.B2(n_160),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_2),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_101),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_90),
.B(n_7),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_123),
.B(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_9),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_112),
.A2(n_9),
.B1(n_101),
.B2(n_126),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_93),
.C(n_111),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g174 ( 
.A(n_89),
.Y(n_174)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_107),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_176),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_93),
.B(n_91),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_SL g177 ( 
.A(n_131),
.B(n_91),
.C(n_116),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_166),
.B(n_168),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_180),
.A2(n_140),
.B1(n_149),
.B2(n_172),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_116),
.B1(n_126),
.B2(n_111),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_181),
.A2(n_192),
.B1(n_214),
.B2(n_197),
.Y(n_250)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_107),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_184),
.B(n_201),
.Y(n_245)
);

CKINVDCx10_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_166),
.A2(n_94),
.B1(n_120),
.B2(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_120),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_196),
.Y(n_221)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_94),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_142),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_219),
.B(n_192),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_218),
.Y(n_237)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_202),
.B1(n_189),
.B2(n_193),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_173),
.B1(n_137),
.B2(n_152),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_175),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_178),
.B(n_157),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_167),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_146),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_227),
.C(n_197),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_207),
.A2(n_177),
.B1(n_146),
.B2(n_162),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_223),
.A2(n_236),
.B1(n_239),
.B2(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_136),
.C(n_175),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_167),
.B1(n_171),
.B2(n_165),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_228),
.A2(n_220),
.B(n_198),
.Y(n_273)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_194),
.B(n_133),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_233),
.B(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_186),
.B(n_143),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_161),
.B1(n_163),
.B2(n_179),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_151),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_243),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_203),
.A2(n_179),
.B1(n_161),
.B2(n_163),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_188),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g244 ( 
.A(n_186),
.B(n_157),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_251),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_248),
.A2(n_250),
.B1(n_217),
.B2(n_212),
.Y(n_284)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_201),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_198),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_220),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_211),
.B(n_196),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_237),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_209),
.B1(n_184),
.B2(n_191),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_267),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_263),
.C(n_265),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_260),
.B(n_229),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_222),
.C(n_237),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_221),
.C(n_210),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_266),
.B(n_278),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_228),
.A2(n_191),
.B1(n_214),
.B2(n_216),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_210),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_185),
.C(n_182),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_221),
.B(n_210),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_270),
.B(n_282),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g271 ( 
.A1(n_223),
.A2(n_218),
.A3(n_185),
.B1(n_215),
.B2(n_182),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_230),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_273),
.A2(n_284),
.B1(n_226),
.B2(n_241),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_252),
.B1(n_239),
.B2(n_238),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_234),
.B1(n_243),
.B2(n_242),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_220),
.B(n_190),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_277),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_225),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_280),
.B(n_274),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_253),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_230),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_224),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_277),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_285),
.B(n_305),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_279),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_288),
.Y(n_318)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_297),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_291),
.B(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_240),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_304),
.C(n_298),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_262),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_264),
.B1(n_258),
.B2(n_261),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_261),
.B1(n_258),
.B2(n_274),
.Y(n_309)
);

A2O1A1O1Ixp25_ASAP7_75t_L g303 ( 
.A1(n_276),
.A2(n_246),
.B(n_190),
.C(n_206),
.D(n_195),
.Y(n_303)
);

OA21x2_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_264),
.B(n_282),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_256),
.B(n_208),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_308),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_290),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_309),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_255),
.B1(n_267),
.B2(n_272),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_272),
.B1(n_271),
.B2(n_275),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_268),
.B1(n_273),
.B2(n_259),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_322),
.C(n_304),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_317),
.A2(n_300),
.B1(n_288),
.B2(n_328),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_291),
.C(n_299),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_265),
.C(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

FAx1_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_269),
.CI(n_232),
.CON(n_325),
.SN(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_328),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_294),
.A2(n_269),
.B1(n_247),
.B2(n_232),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_217),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_298),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_339),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_334),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_332),
.A2(n_313),
.B1(n_309),
.B2(n_327),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_333),
.A2(n_319),
.B(n_326),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_299),
.C(n_297),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_303),
.B(n_296),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_336),
.A2(n_324),
.B(n_310),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_301),
.C(n_293),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_340),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_287),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_289),
.C(n_307),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_307),
.C(n_204),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_345),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_323),
.B(n_204),
.Y(n_343)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_326),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_344),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_208),
.C(n_200),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_316),
.Y(n_346)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_342),
.B1(n_341),
.B2(n_345),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_318),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_325),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_355),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_335),
.A2(n_310),
.B1(n_321),
.B2(n_312),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_347),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_358),
.A2(n_329),
.B(n_340),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_330),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_366),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_362),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_363),
.B(n_364),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_346),
.A2(n_342),
.B1(n_325),
.B2(n_321),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_331),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_365),
.A2(n_350),
.B(n_356),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_SL g367 ( 
.A(n_351),
.B(n_312),
.Y(n_367)
);

AOI21xp33_ASAP7_75t_L g370 ( 
.A1(n_367),
.A2(n_325),
.B(n_351),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_356),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_373),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_370),
.B(n_374),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_354),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_350),
.C(n_373),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_377),
.C(n_379),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_375),
.A2(n_361),
.B(n_368),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_369),
.A2(n_364),
.B1(n_366),
.B2(n_349),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_371),
.Y(n_381)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_381),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_380),
.Y(n_383)
);

MAJx2_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_371),
.C(n_200),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_384),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_385),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_387),
.B(n_382),
.Y(n_388)
);


endmodule