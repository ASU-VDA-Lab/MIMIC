module fake_netlist_1_9710_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
OA21x2_ASAP7_75t_L g11 ( .A1(n_7), .A2(n_0), .B(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_6), .B(n_8), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_13), .B(n_1), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
NAND2x1p5_ASAP7_75t_L g19 ( .A(n_16), .B(n_1), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_13), .B(n_15), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_18), .A2(n_15), .B(n_14), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AND4x1_ASAP7_75t_L g26 ( .A(n_25), .B(n_17), .C(n_23), .D(n_20), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_24), .B(n_19), .Y(n_27) );
O2A1O1Ixp33_ASAP7_75t_SL g28 ( .A1(n_27), .A2(n_24), .B(n_21), .C(n_14), .Y(n_28) );
OAI22xp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_17), .B1(n_11), .B2(n_21), .Y(n_29) );
AOI221xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_16), .B1(n_12), .B2(n_21), .C(n_22), .Y(n_30) );
OAI22xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_16), .B1(n_12), .B2(n_11), .Y(n_31) );
AOI221xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_16), .B1(n_22), .B2(n_11), .C(n_5), .Y(n_32) );
NOR3xp33_ASAP7_75t_L g33 ( .A(n_32), .B(n_22), .C(n_11), .Y(n_33) );
NOR2x1_ASAP7_75t_L g34 ( .A(n_31), .B(n_11), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_30), .Y(n_35) );
OA22x2_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_11), .B1(n_3), .B2(n_4), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
O2A1O1Ixp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_33), .B(n_5), .C(n_6), .Y(n_38) );
OAI222xp33_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_2), .B1(n_9), .B2(n_10), .C1(n_36), .C2(n_37), .Y(n_39) );
endmodule