module fake_aes_5435_n_832 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_832);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_832;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_769;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_613;
wire n_490;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_698;
wire n_555;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_23), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_20), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_65), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_70), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_57), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_54), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_102), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_6), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_92), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_62), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_55), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_84), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_40), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_43), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_60), .Y(n_121) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_18), .B(n_1), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_37), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_6), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_75), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_103), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_34), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_18), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_11), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_8), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_58), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_44), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_100), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_14), .Y(n_135) );
INVxp67_ASAP7_75t_SL g136 ( .A(n_45), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_19), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_10), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_31), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_88), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_99), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_2), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_109), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_140), .B(n_0), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_109), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
CKINVDCx11_ASAP7_75t_R g150 ( .A(n_121), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_140), .B(n_1), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_110), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_116), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_110), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_106), .B(n_2), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_112), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_112), .B(n_24), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_119), .A2(n_49), .B(n_98), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_105), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_125), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_125), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_120), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_117), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_167), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_160), .A2(n_134), .B1(n_114), .B2(n_129), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_167), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_167), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_167), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_163), .B(n_115), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_163), .B(n_108), .Y(n_175) );
AO22x2_ASAP7_75t_L g176 ( .A1(n_160), .A2(n_120), .B1(n_144), .B2(n_143), .Y(n_176) );
NAND2xp33_ASAP7_75t_L g177 ( .A(n_146), .B(n_111), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_150), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_151), .B(n_128), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_151), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_146), .B(n_117), .Y(n_183) );
BUFx6f_ASAP7_75t_SL g184 ( .A(n_160), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_167), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_151), .B(n_106), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_147), .A2(n_107), .B1(n_135), .B2(n_137), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_147), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_154), .B(n_130), .Y(n_195) );
OAI22xp33_ASAP7_75t_L g196 ( .A1(n_155), .A2(n_145), .B1(n_107), .B2(n_135), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_149), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_154), .B(n_137), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_157), .B(n_138), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_149), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_149), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_161), .B(n_113), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_161), .B(n_118), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_172), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_181), .B(n_166), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
O2A1O1Ixp5_ASAP7_75t_L g209 ( .A1(n_205), .A2(n_166), .B(n_155), .C(n_136), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_172), .Y(n_210) );
INVxp67_ASAP7_75t_L g211 ( .A(n_179), .Y(n_211) );
NOR3xp33_ASAP7_75t_L g212 ( .A(n_169), .B(n_124), .C(n_145), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_181), .B(n_123), .Y(n_214) );
NAND2xp33_ASAP7_75t_L g215 ( .A(n_192), .B(n_131), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_186), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_176), .A2(n_165), .B1(n_164), .B2(n_143), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_174), .B(n_139), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_186), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_176), .A2(n_165), .B1(n_164), .B2(n_144), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_194), .B(n_122), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_175), .B(n_142), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_186), .B(n_126), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_186), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_187), .Y(n_225) );
NOR3xp33_ASAP7_75t_L g226 ( .A(n_169), .B(n_126), .C(n_127), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_187), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_201), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_201), .B(n_127), .Y(n_229) );
NOR2xp33_ASAP7_75t_R g230 ( .A(n_178), .B(n_133), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_189), .B(n_133), .Y(n_231) );
INVx4_ASAP7_75t_L g232 ( .A(n_184), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_184), .A2(n_132), .B1(n_141), .B2(n_165), .Y(n_234) );
AO221x1_ASAP7_75t_L g235 ( .A1(n_176), .A2(n_165), .B1(n_164), .B2(n_141), .C(n_132), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_194), .B(n_162), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_196), .B(n_192), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_188), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_189), .B(n_164), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_195), .B(n_164), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_184), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_170), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_176), .B(n_162), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_190), .B(n_3), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_193), .B(n_164), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_204), .B(n_164), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_200), .A2(n_153), .B(n_156), .C(n_158), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_200), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_198), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_198), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_183), .B(n_165), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_177), .B(n_165), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_184), .B(n_165), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_211), .B(n_176), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_228), .B(n_3), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_207), .B(n_162), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_212), .B(n_4), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_252), .A2(n_162), .B1(n_153), .B2(n_156), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_207), .B(n_162), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_229), .B(n_4), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_246), .A2(n_153), .B(n_156), .C(n_158), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_246), .A2(n_168), .B(n_180), .Y(n_264) );
AOI21x1_ASAP7_75t_L g265 ( .A1(n_244), .A2(n_168), .B(n_180), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_251), .B(n_5), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_251), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_231), .B(n_5), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_238), .B(n_7), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_245), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_226), .B(n_7), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_180), .B(n_170), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g274 ( .A(n_217), .B(n_220), .C(n_218), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_245), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_206), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_250), .A2(n_158), .B(n_159), .C(n_182), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_242), .A2(n_159), .B1(n_182), .B2(n_171), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_237), .A2(n_185), .B(n_171), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_244), .A2(n_185), .B1(n_171), .B2(n_173), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_237), .A2(n_185), .B(n_173), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_206), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_242), .A2(n_159), .B1(n_182), .B2(n_173), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_221), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_SL g285 ( .A1(n_234), .A2(n_203), .B(n_199), .C(n_197), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_244), .A2(n_149), .B1(n_199), .B2(n_197), .Y(n_286) );
AOI21x1_ASAP7_75t_L g287 ( .A1(n_244), .A2(n_203), .B(n_199), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_225), .A2(n_203), .B(n_197), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_240), .A2(n_149), .B(n_191), .C(n_202), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_206), .B(n_8), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_221), .B(n_9), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_206), .B(n_9), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_208), .B(n_10), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_244), .A2(n_191), .B1(n_202), .B2(n_13), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_208), .B(n_11), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_208), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_275), .B(n_270), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_267), .B(n_232), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_257), .B(n_214), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_271), .Y(n_300) );
OR2x6_ASAP7_75t_SL g301 ( .A(n_256), .B(n_230), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_257), .B(n_222), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_296), .Y(n_303) );
AOI21x1_ASAP7_75t_L g304 ( .A1(n_260), .A2(n_248), .B(n_253), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_287), .A2(n_255), .B(n_254), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_258), .A2(n_225), .B(n_227), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_266), .B(n_227), .Y(n_307) );
O2A1O1Ixp5_ASAP7_75t_SL g308 ( .A1(n_269), .A2(n_247), .B(n_241), .C(n_235), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_SL g309 ( .A1(n_277), .A2(n_223), .B(n_239), .C(n_236), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_266), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_261), .A2(n_239), .B(n_236), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_284), .B(n_259), .Y(n_312) );
AOI21xp5_ASAP7_75t_SL g313 ( .A1(n_280), .A2(n_232), .B(n_235), .Y(n_313) );
AO31x2_ASAP7_75t_L g314 ( .A1(n_289), .A2(n_239), .A3(n_236), .B(n_232), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_291), .B(n_216), .Y(n_315) );
NOR2xp67_ASAP7_75t_L g316 ( .A(n_262), .B(n_232), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_265), .A2(n_209), .B(n_249), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_262), .B(n_216), .Y(n_318) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_279), .A2(n_224), .B(n_219), .Y(n_319) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_268), .A2(n_215), .B(n_224), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_296), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_281), .A2(n_243), .B(n_191), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_272), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_300), .B(n_293), .Y(n_324) );
AOI22xp33_ASAP7_75t_SL g325 ( .A1(n_300), .A2(n_274), .B1(n_272), .B2(n_292), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_322), .Y(n_326) );
AO31x2_ASAP7_75t_L g327 ( .A1(n_306), .A2(n_310), .A3(n_311), .B(n_277), .Y(n_327) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_298), .B(n_272), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_304), .A2(n_286), .B(n_288), .Y(n_329) );
OAI21x1_ASAP7_75t_L g330 ( .A1(n_304), .A2(n_294), .B(n_290), .Y(n_330) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_313), .A2(n_285), .B(n_289), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_297), .B(n_295), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_308), .A2(n_273), .B(n_264), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_308), .A2(n_283), .B(n_278), .Y(n_334) );
OAI21x1_ASAP7_75t_L g335 ( .A1(n_322), .A2(n_282), .B(n_276), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_298), .B(n_276), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g337 ( .A(n_303), .B(n_282), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_312), .B(n_219), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_307), .B(n_216), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_303), .Y(n_340) );
INVx4_ASAP7_75t_L g341 ( .A(n_298), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_321), .B(n_323), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_305), .A2(n_285), .B(n_243), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_318), .Y(n_344) );
NAND3xp33_ASAP7_75t_L g345 ( .A(n_313), .B(n_263), .C(n_202), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_321), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
AOI21xp5_ASAP7_75t_SL g348 ( .A1(n_315), .A2(n_263), .B(n_213), .Y(n_348) );
AO21x2_ASAP7_75t_L g349 ( .A1(n_345), .A2(n_309), .B(n_305), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_344), .B(n_314), .Y(n_350) );
INVxp67_ASAP7_75t_L g351 ( .A(n_347), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_328), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_326), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_344), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_327), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_343), .A2(n_317), .B(n_319), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_346), .B(n_314), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_327), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_327), .B(n_314), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_346), .B(n_314), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_327), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_341), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_335), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_346), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_335), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_341), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_347), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_341), .B(n_314), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_339), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_343), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_340), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_339), .Y(n_380) );
OR2x6_ASAP7_75t_L g381 ( .A(n_345), .B(n_316), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_343), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_331), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_331), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_337), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_342), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_374), .B(n_355), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_361), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_350), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_350), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_354), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_351), .A2(n_324), .B(n_325), .C(n_302), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_374), .B(n_331), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_355), .B(n_332), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_374), .B(n_356), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_356), .B(n_331), .Y(n_397) );
BUFx2_ASAP7_75t_L g398 ( .A(n_359), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_366), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_358), .B(n_336), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_361), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_354), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_358), .B(n_336), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_351), .B(n_338), .C(n_332), .D(n_299), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_367), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_352), .Y(n_406) );
BUFx2_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_367), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_367), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_360), .B(n_336), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_360), .B(n_336), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_364), .B(n_328), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_364), .B(n_342), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_375), .Y(n_414) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_366), .B(n_348), .Y(n_415) );
AOI322xp5_ASAP7_75t_L g416 ( .A1(n_379), .A2(n_301), .A3(n_13), .B1(n_14), .B2(n_15), .C1(n_16), .C2(n_17), .Y(n_416) );
AO21x2_ASAP7_75t_L g417 ( .A1(n_383), .A2(n_348), .B(n_330), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_376), .B(n_337), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_376), .A2(n_320), .B1(n_323), .B2(n_342), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_365), .B(n_333), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_361), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_359), .B(n_333), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_361), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_352), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_379), .B(n_334), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_352), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_380), .B(n_334), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_375), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_373), .B(n_12), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_380), .B(n_334), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_372), .B(n_333), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_365), .B(n_330), .Y(n_432) );
NAND4xp25_ASAP7_75t_L g433 ( .A(n_362), .B(n_12), .C(n_15), .D(n_16), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_362), .B(n_330), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_359), .B(n_363), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_372), .B(n_17), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_368), .B(n_329), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_359), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_372), .B(n_19), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_361), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_386), .B(n_329), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_363), .B(n_20), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_363), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_366), .B(n_21), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_366), .A2(n_213), .B1(n_210), .B2(n_23), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_363), .B(n_317), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_361), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_363), .B(n_21), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_361), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_368), .B(n_22), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_404), .A2(n_384), .B1(n_383), .B2(n_385), .C(n_370), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_395), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_435), .B(n_383), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_399), .Y(n_454) );
INVxp67_ASAP7_75t_L g455 ( .A(n_444), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_396), .B(n_384), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_396), .B(n_384), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_393), .B(n_369), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_393), .B(n_387), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_387), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_389), .B(n_390), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_435), .B(n_369), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_400), .B(n_378), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_442), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_442), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_448), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_422), .B(n_381), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_422), .B(n_381), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_422), .B(n_381), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_400), .B(n_378), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_414), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_403), .B(n_378), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_394), .B(n_386), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_422), .B(n_381), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_403), .B(n_382), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_410), .B(n_382), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_410), .B(n_382), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_411), .B(n_371), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_411), .B(n_371), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_389), .B(n_385), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_399), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_399), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_390), .B(n_370), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_448), .B(n_366), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_397), .B(n_371), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_414), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_399), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_397), .B(n_371), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_406), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_398), .B(n_371), .Y(n_490) );
AND2x4_ASAP7_75t_SL g491 ( .A(n_406), .B(n_377), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_424), .Y(n_492) );
INVx5_ASAP7_75t_L g493 ( .A(n_388), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_398), .B(n_371), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_428), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_407), .B(n_371), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_395), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_428), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_426), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_388), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_418), .Y(n_501) );
CKINVDCx14_ASAP7_75t_R g502 ( .A(n_429), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_395), .Y(n_503) );
BUFx2_ASAP7_75t_SL g504 ( .A(n_426), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_407), .B(n_381), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_404), .B(n_377), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_438), .B(n_357), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_450), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_438), .B(n_357), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_443), .B(n_381), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_443), .B(n_357), .Y(n_511) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_424), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_420), .B(n_349), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_450), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_420), .B(n_349), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_391), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_412), .B(n_349), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_391), .Y(n_518) );
INVxp67_ASAP7_75t_SL g519 ( .A(n_405), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_405), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_408), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_412), .B(n_349), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_413), .B(n_377), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_426), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_402), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_402), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_408), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_413), .B(n_416), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_416), .B(n_377), .C(n_353), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_432), .B(n_349), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_433), .B(n_427), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_402), .Y(n_532) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_409), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_409), .Y(n_534) );
INVx4_ASAP7_75t_L g535 ( .A(n_388), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_427), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_432), .B(n_377), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_430), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_446), .B(n_353), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_430), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_437), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_421), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_459), .B(n_446), .Y(n_543) );
NAND2x1_ASAP7_75t_L g544 ( .A(n_454), .B(n_415), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_489), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_459), .B(n_446), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_452), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_460), .B(n_425), .Y(n_548) );
OR3x2_ASAP7_75t_L g549 ( .A(n_502), .B(n_433), .C(n_425), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_492), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_536), .B(n_434), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_458), .B(n_434), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_536), .B(n_431), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_538), .B(n_437), .Y(n_554) );
OR2x2_ASAP7_75t_SL g555 ( .A(n_487), .B(n_436), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
INVxp33_ASAP7_75t_L g557 ( .A(n_454), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_480), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_462), .B(n_458), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_519), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_481), .B(n_415), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_455), .B(n_392), .C(n_439), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_471), .Y(n_563) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_481), .B(n_445), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_462), .B(n_446), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_538), .B(n_419), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_471), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_482), .B(n_445), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_452), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_482), .B(n_441), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_456), .B(n_388), .Y(n_571) );
NOR2x1p5_ASAP7_75t_L g572 ( .A(n_529), .B(n_353), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_456), .B(n_401), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_457), .B(n_401), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_486), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_457), .B(n_441), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_540), .B(n_419), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_461), .B(n_449), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_540), .B(n_417), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_461), .B(n_417), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_497), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_501), .B(n_449), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_533), .B(n_449), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_495), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_495), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_539), .B(n_401), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_541), .B(n_417), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_539), .B(n_401), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_464), .B(n_447), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_498), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_497), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_505), .B(n_447), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_505), .B(n_447), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_528), .A2(n_440), .B1(n_423), .B2(n_421), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_498), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_465), .B(n_440), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_466), .B(n_440), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_503), .Y(n_599) );
AND2x2_ASAP7_75t_SL g600 ( .A(n_491), .B(n_423), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_503), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_491), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_516), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_537), .B(n_423), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_516), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_523), .B(n_421), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_537), .B(n_512), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_478), .B(n_417), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_531), .A2(n_22), .B(n_210), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_520), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_520), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_478), .B(n_25), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_479), .B(n_453), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_524), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_541), .B(n_26), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_521), .B(n_27), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_521), .B(n_28), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_527), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_504), .B(n_29), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_504), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_527), .B(n_30), .Y(n_621) );
OAI31xp33_ASAP7_75t_SL g622 ( .A1(n_451), .A2(n_32), .A3(n_33), .B(n_35), .Y(n_622) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_506), .A2(n_202), .B(n_243), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_518), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_479), .B(n_36), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_534), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_453), .B(n_38), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_508), .B(n_39), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_473), .B(n_42), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_513), .B(n_46), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_513), .B(n_47), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_499), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_453), .B(n_48), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_483), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_463), .B(n_50), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_515), .B(n_51), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_515), .B(n_52), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_525), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_530), .B(n_53), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_535), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_530), .B(n_56), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_560), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_562), .B(n_514), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_560), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_556), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_613), .B(n_488), .Y(n_646) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_614), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_622), .A2(n_499), .B(n_484), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_558), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_547), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_624), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_634), .B(n_485), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_622), .A2(n_505), .B(n_510), .Y(n_653) );
INVxp33_ASAP7_75t_L g654 ( .A(n_564), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_640), .B(n_467), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_545), .B(n_550), .Y(n_656) );
NOR2xp67_ASAP7_75t_L g657 ( .A(n_640), .B(n_535), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_568), .A2(n_535), .B1(n_507), .B2(n_509), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_559), .B(n_485), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_543), .B(n_488), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_569), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_584), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_595), .A2(n_507), .B(n_509), .C(n_511), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_546), .B(n_607), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_632), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_552), .B(n_463), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_581), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_551), .B(n_517), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_565), .B(n_467), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_592), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_551), .B(n_517), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_626), .Y(n_672) );
OAI32xp33_ASAP7_75t_L g673 ( .A1(n_557), .A2(n_483), .A3(n_500), .B1(n_511), .B2(n_490), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_599), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_601), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_563), .Y(n_676) );
INVx5_ASAP7_75t_L g677 ( .A(n_561), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_620), .B(n_493), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_587), .B(n_589), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_609), .A2(n_510), .B(n_468), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_571), .B(n_467), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_567), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_553), .B(n_522), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_553), .B(n_522), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_576), .B(n_476), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_566), .B(n_476), .Y(n_686) );
OAI322xp33_ASAP7_75t_L g687 ( .A1(n_548), .A2(n_470), .A3(n_475), .B1(n_472), .B2(n_477), .C1(n_525), .C2(n_526), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_566), .B(n_577), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_573), .B(n_468), .Y(n_689) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_609), .A2(n_510), .B1(n_493), .B2(n_468), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_580), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_575), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_583), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_585), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_574), .B(n_469), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_586), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_578), .B(n_477), .Y(n_697) );
BUFx2_ASAP7_75t_L g698 ( .A(n_602), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_577), .B(n_475), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_554), .B(n_591), .Y(n_700) );
OR2x2_ASAP7_75t_L g701 ( .A(n_606), .B(n_472), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_596), .Y(n_702) );
NOR2x2_ASAP7_75t_L g703 ( .A(n_549), .B(n_532), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_600), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_572), .A2(n_469), .B(n_474), .C(n_494), .Y(n_705) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_632), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_603), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_582), .B(n_470), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_604), .B(n_469), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_554), .B(n_496), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_605), .B(n_496), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_608), .B(n_474), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_638), .Y(n_713) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_580), .A2(n_474), .B(n_494), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_610), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_611), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_620), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_618), .B(n_490), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_570), .B(n_500), .Y(n_719) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_588), .Y(n_720) );
INVx1_ASAP7_75t_SL g721 ( .A(n_698), .Y(n_721) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_647), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_643), .A2(n_561), .B1(n_570), .B2(n_594), .Y(n_723) );
INVxp67_ASAP7_75t_L g724 ( .A(n_647), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_654), .A2(n_544), .B1(n_639), .B2(n_637), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_642), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_662), .B(n_597), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_644), .Y(n_728) );
OAI321xp33_ASAP7_75t_L g729 ( .A1(n_658), .A2(n_641), .A3(n_639), .B1(n_637), .B2(n_636), .C(n_630), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_662), .Y(n_730) );
NAND2x1_ASAP7_75t_L g731 ( .A(n_704), .B(n_619), .Y(n_731) );
NAND2x1_ASAP7_75t_L g732 ( .A(n_704), .B(n_594), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_651), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_672), .Y(n_734) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_665), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_700), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_665), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_653), .A2(n_555), .B1(n_636), .B2(n_631), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_676), .Y(n_739) );
INVx1_ASAP7_75t_SL g740 ( .A(n_717), .Y(n_740) );
NOR3xp33_ASAP7_75t_L g741 ( .A(n_643), .B(n_641), .C(n_630), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_688), .B(n_579), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_687), .A2(n_579), .B1(n_588), .B2(n_631), .C(n_628), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g744 ( .A1(n_654), .A2(n_629), .B(n_615), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_705), .A2(n_633), .B1(n_627), .B2(n_593), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_691), .B(n_598), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_691), .B(n_590), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_645), .B(n_593), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_649), .B(n_615), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_682), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_680), .A2(n_625), .B1(n_612), .B2(n_635), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_692), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_705), .A2(n_657), .B1(n_648), .B2(n_690), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_693), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_694), .Y(n_755) );
OAI21xp33_ASAP7_75t_L g756 ( .A1(n_714), .A2(n_623), .B(n_621), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_696), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_712), .B(n_500), .Y(n_758) );
AOI21xp33_ASAP7_75t_L g759 ( .A1(n_658), .A2(n_621), .B(n_617), .Y(n_759) );
OAI21xp33_ASAP7_75t_L g760 ( .A1(n_663), .A2(n_617), .B(n_616), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_690), .A2(n_493), .B1(n_616), .B2(n_542), .Y(n_761) );
O2A1O1Ixp5_ASAP7_75t_L g762 ( .A1(n_678), .A2(n_532), .B(n_526), .C(n_542), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_683), .B(n_493), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_709), .B(n_493), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_702), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_656), .A2(n_202), .B1(n_61), .B2(n_63), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_681), .B(n_59), .Y(n_767) );
AOI222xp33_ASAP7_75t_L g768 ( .A1(n_743), .A2(n_656), .B1(n_720), .B2(n_706), .C1(n_673), .C2(n_684), .Y(n_768) );
AOI211xp5_ASAP7_75t_L g769 ( .A1(n_753), .A2(n_678), .B(n_706), .C(n_655), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_721), .B(n_689), .Y(n_770) );
OAI222xp33_ASAP7_75t_L g771 ( .A1(n_738), .A2(n_703), .B1(n_677), .B2(n_655), .C1(n_666), .C2(n_686), .Y(n_771) );
OAI32xp33_ASAP7_75t_L g772 ( .A1(n_745), .A2(n_703), .A3(n_685), .B1(n_701), .B2(n_708), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_730), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g774 ( .A1(n_731), .A2(n_677), .B(n_720), .C(n_671), .Y(n_774) );
A2O1A1Ixp33_ASAP7_75t_L g775 ( .A1(n_732), .A2(n_677), .B(n_669), .C(n_664), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g776 ( .A1(n_736), .A2(n_699), .B1(n_668), .B2(n_652), .C(n_710), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_723), .A2(n_677), .B1(n_697), .B2(n_695), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_SL g778 ( .A1(n_724), .A2(n_718), .B(n_711), .C(n_716), .Y(n_778) );
INVx2_ASAP7_75t_SL g779 ( .A(n_740), .Y(n_779) );
AOI32xp33_ASAP7_75t_L g780 ( .A1(n_725), .A2(n_719), .A3(n_659), .B1(n_679), .B2(n_646), .Y(n_780) );
OAI332xp33_ASAP7_75t_L g781 ( .A1(n_725), .A2(n_715), .A3(n_707), .B1(n_670), .B2(n_675), .B3(n_674), .C1(n_667), .C2(n_661), .Y(n_781) );
AOI221xp5_ASAP7_75t_L g782 ( .A1(n_724), .A2(n_660), .B1(n_675), .B2(n_674), .C(n_670), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_722), .A2(n_667), .B(n_661), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_741), .A2(n_650), .B1(n_713), .B2(n_202), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_733), .B(n_650), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_758), .B(n_64), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g787 ( .A(n_762), .B(n_233), .Y(n_787) );
O2A1O1Ixp33_ASAP7_75t_L g788 ( .A1(n_722), .A2(n_66), .B(n_67), .C(n_68), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_746), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_742), .B(n_69), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_734), .B(n_71), .Y(n_791) );
OAI21xp5_ASAP7_75t_SL g792 ( .A1(n_741), .A2(n_72), .B(n_73), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_764), .B(n_74), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_789), .B(n_735), .Y(n_794) );
NAND2xp33_ASAP7_75t_L g795 ( .A(n_780), .B(n_760), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_776), .B(n_735), .Y(n_796) );
AOI221x1_ASAP7_75t_L g797 ( .A1(n_777), .A2(n_726), .B1(n_728), .B2(n_737), .C(n_759), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g798 ( .A(n_769), .B(n_729), .Y(n_798) );
OAI211xp5_ASAP7_75t_L g799 ( .A1(n_772), .A2(n_768), .B(n_774), .C(n_792), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_771), .A2(n_754), .B1(n_765), .B2(n_750), .C(n_752), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_781), .B(n_755), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_771), .A2(n_762), .B(n_756), .Y(n_802) );
AOI211x1_ASAP7_75t_SL g803 ( .A1(n_783), .A2(n_744), .B(n_749), .C(n_748), .Y(n_803) );
O2A1O1Ixp33_ASAP7_75t_L g804 ( .A1(n_779), .A2(n_757), .B(n_739), .C(n_747), .Y(n_804) );
OAI21xp33_ASAP7_75t_L g805 ( .A1(n_775), .A2(n_763), .B(n_761), .Y(n_805) );
O2A1O1Ixp33_ASAP7_75t_SL g806 ( .A1(n_782), .A2(n_727), .B(n_766), .C(n_751), .Y(n_806) );
NOR3xp33_ASAP7_75t_L g807 ( .A(n_788), .B(n_767), .C(n_77), .Y(n_807) );
OAI21xp5_ASAP7_75t_L g808 ( .A1(n_798), .A2(n_778), .B(n_784), .Y(n_808) );
NOR3xp33_ASAP7_75t_L g809 ( .A(n_799), .B(n_790), .C(n_787), .Y(n_809) );
NAND4xp25_ASAP7_75t_SL g810 ( .A(n_800), .B(n_770), .C(n_793), .D(n_786), .Y(n_810) );
OAI322xp33_ASAP7_75t_L g811 ( .A1(n_796), .A2(n_801), .A3(n_794), .B1(n_804), .B2(n_803), .C1(n_795), .C2(n_773), .Y(n_811) );
NAND4xp75_ASAP7_75t_L g812 ( .A(n_797), .B(n_791), .C(n_785), .D(n_79), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g813 ( .A(n_802), .B(n_785), .Y(n_813) );
INVx2_ASAP7_75t_SL g814 ( .A(n_805), .Y(n_814) );
NOR3x1_ASAP7_75t_L g815 ( .A(n_814), .B(n_806), .C(n_807), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_813), .Y(n_816) );
NOR3xp33_ASAP7_75t_L g817 ( .A(n_811), .B(n_791), .C(n_78), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_808), .B(n_76), .Y(n_818) );
NOR3xp33_ASAP7_75t_L g819 ( .A(n_817), .B(n_816), .C(n_818), .Y(n_819) );
NOR4xp75_ASAP7_75t_L g820 ( .A(n_815), .B(n_812), .C(n_809), .D(n_810), .Y(n_820) );
NOR2x1_ASAP7_75t_L g821 ( .A(n_817), .B(n_80), .Y(n_821) );
XNOR2x1_ASAP7_75t_L g822 ( .A(n_820), .B(n_81), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_819), .B(n_82), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_823), .B(n_821), .Y(n_824) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_822), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_825), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_824), .A2(n_233), .B1(n_86), .B2(n_87), .Y(n_827) );
INVx1_ASAP7_75t_SL g828 ( .A(n_826), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_828), .A2(n_827), .B1(n_233), .B2(n_91), .Y(n_829) );
AOI221x1_ASAP7_75t_L g830 ( .A1(n_829), .A2(n_85), .B1(n_89), .B2(n_94), .C(n_95), .Y(n_830) );
AOI21xp33_ASAP7_75t_L g831 ( .A1(n_830), .A2(n_96), .B(n_97), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_831), .A2(n_101), .B1(n_233), .B2(n_828), .Y(n_832) );
endmodule