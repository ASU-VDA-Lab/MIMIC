module real_jpeg_23049_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_1),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_10)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_1),
.A2(n_12),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_11),
.B1(n_13),
.B2(n_20),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_20),
.B1(n_42),
.B2(n_44),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_3),
.B(n_11),
.C(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_10),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_34),
.Y(n_6)
);

AOI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_24),
.B(n_33),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_21),
.Y(n_8)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_14),
.B(n_16),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_22),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_11),
.A2(n_13),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_19),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_40),
.B(n_45),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_48),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_29),
.B1(n_42),
.B2(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_53),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_50),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);


endmodule