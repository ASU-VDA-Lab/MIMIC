module real_jpeg_7085_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_525;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g197 ( 
.A(n_0),
.Y(n_197)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g285 ( 
.A(n_0),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_0),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_2),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_2),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_2),
.Y(n_328)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_2),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_2),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_3),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_3),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_3),
.A2(n_282),
.B1(n_364),
.B2(n_366),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_3),
.A2(n_282),
.B1(n_287),
.B2(n_390),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_L g454 ( 
.A1(n_3),
.A2(n_50),
.B1(n_282),
.B2(n_455),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_4),
.A2(n_211),
.B1(n_215),
.B2(n_216),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_4),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_4),
.A2(n_203),
.B1(n_215),
.B2(n_237),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_4),
.A2(n_89),
.B1(n_215),
.B2(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_4),
.A2(n_215),
.B1(n_327),
.B2(n_427),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_5),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_5),
.A2(n_99),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_5),
.A2(n_58),
.B1(n_99),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_5),
.A2(n_99),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_131),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_8),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_8),
.A2(n_171),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_8),
.A2(n_171),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_8),
.A2(n_150),
.B1(n_171),
.B2(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_11),
.A2(n_162),
.B1(n_164),
.B2(n_167),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_11),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_11),
.B(n_178),
.C(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_11),
.B(n_76),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_11),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_129),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_14),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_14),
.A2(n_92),
.B1(n_139),
.B2(n_144),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_14),
.A2(n_92),
.B1(n_180),
.B2(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_14),
.A2(n_92),
.B1(n_405),
.B2(n_409),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_15),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_15),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_15),
.A2(n_131),
.B1(n_190),
.B2(n_212),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_15),
.A2(n_190),
.B1(n_287),
.B2(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_15),
.A2(n_53),
.B1(n_60),
.B2(n_190),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_16),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_16),
.A2(n_54),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_16),
.A2(n_54),
.B1(n_211),
.B2(n_366),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_16),
.A2(n_54),
.B1(n_394),
.B2(n_396),
.Y(n_393)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_18),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_18),
.A2(n_61),
.B1(n_340),
.B2(n_342),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_18),
.A2(n_61),
.B1(n_133),
.B2(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_18),
.A2(n_61),
.B1(n_390),
.B2(n_440),
.Y(n_439)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_532),
.B(n_535),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_151),
.B(n_531),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_148),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_27),
.B(n_148),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_137),
.C(n_145),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_28),
.A2(n_29),
.B1(n_527),
.B2(n_528),
.Y(n_526)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_62),
.C(n_100),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_30),
.B(n_519),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_31),
.A2(n_55),
.B1(n_57),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_31),
.A2(n_55),
.B1(n_138),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_31),
.A2(n_352),
.B(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_31),
.A2(n_55),
.B1(n_400),
.B2(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_31),
.A2(n_49),
.B1(n_55),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_32),
.A2(n_349),
.B(n_351),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_32),
.B(n_353),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_32),
.A2(n_56),
.B(n_534),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_34),
.Y(n_330)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx8_ASAP7_75t_L g350 ( 
.A(n_35),
.Y(n_350)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_41),
.Y(n_332)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_44),
.Y(n_271)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_55),
.B(n_167),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_55),
.A2(n_426),
.B(n_458),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_56),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_56),
.B(n_454),
.Y(n_453)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_62),
.A2(n_100),
.B1(n_101),
.B2(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_62),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_85),
.B1(n_93),
.B2(n_94),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_63),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_63),
.A2(n_93),
.B1(n_305),
.B2(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_63),
.A2(n_93),
.B1(n_389),
.B2(n_393),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_63),
.A2(n_85),
.B1(n_93),
.B2(n_508),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_76),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_71),
.B2(n_74),
.Y(n_64)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_65),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_67),
.Y(n_274)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_70),
.Y(n_266)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_70),
.Y(n_326)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_70),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_77),
.B1(n_81),
.B2(n_83),
.Y(n_76)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_73),
.Y(n_292)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_75),
.Y(n_398)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_76),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

AOI22x1_ASAP7_75t_L g429 ( 
.A1(n_76),
.A2(n_146),
.B1(n_308),
.B2(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_76),
.A2(n_146),
.B1(n_438),
.B2(n_439),
.Y(n_437)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g408 ( 
.A(n_80),
.Y(n_408)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_86),
.B(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_88),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_88),
.Y(n_395)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_90),
.Y(n_275)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_93),
.B(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_93),
.A2(n_305),
.B(n_307),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_95),
.Y(n_287)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_100),
.A2(n_101),
.B1(n_506),
.B2(n_507),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_100),
.B(n_503),
.C(n_506),
.Y(n_514)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_128),
.B(n_130),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_161),
.B(n_168),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_102),
.A2(n_128),
.B1(n_210),
.B2(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_102),
.A2(n_168),
.B(n_262),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_102),
.A2(n_128),
.B1(n_363),
.B2(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_103),
.B(n_169),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_103),
.A2(n_129),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_103),
.A2(n_129),
.B1(n_385),
.B2(n_404),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_103),
.A2(n_129),
.B1(n_404),
.B2(n_445),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_110),
.B2(n_113),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g366 ( 
.A(n_105),
.Y(n_366)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_106),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_114),
.Y(n_290)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_115),
.A2(n_210),
.B(n_219),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_122),
.B2(n_124),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_121),
.Y(n_284)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_121),
.Y(n_313)
);

BUFx8_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_123),
.Y(n_239)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_128),
.A2(n_219),
.B(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_129),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_130),
.Y(n_445)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g293 ( 
.A(n_134),
.B(n_294),
.Y(n_293)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_136),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_136),
.Y(n_365)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_136),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_137),
.B(n_145),
.Y(n_528)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_140),
.B(n_167),
.Y(n_333)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_143),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_146),
.A2(n_265),
.B(n_272),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_146),
.B(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_146),
.A2(n_272),
.B(n_471),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_148),
.B(n_533),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_148),
.B(n_533),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_149),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_525),
.B(n_530),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_497),
.B(n_522),
.Y(n_152)
);

OAI311xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_369),
.A3(n_473),
.B1(n_491),
.C1(n_492),
.Y(n_153)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_319),
.B(n_368),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_296),
.B(n_318),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_256),
.B(n_295),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_222),
.B(n_255),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_185),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_159),
.B(n_185),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_172),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_160),
.A2(n_172),
.B1(n_173),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_160),
.Y(n_253)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_167),
.A2(n_194),
.B(n_200),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_SL g265 ( 
.A1(n_167),
.A2(n_266),
.B(n_267),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_SL g349 ( 
.A1(n_167),
.A2(n_333),
.B(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_182),
.Y(n_341)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_207),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_208),
.C(n_221),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_194),
.B(n_200),
.Y(n_186)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_193),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_194),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_194),
.A2(n_250),
.B1(n_375),
.B2(n_379),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_194),
.A2(n_379),
.B(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_202),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_195),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_195),
.A2(n_279),
.B1(n_312),
.B2(n_315),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_195),
.A2(n_315),
.B1(n_339),
.B2(n_423),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_197),
.Y(n_316)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_205),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_220),
.B2(n_221),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_245),
.B(n_254),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_234),
.B(n_244),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_233),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_230),
.Y(n_281)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_230),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_243),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_243),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_242),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_278),
.B(n_285),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_252),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_252),
.Y(n_254)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_258),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_276),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_263),
.C(n_276),
.Y(n_297)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI32xp33_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_287),
.A3(n_288),
.B1(n_291),
.B2(n_293),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx5_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_297),
.B(n_298),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_317),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_302),
.C(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_309),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_310),
.C(n_311),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_312),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_320),
.B(n_321),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_346),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_322)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_323),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_334),
.B2(n_335),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_325),
.B(n_334),
.Y(n_469)
);

OAI32xp33_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.A3(n_329),
.B1(n_331),
.B2(n_333),
.Y(n_325)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_340),
.Y(n_380)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_343),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_343),
.B(n_344),
.C(n_346),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_357),
.B2(n_367),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_347),
.B(n_358),
.C(n_362),
.Y(n_482)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_359),
.Y(n_471)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_459),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_370),
.A2(n_459),
.B(n_493),
.C(n_496),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_431),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_371),
.B(n_431),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_401),
.C(n_418),
.Y(n_371)
);

FAx1_ASAP7_75t_L g472 ( 
.A(n_372),
.B(n_401),
.CI(n_418),
.CON(n_472),
.SN(n_472)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_387),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_373),
.B(n_388),
.C(n_399),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_383),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_374),
.B(n_383),
.Y(n_465)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_375),
.Y(n_423)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_399),
.Y(n_387)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_413),
.B2(n_417),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_413),
.Y(n_449)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx8_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_413),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_413),
.A2(n_417),
.B1(n_451),
.B2(n_452),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_413),
.A2(n_449),
.B(n_452),
.Y(n_500)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_424),
.C(n_429),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_419),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_422),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_420),
.B(n_422),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_424),
.A2(n_425),
.B1(n_429),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx6_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_429),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_432),
.B(n_435),
.C(n_447),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_447),
.B2(n_448),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_443),
.B(n_446),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_444),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_439),
.Y(n_508)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_446),
.B(n_500),
.CI(n_501),
.CON(n_499),
.SN(n_499)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_446),
.B(n_500),
.C(n_501),
.Y(n_521)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_458),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_454),
.Y(n_504)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_472),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_472),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.C(n_466),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_461),
.A2(n_462),
.B1(n_465),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_465),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_484),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_469),
.C(n_470),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_467),
.A2(n_468),
.B1(n_470),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_472),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_486),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_475),
.A2(n_494),
.B(n_495),
.Y(n_493)
);

NOR2x1_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_483),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_483),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_480),
.C(n_482),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_489),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_480),
.A2(n_481),
.B1(n_482),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_482),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_488),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_511),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_510),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_499),
.B(n_510),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_499),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_503),
.B1(n_505),
.B2(n_509),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_502),
.A2(n_503),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_513),
.C(n_517),
.Y(n_529)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_505),
.Y(n_509)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_511),
.A2(n_523),
.B(n_524),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_512),
.B(n_521),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_521),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_529),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_529),
.Y(n_530)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

CKINVDCx14_ASAP7_75t_R g535 ( 
.A(n_536),
.Y(n_535)
);


endmodule