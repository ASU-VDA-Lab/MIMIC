module fake_netlist_6_2949_n_4429 (n_992, n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_968, n_909, n_580, n_762, n_1030, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_1008, n_1027, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_1033, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_1038, n_578, n_703, n_1003, n_144, n_365, n_978, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_951, n_783, n_106, n_725, n_952, n_999, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_994, n_677, n_969, n_988, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_974, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_1020, n_180, n_1009, n_1042, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_1032, n_845, n_255, n_807, n_1036, n_739, n_284, n_400, n_140, n_337, n_955, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_1026, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_963, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_1024, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_1018, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_1037, n_72, n_721, n_996, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_1015, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_360, n_945, n_977, n_603, n_1005, n_119, n_991, n_957, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_971, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_987, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_989, n_797, n_666, n_1016, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_1035, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_953, n_20, n_1004, n_1017, n_494, n_539, n_493, n_397, n_155, n_1022, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_576, n_1028, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_976, n_490, n_803, n_290, n_220, n_809, n_1011, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_986, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_990, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_998, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_972, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_962, n_1000, n_279, n_686, n_796, n_1041, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_984, n_411, n_503, n_716, n_152, n_623, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_1021, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_958, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_981, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_985, n_589, n_860, n_481, n_788, n_819, n_939, n_997, n_821, n_325, n_938, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_964, n_982, n_561, n_33, n_477, n_549, n_980, n_533, n_954, n_408, n_932, n_806, n_864, n_879, n_959, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_979, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_993, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_966, n_546, n_562, n_249, n_201, n_386, n_764, n_1039, n_556, n_159, n_1034, n_157, n_162, n_692, n_733, n_754, n_941, n_975, n_1031, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_970, n_560, n_1014, n_753, n_642, n_995, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_973, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_1029, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_967, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_1010, n_355, n_426, n_317, n_149, n_1040, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_1006, n_373, n_1012, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_1002, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_1019, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_965, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_983, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_961, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_950, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_956, n_960, n_531, n_827, n_1001, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_1025, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_1013, n_1023, n_194, n_664, n_171, n_949, n_678, n_192, n_57, n_169, n_1007, n_51, n_649, n_283, n_4429);

input n_992;
input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_968;
input n_909;
input n_580;
input n_762;
input n_1030;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_1008;
input n_1027;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_1033;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_1038;
input n_578;
input n_703;
input n_1003;
input n_144;
input n_365;
input n_978;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_951;
input n_783;
input n_106;
input n_725;
input n_952;
input n_999;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_994;
input n_677;
input n_969;
input n_988;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_974;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_1020;
input n_180;
input n_1009;
input n_1042;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_1032;
input n_845;
input n_255;
input n_807;
input n_1036;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_955;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_1026;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_963;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_1024;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_1018;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_1037;
input n_72;
input n_721;
input n_996;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_1015;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_945;
input n_977;
input n_603;
input n_1005;
input n_119;
input n_991;
input n_957;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_971;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_987;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_989;
input n_797;
input n_666;
input n_1016;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_1035;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_953;
input n_20;
input n_1004;
input n_1017;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_1022;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_576;
input n_1028;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_976;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_1011;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_986;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_990;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_998;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_972;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_962;
input n_1000;
input n_279;
input n_686;
input n_796;
input n_1041;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_984;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_1021;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_958;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_981;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_985;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_997;
input n_821;
input n_325;
input n_938;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_964;
input n_982;
input n_561;
input n_33;
input n_477;
input n_549;
input n_980;
input n_533;
input n_954;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_959;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_979;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_993;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_966;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_1039;
input n_556;
input n_159;
input n_1034;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_975;
input n_1031;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_970;
input n_560;
input n_1014;
input n_753;
input n_642;
input n_995;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_973;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_1029;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_967;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_1010;
input n_355;
input n_426;
input n_317;
input n_149;
input n_1040;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_1006;
input n_373;
input n_1012;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_1002;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_1019;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_965;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_983;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_961;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_950;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_956;
input n_960;
input n_531;
input n_827;
input n_1001;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_1025;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_1013;
input n_1023;
input n_194;
input n_664;
input n_171;
input n_949;
input n_678;
input n_192;
input n_57;
input n_169;
input n_1007;
input n_51;
input n_649;
input n_283;

output n_4429;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_2576;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1581;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_4372;
wire n_2451;
wire n_1620;
wire n_1738;
wire n_2243;
wire n_2324;
wire n_1575;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_2260;
wire n_1387;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_2847;
wire n_2557;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_2211;
wire n_1415;
wire n_1555;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_2247;
wire n_1711;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_2356;
wire n_1143;
wire n_1511;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_3979;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_2739;
wire n_2044;
wire n_1954;
wire n_2510;
wire n_1735;
wire n_1541;
wire n_2480;
wire n_1300;
wire n_3023;
wire n_3890;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_3063;
wire n_3048;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1455;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_4187;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2603;
wire n_2090;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_4125;
wire n_2625;
wire n_1400;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_4102;
wire n_4297;
wire n_2113;
wire n_1641;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_4314;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_3910;
wire n_1699;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_1530;
wire n_3798;
wire n_3488;
wire n_2811;
wire n_1543;
wire n_1302;
wire n_1068;
wire n_3732;
wire n_1599;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_2692;
wire n_1680;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_2714;
wire n_3092;
wire n_2245;
wire n_3055;
wire n_1289;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_1912;
wire n_1563;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_2818;
wire n_1359;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_3069;
wire n_3921;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_2311;
wire n_1386;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_1747;
wire n_3691;
wire n_4427;
wire n_3861;
wire n_2624;
wire n_4066;
wire n_4386;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_1801;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1214;
wire n_1654;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_4313;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_4169;
wire n_4055;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_2271;
wire n_3192;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3780;
wire n_3696;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_3337;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3431;
wire n_1767;
wire n_3450;
wire n_4002;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_3953;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_2913;
wire n_3614;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_4385;
wire n_1952;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_1932;
wire n_1101;
wire n_2535;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_2693;
wire n_1293;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_2767;
wire n_3793;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_3293;
wire n_1646;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_2897;
wire n_2537;
wire n_3970;
wire n_4389;
wire n_4345;
wire n_2554;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_2747;
wire n_1513;
wire n_3924;
wire n_3171;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_4284;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_2316;
wire n_1771;
wire n_4103;
wire n_4058;
wire n_3104;
wire n_3435;
wire n_3148;
wire n_2262;
wire n_3348;
wire n_3229;
wire n_4022;
wire n_2239;
wire n_3082;
wire n_1707;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_2842;
wire n_3580;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3775;
wire n_3537;
wire n_1176;
wire n_2134;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_3887;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4123;
wire n_1431;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_3835;
wire n_1571;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_2948;
wire n_1577;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_3996;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_4218;
wire n_4402;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_2372;
wire n_1490;
wire n_1568;
wire n_1299;
wire n_2896;
wire n_3837;
wire n_1650;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_2127;
wire n_1178;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_3191;
wire n_1626;
wire n_4005;
wire n_2482;
wire n_1507;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_2296;
wire n_2424;
wire n_1604;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_1774;
wire n_1475;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_1791;
wire n_3480;
wire n_1368;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_3641;
wire n_1837;
wire n_1314;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_4419;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1736;
wire n_1564;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_2416;
wire n_1427;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_3944;
wire n_3909;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3724;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_1286;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_1093;
wire n_4428;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3364;
wire n_3226;
wire n_3323;
wire n_4020;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_4404;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2502;
wire n_2131;
wire n_2226;
wire n_3646;
wire n_2801;
wire n_2920;
wire n_4015;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_3188;
wire n_3742;
wire n_1614;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_3284;
wire n_1806;
wire n_1267;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_2289;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2863;
wire n_1419;
wire n_1390;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_2627;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_3917;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3688;
wire n_3566;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_2181;
wire n_3751;
wire n_1594;
wire n_1869;
wire n_3625;
wire n_2911;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_2942;
wire n_1635;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_2327;
wire n_4374;
wire n_2201;
wire n_3919;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3194;
wire n_3250;
wire n_3276;
wire n_1934;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_3886;
wire n_2924;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_4420;
wire n_1510;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_2598;
wire n_1916;
wire n_1683;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_4234;
wire n_4304;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_3592;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_1108;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_4155;
wire n_2740;
wire n_4238;
wire n_3011;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_3137;
wire n_1535;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_3177;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_3238;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3529;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_2392;
wire n_1272;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_2050;
wire n_1472;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_3475;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_2789;
wire n_1352;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_2017;
wire n_1682;
wire n_1828;
wire n_2699;
wire n_2046;
wire n_2272;
wire n_3029;
wire n_2200;
wire n_1695;
wire n_4258;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_2376;
wire n_1405;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_2670;
wire n_1332;
wire n_2700;
wire n_4323;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_4209;
wire n_2871;
wire n_4135;
wire n_4279;
wire n_2688;
wire n_3858;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_2258;
wire n_1485;
wire n_1544;
wire n_1640;
wire n_4040;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_2390;
wire n_4007;
wire n_3712;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_3221;
wire n_1758;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3932;
wire n_3469;
wire n_3958;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_4205;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_2083;
wire n_1931;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1941;
wire n_1375;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_1045;
wire n_1794;
wire n_1962;
wire n_1236;
wire n_3506;
wire n_2398;
wire n_1725;
wire n_1928;
wire n_1559;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2888;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4170;
wire n_4143;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_4421;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_3621;
wire n_1476;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_2369;
wire n_1378;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_3343;
wire n_3303;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_4408;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_3027;
wire n_3231;
wire n_1554;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_4295;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_2020;
wire n_1643;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_2385;
wire n_1283;
wire n_4112;
wire n_1848;
wire n_1785;
wire n_1114;
wire n_1147;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3701;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_3473;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_2769;
wire n_1303;
wire n_4342;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1721;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_2180;
wire n_1689;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1347;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_4373;
wire n_1245;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_3811;
wire n_1656;
wire n_3494;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_2430;
wire n_1464;
wire n_1737;
wire n_3486;
wire n_1414;
wire n_3584;
wire n_4086;
wire n_2649;
wire n_2721;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_2743;
wire n_3962;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_4166;
wire n_1500;
wire n_1821;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_1253;
wire n_2242;
wire n_3362;
wire n_1266;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_1156;
wire n_1362;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_3285;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_3596;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_4316;
wire n_2233;
wire n_2723;
wire n_2440;
wire n_3521;
wire n_3233;
wire n_2800;
wire n_1710;
wire n_2161;
wire n_3496;
wire n_2805;
wire n_1301;
wire n_3310;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_3101;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_1574;
wire n_3989;
wire n_2478;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_4332;
wire n_4108;
wire n_1133;
wire n_3374;
wire n_1194;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_4293;
wire n_3552;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_1675;
wire n_2065;
wire n_2879;
wire n_3717;
wire n_4148;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_4263;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_3555;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1861;
wire n_3110;
wire n_1890;
wire n_1632;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_2280;
wire n_1557;
wire n_1833;
wire n_3903;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_1612;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_4129;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_2813;
wire n_1423;
wire n_1935;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_4030;
wire n_3113;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_155),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_959),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_568),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_470),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_98),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_814),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_831),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_846),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_981),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_133),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_784),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_834),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_781),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_239),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_38),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_346),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_172),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_1000),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_914),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_304),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_926),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_908),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_922),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_949),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_752),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_202),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_697),
.Y(n_1069)
);

BUFx10_ASAP7_75t_L g1070 ( 
.A(n_953),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_198),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_983),
.Y(n_1072)
);

CKINVDCx14_ASAP7_75t_R g1073 ( 
.A(n_89),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_848),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_771),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_1036),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1041),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_307),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_966),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_699),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_51),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_87),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_808),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_796),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_629),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_619),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_403),
.Y(n_1087)
);

CKINVDCx16_ASAP7_75t_R g1088 ( 
.A(n_634),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_458),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_925),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_755),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_901),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_927),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_821),
.Y(n_1094)
);

CKINVDCx16_ASAP7_75t_R g1095 ( 
.A(n_818),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_95),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_152),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_895),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_2),
.Y(n_1099)
);

CKINVDCx11_ASAP7_75t_R g1100 ( 
.A(n_548),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_732),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_616),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1016),
.Y(n_1103)
);

BUFx10_ASAP7_75t_L g1104 ( 
.A(n_83),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_820),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_954),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_210),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_412),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_943),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_297),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_178),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_98),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_854),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_946),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_505),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_859),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_944),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1030),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1001),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_241),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_254),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_786),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_32),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_493),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_802),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_454),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_647),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_94),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_920),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_891),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_333),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_550),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_731),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_720),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_27),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_969),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1020),
.Y(n_1137)
);

CKINVDCx16_ASAP7_75t_R g1138 ( 
.A(n_909),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_342),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_871),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_801),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_72),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_948),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_940),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_641),
.Y(n_1145)
);

BUFx10_ASAP7_75t_L g1146 ( 
.A(n_797),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_919),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1012),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_806),
.Y(n_1149)
);

BUFx10_ASAP7_75t_L g1150 ( 
.A(n_540),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_127),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_541),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_868),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_55),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_730),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_319),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1014),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_898),
.Y(n_1158)
);

CKINVDCx14_ASAP7_75t_R g1159 ( 
.A(n_692),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_960),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_701),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_313),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1002),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_842),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_826),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_825),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_776),
.Y(n_1167)
);

CKINVDCx16_ASAP7_75t_R g1168 ( 
.A(n_631),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_838),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_232),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_545),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_179),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1028),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_413),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_601),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_764),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_758),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_119),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_765),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_159),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_673),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_106),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_497),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_870),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_836),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_500),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_676),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_492),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_162),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_856),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_775),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_725),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_320),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_748),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_777),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_217),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_935),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_303),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_408),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_439),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_885),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_961),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_760),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_886),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_711),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_809),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_867),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_811),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_512),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_890),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_945),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_82),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_180),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_167),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_862),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_215),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_710),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_267),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_987),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_495),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_242),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_20),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_804),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_536),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_729),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_372),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_16),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_999),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_717),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_557),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_687),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_988),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_652),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_32),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_897),
.Y(n_1235)
);

CKINVDCx16_ASAP7_75t_R g1236 ( 
.A(n_572),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_298),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_882),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_718),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_253),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_912),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_979),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_719),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_104),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_994),
.Y(n_1245)
);

CKINVDCx16_ASAP7_75t_R g1246 ( 
.A(n_659),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_700),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_428),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_532),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_481),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1027),
.Y(n_1251)
);

BUFx10_ASAP7_75t_L g1252 ( 
.A(n_500),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_6),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_566),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_532),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_312),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_414),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_933),
.Y(n_1258)
);

BUFx10_ASAP7_75t_L g1259 ( 
.A(n_315),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_102),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_751),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_385),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_248),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_875),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_894),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_989),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1039),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_501),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_649),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_174),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_112),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_335),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_505),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_709),
.Y(n_1274)
);

BUFx2_ASAP7_75t_SL g1275 ( 
.A(n_575),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_726),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_513),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_887),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_321),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_478),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_990),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_602),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_447),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_918),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_923),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_191),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_829),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_782),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1017),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_26),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_975),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_739),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_29),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_696),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_300),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_789),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_850),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_16),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_156),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_233),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_337),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_851),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_228),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_90),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_873),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_996),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_600),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_705),
.Y(n_1308)
);

CKINVDCx16_ASAP7_75t_R g1309 ( 
.A(n_309),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_400),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_624),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_30),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_794),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_448),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_160),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1042),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_968),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_89),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_917),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_244),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1032),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_231),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_998),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_963),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_203),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_600),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_333),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_708),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_905),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_386),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_358),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_625),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1011),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_55),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_971),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1022),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_936),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_876),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_99),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_587),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1023),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_807),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1040),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_840),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_861),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_673),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_772),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_892),
.Y(n_1348)
);

CKINVDCx14_ASAP7_75t_R g1349 ( 
.A(n_767),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_586),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_422),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_587),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_26),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_900),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_783),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_938),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_835),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_56),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_972),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_924),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1024),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_294),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1033),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1013),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_992),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_141),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_640),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_947),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_409),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_795),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_565),
.Y(n_1371)
);

BUFx5_ASAP7_75t_L g1372 ( 
.A(n_881),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_866),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1034),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_617),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_932),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_203),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_693),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_770),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_292),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_93),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_52),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_958),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_478),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_986),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_49),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_196),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_627),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_787),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_553),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_658),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_727),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_827),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_910),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_965),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_941),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_125),
.Y(n_1397)
);

CKINVDCx14_ASAP7_75t_R g1398 ( 
.A(n_340),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_307),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_290),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_832),
.Y(n_1401)
);

BUFx10_ASAP7_75t_L g1402 ( 
.A(n_92),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_753),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_166),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_186),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_937),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_790),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_763),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_913),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_830),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_984),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_675),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_196),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_491),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_14),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_25),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_701),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1037),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_779),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_49),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_278),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_390),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_126),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_583),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_921),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_172),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_817),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_145),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_716),
.Y(n_1429)
);

INVx2_ASAP7_75t_SL g1430 ( 
.A(n_619),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_525),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_691),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_398),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_810),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_967),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_696),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_889),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_762),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_823),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_99),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_27),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_931),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_208),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_792),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_241),
.Y(n_1445)
);

BUFx8_ASAP7_75t_SL g1446 ( 
.A(n_877),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_644),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_844),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_843),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_915),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_85),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_691),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_952),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_930),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_880),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_675),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_734),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_833),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_855),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_712),
.Y(n_1460)
);

BUFx10_ASAP7_75t_L g1461 ( 
.A(n_1025),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_198),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_238),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_604),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_377),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_528),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_433),
.Y(n_1467)
);

BUFx10_ASAP7_75t_L g1468 ( 
.A(n_1007),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_341),
.Y(n_1469)
);

BUFx10_ASAP7_75t_L g1470 ( 
.A(n_51),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_857),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_815),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_982),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_363),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_956),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_813),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_819),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_929),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_302),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_991),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_962),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_688),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_759),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1004),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_189),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_893),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1029),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_538),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_544),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_403),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_757),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_899),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_303),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_158),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_481),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_255),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_535),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_476),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1010),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_476),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_614),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_471),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_828),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_487),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_139),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_108),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_837),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_275),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1026),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_768),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_416),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_896),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_452),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_653),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_120),
.Y(n_1515)
);

CKINVDCx16_ASAP7_75t_R g1516 ( 
.A(n_699),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_42),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1031),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_550),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_43),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_158),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_697),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_467),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_147),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_977),
.Y(n_1525)
);

CKINVDCx14_ASAP7_75t_R g1526 ( 
.A(n_687),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_741),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_494),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_995),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_703),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_242),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_179),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_793),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_443),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_47),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1005),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_452),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_656),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_706),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_566),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_799),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_847),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_197),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_140),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_798),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_902),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_54),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_409),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_774),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_502),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_483),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_335),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_578),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_883),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_705),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_845),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_531),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_597),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_997),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_525),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_708),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_985),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_282),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_375),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_791),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_146),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_724),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_46),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_442),
.Y(n_1569)
);

BUFx10_ASAP7_75t_L g1570 ( 
.A(n_978),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_744),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_432),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_124),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_928),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_389),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_750),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_147),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_800),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_723),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_644),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_297),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1009),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_803),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_288),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_336),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_274),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_119),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_146),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_102),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_400),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_974),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_110),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_865),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_746),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_816),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_571),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_955),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_278),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_869),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_159),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_300),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_373),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_904),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_993),
.Y(n_1604)
);

CKINVDCx14_ASAP7_75t_R g1605 ( 
.A(n_534),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_87),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_633),
.Y(n_1607)
);

CKINVDCx16_ASAP7_75t_R g1608 ( 
.A(n_878),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_137),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_521),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_721),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_217),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_308),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_907),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_860),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_839),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_471),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_510),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_864),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_745),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_389),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_580),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_264),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_470),
.Y(n_1624)
);

CKINVDCx20_ASAP7_75t_R g1625 ( 
.A(n_950),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_349),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_511),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_567),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_554),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_373),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_934),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_113),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_553),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_853),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_378),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_161),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_668),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_888),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_747),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_396),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_528),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_96),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_343),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_858),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_253),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_91),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1021),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_903),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_736),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_884),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_714),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_489),
.Y(n_1652)
);

BUFx10_ASAP7_75t_L g1653 ( 
.A(n_2),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_265),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_165),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_79),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_824),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_190),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_484),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_202),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_50),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_841),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_156),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_357),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_970),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_513),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_366),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_323),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_714),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_615),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_421),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_498),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_715),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_209),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_805),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_707),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_187),
.Y(n_1677)
);

CKINVDCx16_ASAP7_75t_R g1678 ( 
.A(n_728),
.Y(n_1678)
);

CKINVDCx16_ASAP7_75t_R g1679 ( 
.A(n_766),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1038),
.Y(n_1680)
);

CKINVDCx20_ASAP7_75t_R g1681 ( 
.A(n_287),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_348),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_976),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_852),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_493),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_19),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_957),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_662),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_260),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_365),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_980),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_647),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_410),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_638),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_879),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_291),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_135),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_495),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_724),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_171),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_874),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_740),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_186),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_906),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_812),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_267),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_301),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_720),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_330),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_916),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_773),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_951),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_973),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_351),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_14),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_340),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_822),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_213),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1035),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1019),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_646),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_184),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_964),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1018),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_594),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_713),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_540),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_756),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_357),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_402),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_501),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_84),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_375),
.Y(n_1733)
);

CKINVDCx20_ASAP7_75t_R g1734 ( 
.A(n_334),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_106),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_227),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_249),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_743),
.Y(n_1738)
);

CKINVDCx20_ASAP7_75t_R g1739 ( 
.A(n_255),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_939),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_221),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_780),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_514),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_849),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_453),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_325),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_411),
.Y(n_1747)
);

BUFx3_ASAP7_75t_L g1748 ( 
.A(n_722),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_620),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1003),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1015),
.Y(n_1751)
);

CKINVDCx20_ASAP7_75t_R g1752 ( 
.A(n_280),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_175),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_769),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_778),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_559),
.Y(n_1756)
);

CKINVDCx16_ASAP7_75t_R g1757 ( 
.A(n_788),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_243),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_754),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_162),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_309),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_761),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_143),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_239),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_607),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_282),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_863),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_742),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_942),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_785),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_735),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_749),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_372),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_690),
.Y(n_1774)
);

CKINVDCx5p33_ASAP7_75t_R g1775 ( 
.A(n_441),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1006),
.Y(n_1776)
);

CKINVDCx20_ASAP7_75t_R g1777 ( 
.A(n_911),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_872),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_618),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_593),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1008),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_522),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_1064),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1523),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1523),
.Y(n_1785)
);

CKINVDCx16_ASAP7_75t_R g1786 ( 
.A(n_1088),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1131),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1131),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1081),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1131),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1180),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1180),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1180),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1496),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1496),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1496),
.Y(n_1796)
);

INVxp33_ASAP7_75t_SL g1797 ( 
.A(n_1268),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1587),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1587),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1587),
.Y(n_1800)
);

BUFx3_ASAP7_75t_L g1801 ( 
.A(n_1070),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1446),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1100),
.Y(n_1803)
);

INVxp33_ASAP7_75t_SL g1804 ( 
.A(n_1413),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1645),
.Y(n_1805)
);

CKINVDCx20_ASAP7_75t_R g1806 ( 
.A(n_1777),
.Y(n_1806)
);

INVxp33_ASAP7_75t_SL g1807 ( 
.A(n_1515),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1645),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1645),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1126),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1125),
.Y(n_1811)
);

INVxp67_ASAP7_75t_SL g1812 ( 
.A(n_1356),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_1065),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1070),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1087),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1156),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1372),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1135),
.Y(n_1818)
);

CKINVDCx16_ASAP7_75t_R g1819 ( 
.A(n_1168),
.Y(n_1819)
);

INVxp67_ASAP7_75t_SL g1820 ( 
.A(n_1075),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1044),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1206),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1048),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1187),
.Y(n_1824)
);

INVxp33_ASAP7_75t_L g1825 ( 
.A(n_1573),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1193),
.Y(n_1826)
);

INVxp33_ASAP7_75t_SL g1827 ( 
.A(n_1579),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1200),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1218),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1372),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1049),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1050),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1271),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1330),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1351),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_1079),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1421),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1500),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1589),
.Y(n_1839)
);

INVxp33_ASAP7_75t_SL g1840 ( 
.A(n_1607),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1164),
.Y(n_1841)
);

INVxp67_ASAP7_75t_SL g1842 ( 
.A(n_1338),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1051),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1622),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1666),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1694),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1236),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1730),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1748),
.Y(n_1849)
);

CKINVDCx20_ASAP7_75t_R g1850 ( 
.A(n_1167),
.Y(n_1850)
);

CKINVDCx14_ASAP7_75t_R g1851 ( 
.A(n_1073),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1774),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1054),
.Y(n_1853)
);

INVxp67_ASAP7_75t_SL g1854 ( 
.A(n_1492),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1045),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1055),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1046),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1372),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1372),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1062),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1253),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1069),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1097),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1111),
.Y(n_1864)
);

INVxp33_ASAP7_75t_SL g1865 ( 
.A(n_1290),
.Y(n_1865)
);

CKINVDCx20_ASAP7_75t_R g1866 ( 
.A(n_1194),
.Y(n_1866)
);

INVxp33_ASAP7_75t_SL g1867 ( 
.A(n_1346),
.Y(n_1867)
);

INVxp67_ASAP7_75t_SL g1868 ( 
.A(n_1638),
.Y(n_1868)
);

CKINVDCx20_ASAP7_75t_R g1869 ( 
.A(n_1335),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1120),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1124),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1128),
.Y(n_1872)
);

INVxp67_ASAP7_75t_SL g1873 ( 
.A(n_1265),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1159),
.B(n_1),
.Y(n_1874)
);

INVxp67_ASAP7_75t_SL g1875 ( 
.A(n_1265),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1142),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1060),
.Y(n_1877)
);

CKINVDCx14_ASAP7_75t_R g1878 ( 
.A(n_1398),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1152),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1170),
.Y(n_1880)
);

CKINVDCx16_ASAP7_75t_R g1881 ( 
.A(n_1246),
.Y(n_1881)
);

INVxp33_ASAP7_75t_SL g1882 ( 
.A(n_1388),
.Y(n_1882)
);

CKINVDCx20_ASAP7_75t_R g1883 ( 
.A(n_1354),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1309),
.Y(n_1884)
);

INVxp33_ASAP7_75t_L g1885 ( 
.A(n_1432),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1171),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1067),
.Y(n_1887)
);

INVx1_ASAP7_75t_SL g1888 ( 
.A(n_1519),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1172),
.Y(n_1889)
);

INVxp67_ASAP7_75t_SL g1890 ( 
.A(n_1106),
.Y(n_1890)
);

INVxp33_ASAP7_75t_SL g1891 ( 
.A(n_1709),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1174),
.Y(n_1892)
);

INVxp67_ASAP7_75t_SL g1893 ( 
.A(n_1190),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_1408),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1074),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1182),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1192),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1795),
.Y(n_1898)
);

AOI22x1_ASAP7_75t_SL g1899 ( 
.A1(n_1783),
.A2(n_1085),
.B1(n_1133),
.B2(n_1080),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1801),
.B(n_1305),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1821),
.B(n_1349),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1851),
.B(n_1526),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1787),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1788),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1865),
.A2(n_1605),
.B1(n_1678),
.B2(n_1516),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1878),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1796),
.Y(n_1907)
);

XNOR2xp5_ASAP7_75t_L g1908 ( 
.A(n_1806),
.B(n_1154),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1790),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1814),
.B(n_1406),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1791),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1867),
.A2(n_1138),
.B1(n_1608),
.B2(n_1095),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1890),
.B(n_1679),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1882),
.A2(n_1757),
.B1(n_1308),
.B2(n_1520),
.Y(n_1914)
);

OA21x2_ASAP7_75t_L g1915 ( 
.A1(n_1873),
.A2(n_1662),
.B(n_1472),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1893),
.B(n_1437),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1823),
.B(n_1831),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1792),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1796),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1793),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_SL g1921 ( 
.A(n_1789),
.B(n_1146),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1847),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1832),
.B(n_1166),
.Y(n_1923)
);

AOI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1891),
.A2(n_1459),
.B1(n_1471),
.B2(n_1434),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1843),
.B(n_1853),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1794),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1810),
.B(n_1240),
.Y(n_1927)
);

CKINVDCx8_ASAP7_75t_R g1928 ( 
.A(n_1786),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1798),
.Y(n_1929)
);

BUFx2_ASAP7_75t_L g1930 ( 
.A(n_1803),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1799),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1820),
.B(n_1822),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1884),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1797),
.A2(n_1198),
.B1(n_1227),
.B2(n_1188),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1800),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1818),
.Y(n_1936)
);

INVx5_ASAP7_75t_L g1937 ( 
.A(n_1861),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1805),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1808),
.Y(n_1939)
);

INVx6_ASAP7_75t_L g1940 ( 
.A(n_1819),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1842),
.B(n_1525),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1809),
.Y(n_1942)
);

BUFx6f_ASAP7_75t_L g1943 ( 
.A(n_1852),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1815),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1784),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1855),
.Y(n_1946)
);

AOI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1804),
.A2(n_1510),
.B1(n_1512),
.B2(n_1475),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1807),
.A2(n_1668),
.B1(n_1685),
.B2(n_1248),
.Y(n_1948)
);

AND2x2_ASAP7_75t_SL g1949 ( 
.A(n_1881),
.B(n_1047),
.Y(n_1949)
);

INVx4_ASAP7_75t_L g1950 ( 
.A(n_1856),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1877),
.B(n_1518),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1854),
.B(n_1631),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1857),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1868),
.B(n_1179),
.Y(n_1954)
);

OA21x2_ASAP7_75t_L g1955 ( 
.A1(n_1875),
.A2(n_1061),
.B(n_1053),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1811),
.B(n_1297),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1887),
.Y(n_1957)
);

OA21x2_ASAP7_75t_L g1958 ( 
.A1(n_1785),
.A2(n_1066),
.B(n_1063),
.Y(n_1958)
);

NOR2x1_ASAP7_75t_L g1959 ( 
.A(n_1817),
.B(n_1072),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1860),
.Y(n_1960)
);

XNOR2xp5_ASAP7_75t_L g1961 ( 
.A(n_1813),
.B(n_1229),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1895),
.B(n_1191),
.Y(n_1962)
);

OA21x2_ASAP7_75t_L g1963 ( 
.A1(n_1830),
.A2(n_1084),
.B(n_1077),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1812),
.B(n_1146),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1816),
.B(n_1219),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1862),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1863),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1824),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1826),
.B(n_1251),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1864),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1870),
.Y(n_1971)
);

AND2x2_ASAP7_75t_SL g1972 ( 
.A(n_1874),
.B(n_1071),
.Y(n_1972)
);

CKINVDCx20_ASAP7_75t_R g1973 ( 
.A(n_1836),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1888),
.B(n_1345),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1828),
.B(n_1284),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1871),
.Y(n_1976)
);

INVx4_ASAP7_75t_L g1977 ( 
.A(n_1802),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1829),
.B(n_1306),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1833),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1834),
.B(n_1324),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1835),
.B(n_1343),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1837),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1872),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1838),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1876),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1879),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1880),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1858),
.A2(n_1859),
.B(n_1450),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1827),
.A2(n_1625),
.B1(n_1649),
.B2(n_1582),
.Y(n_1989)
);

AND2x2_ASAP7_75t_SL g1990 ( 
.A(n_1839),
.B(n_1257),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1886),
.Y(n_1991)
);

BUFx6f_ASAP7_75t_L g1992 ( 
.A(n_1889),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1841),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1892),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1844),
.B(n_1453),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1896),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1845),
.Y(n_1997)
);

OAI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1840),
.A2(n_1052),
.B1(n_1056),
.B2(n_1043),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1897),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1846),
.B(n_1401),
.Y(n_2000)
);

BUFx8_ASAP7_75t_SL g2001 ( 
.A(n_1894),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1848),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1849),
.B(n_1177),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1850),
.Y(n_2004)
);

INVxp67_ASAP7_75t_L g2005 ( 
.A(n_1885),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1825),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1866),
.B(n_1461),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1869),
.B(n_1461),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1883),
.B(n_1509),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1795),
.Y(n_2010)
);

NAND2xp33_ASAP7_75t_L g2011 ( 
.A(n_1821),
.B(n_1057),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1801),
.B(n_1776),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1851),
.B(n_1468),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1795),
.Y(n_2014)
);

OA21x2_ASAP7_75t_L g2015 ( 
.A1(n_1873),
.A2(n_1094),
.B(n_1093),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1796),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1801),
.Y(n_2017)
);

BUFx2_ASAP7_75t_L g2018 ( 
.A(n_1851),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1795),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1795),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1795),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1801),
.B(n_1103),
.Y(n_2022)
);

BUFx8_ASAP7_75t_L g2023 ( 
.A(n_1818),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1821),
.B(n_1533),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1851),
.B(n_1468),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1821),
.B(n_1647),
.Y(n_2026)
);

BUFx8_ASAP7_75t_L g2027 ( 
.A(n_1818),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1865),
.A2(n_1704),
.B1(n_1720),
.B2(n_1717),
.Y(n_2028)
);

OAI21x1_ASAP7_75t_L g2029 ( 
.A1(n_1817),
.A2(n_1778),
.B(n_1772),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1821),
.B(n_1116),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1795),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1821),
.B(n_1119),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1821),
.B(n_1122),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1821),
.B(n_1130),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1795),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1801),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1801),
.B(n_1137),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_1847),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1795),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1847),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1795),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1795),
.Y(n_2042)
);

OAI21x1_ASAP7_75t_L g2043 ( 
.A1(n_1817),
.A2(n_1148),
.B(n_1147),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_SL g2044 ( 
.A1(n_1865),
.A2(n_1249),
.B1(n_1294),
.B2(n_1237),
.Y(n_2044)
);

BUFx2_ASAP7_75t_L g2045 ( 
.A(n_1851),
.Y(n_2045)
);

OAI22xp5_ASAP7_75t_SL g2046 ( 
.A1(n_1865),
.A2(n_1315),
.B1(n_1320),
.B2(n_1314),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1795),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1851),
.B(n_1570),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1865),
.A2(n_1723),
.B1(n_1672),
.B2(n_1059),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1795),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1795),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1865),
.A2(n_1068),
.B1(n_1078),
.B2(n_1058),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1795),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1817),
.A2(n_1158),
.B(n_1149),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_1801),
.B(n_1163),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_1851),
.B(n_1570),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1796),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1865),
.A2(n_1082),
.B1(n_1089),
.B2(n_1086),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1795),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1821),
.B(n_1173),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1821),
.B(n_1185),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1795),
.Y(n_2062)
);

BUFx6f_ASAP7_75t_L g2063 ( 
.A(n_1795),
.Y(n_2063)
);

BUFx8_ASAP7_75t_L g2064 ( 
.A(n_1818),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1795),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1795),
.Y(n_2066)
);

AOI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_1865),
.A2(n_1099),
.B1(n_1102),
.B2(n_1096),
.Y(n_2067)
);

INVx3_ASAP7_75t_L g2068 ( 
.A(n_1796),
.Y(n_2068)
);

CKINVDCx20_ASAP7_75t_R g2069 ( 
.A(n_1783),
.Y(n_2069)
);

HB1xp67_ASAP7_75t_L g2070 ( 
.A(n_1847),
.Y(n_2070)
);

BUFx8_ASAP7_75t_L g2071 ( 
.A(n_1818),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1795),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_1801),
.B(n_1195),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1795),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_L g2075 ( 
.A(n_1795),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1851),
.B(n_1255),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1795),
.Y(n_2077)
);

OAI22xp5_ASAP7_75t_SL g2078 ( 
.A1(n_1865),
.A2(n_1382),
.B1(n_1452),
.B2(n_1353),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1795),
.Y(n_2079)
);

CKINVDCx6p67_ASAP7_75t_R g2080 ( 
.A(n_1786),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1821),
.Y(n_2081)
);

INVx4_ASAP7_75t_L g2082 ( 
.A(n_1821),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1821),
.B(n_1201),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1795),
.Y(n_2084)
);

BUFx8_ASAP7_75t_SL g2085 ( 
.A(n_1803),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1795),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1851),
.B(n_1414),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1795),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1795),
.Y(n_2089)
);

BUFx8_ASAP7_75t_L g2090 ( 
.A(n_1818),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_1795),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1851),
.B(n_1422),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1795),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1801),
.B(n_1202),
.Y(n_2094)
);

INVx4_ASAP7_75t_L g2095 ( 
.A(n_1821),
.Y(n_2095)
);

BUFx12f_ASAP7_75t_L g2096 ( 
.A(n_1802),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1795),
.Y(n_2097)
);

BUFx6f_ASAP7_75t_L g2098 ( 
.A(n_1795),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1795),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1795),
.Y(n_2100)
);

CKINVDCx20_ASAP7_75t_R g2101 ( 
.A(n_1783),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1795),
.Y(n_2102)
);

INVx3_ASAP7_75t_L g2103 ( 
.A(n_1796),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1786),
.B(n_1104),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1821),
.B(n_1215),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1795),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1795),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_1821),
.B(n_1238),
.Y(n_2108)
);

INVx3_ASAP7_75t_L g2109 ( 
.A(n_1796),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_1847),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1796),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1821),
.B(n_1241),
.Y(n_2112)
);

BUFx3_ASAP7_75t_L g2113 ( 
.A(n_1815),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1821),
.B(n_1242),
.Y(n_2114)
);

INVx3_ASAP7_75t_L g2115 ( 
.A(n_1796),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1795),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1795),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1795),
.Y(n_2118)
);

INVx2_ASAP7_75t_SL g2119 ( 
.A(n_1801),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1801),
.B(n_1245),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1795),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1821),
.B(n_1261),
.Y(n_2122)
);

CKINVDCx5p33_ASAP7_75t_R g2123 ( 
.A(n_1821),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1786),
.B(n_1104),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1821),
.B(n_1281),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_1796),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1795),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1851),
.B(n_1429),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1821),
.B(n_1296),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_1795),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_SL g2131 ( 
.A1(n_1865),
.A2(n_1467),
.B1(n_1504),
.B2(n_1465),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1795),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1795),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_1796),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1795),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1795),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1795),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1795),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1795),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_1796),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1795),
.Y(n_2141)
);

INVx3_ASAP7_75t_L g2142 ( 
.A(n_1796),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1795),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_1801),
.B(n_1329),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1795),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1795),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1795),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1795),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1795),
.Y(n_2149)
);

XNOR2xp5_ASAP7_75t_L g2150 ( 
.A(n_1783),
.B(n_1506),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1851),
.B(n_1430),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1795),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1795),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1795),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1851),
.B(n_1600),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_1821),
.B(n_1333),
.Y(n_2156)
);

OA21x2_ASAP7_75t_L g2157 ( 
.A1(n_1873),
.A2(n_1341),
.B(n_1336),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1795),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_1796),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1795),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1796),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1851),
.B(n_1692),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1821),
.B(n_1357),
.Y(n_2163)
);

INVx3_ASAP7_75t_L g2164 ( 
.A(n_1796),
.Y(n_2164)
);

INVx4_ASAP7_75t_L g2165 ( 
.A(n_1821),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1795),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1795),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_1847),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1821),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2014),
.Y(n_2170)
);

AND3x2_ASAP7_75t_L g2171 ( 
.A(n_1921),
.B(n_1399),
.C(n_1322),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2014),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1960),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_1927),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_1907),
.Y(n_2175)
);

OAI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2049),
.A2(n_1108),
.B1(n_1110),
.B2(n_1107),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2041),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1913),
.B(n_1076),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1962),
.B(n_1112),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1907),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1966),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2024),
.B(n_1083),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1974),
.B(n_1090),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1932),
.B(n_1150),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2026),
.B(n_1091),
.Y(n_2185)
);

INVx3_ASAP7_75t_L g2186 ( 
.A(n_1919),
.Y(n_2186)
);

NAND2xp33_ASAP7_75t_SL g2187 ( 
.A(n_1912),
.B(n_1521),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2041),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_2005),
.B(n_2006),
.Y(n_2189)
);

INVx2_ASAP7_75t_SL g2190 ( 
.A(n_1940),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2063),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1967),
.Y(n_2192)
);

BUFx3_ASAP7_75t_L g2193 ( 
.A(n_1968),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2063),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2066),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_1916),
.B(n_1150),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2066),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2075),
.Y(n_2198)
);

CKINVDCx20_ASAP7_75t_R g2199 ( 
.A(n_1973),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_1919),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2075),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2089),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2089),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_2091),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1971),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1985),
.Y(n_2206)
);

BUFx6f_ASAP7_75t_L g2207 ( 
.A(n_2091),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2033),
.B(n_1092),
.Y(n_2208)
);

OR2x6_ASAP7_75t_L g2209 ( 
.A(n_2096),
.B(n_1275),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1991),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2098),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2098),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1954),
.B(n_1098),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2102),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2102),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2118),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2118),
.Y(n_2217)
);

BUFx6f_ASAP7_75t_L g2218 ( 
.A(n_2130),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_1937),
.Y(n_2219)
);

INVx3_ASAP7_75t_L g2220 ( 
.A(n_2130),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2002),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2132),
.Y(n_2222)
);

INVx4_ASAP7_75t_L g2223 ( 
.A(n_1957),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2132),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_SL g2225 ( 
.A(n_1956),
.B(n_1101),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2002),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2060),
.B(n_1105),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1949),
.B(n_1109),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_1937),
.B(n_1113),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2139),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2139),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2113),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2010),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2031),
.Y(n_2234)
);

OR2x6_ASAP7_75t_L g2235 ( 
.A(n_1906),
.B(n_1216),
.Y(n_2235)
);

INVx2_ASAP7_75t_SL g2236 ( 
.A(n_2076),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2047),
.Y(n_2237)
);

BUFx10_ASAP7_75t_L g2238 ( 
.A(n_2081),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2108),
.B(n_1114),
.Y(n_2239)
);

OAI22xp5_ASAP7_75t_SL g2240 ( 
.A1(n_1934),
.A2(n_1531),
.B1(n_1584),
.B2(n_1524),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2050),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_2030),
.B(n_1115),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_1995),
.B(n_1117),
.Y(n_2243)
);

NAND2xp33_ASAP7_75t_SL g2244 ( 
.A(n_1905),
.B(n_1629),
.Y(n_2244)
);

INVx3_ASAP7_75t_L g2245 ( 
.A(n_1943),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_1943),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1953),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1953),
.Y(n_2248)
);

NAND2xp33_ASAP7_75t_L g2249 ( 
.A(n_2032),
.B(n_1285),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1987),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1964),
.B(n_1196),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2051),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2059),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2156),
.B(n_1118),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_2034),
.B(n_1121),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2077),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2084),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_2013),
.B(n_1129),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1987),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_1992),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1992),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_1999),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1999),
.Y(n_2263)
);

NOR2xp33_ASAP7_75t_L g2264 ( 
.A(n_2061),
.B(n_1123),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_L g2265 ( 
.A(n_2083),
.B(n_1127),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2105),
.B(n_1136),
.Y(n_2266)
);

BUFx10_ASAP7_75t_L g2267 ( 
.A(n_2123),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2112),
.B(n_1140),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2086),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1945),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_1920),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_2025),
.B(n_1141),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2088),
.Y(n_2273)
);

AND3x2_ASAP7_75t_L g2274 ( 
.A(n_2018),
.B(n_2045),
.C(n_1930),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1946),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_2048),
.B(n_1143),
.Y(n_2276)
);

NAND2xp33_ASAP7_75t_L g2277 ( 
.A(n_2114),
.B(n_1285),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2093),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2056),
.B(n_1144),
.Y(n_2279)
);

INVxp67_ASAP7_75t_SL g2280 ( 
.A(n_1982),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2122),
.B(n_1153),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1970),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1976),
.Y(n_2283)
);

AOI21x1_ASAP7_75t_L g2284 ( 
.A1(n_1959),
.A2(n_1374),
.B(n_1363),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1983),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2100),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1920),
.Y(n_2287)
);

BUFx10_ASAP7_75t_L g2288 ( 
.A(n_2169),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1986),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_L g2290 ( 
.A(n_2125),
.B(n_1132),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1994),
.Y(n_2291)
);

NAND2xp33_ASAP7_75t_L g2292 ( 
.A(n_2129),
.B(n_1285),
.Y(n_2292)
);

BUFx10_ASAP7_75t_L g2293 ( 
.A(n_1900),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1996),
.Y(n_2294)
);

HB1xp67_ASAP7_75t_L g2295 ( 
.A(n_1922),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_2017),
.B(n_1157),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_2087),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1902),
.B(n_1196),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2016),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2036),
.B(n_1160),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2106),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2163),
.B(n_1165),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2119),
.B(n_1169),
.Y(n_2303)
);

OR2x6_ASAP7_75t_L g2304 ( 
.A(n_2004),
.B(n_1977),
.Y(n_2304)
);

HB1xp67_ASAP7_75t_L g2305 ( 
.A(n_1933),
.Y(n_2305)
);

INVx2_ASAP7_75t_SL g2306 ( 
.A(n_2092),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2107),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2127),
.Y(n_2308)
);

INVx3_ASAP7_75t_L g2309 ( 
.A(n_1931),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2136),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2146),
.Y(n_2311)
);

CKINVDCx6p67_ASAP7_75t_R g2312 ( 
.A(n_2080),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2147),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2009),
.B(n_1176),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2057),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2149),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1915),
.B(n_1184),
.Y(n_2317)
);

INVx3_ASAP7_75t_L g2318 ( 
.A(n_1931),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1901),
.B(n_1197),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2012),
.B(n_1203),
.Y(n_2320)
);

AOI21x1_ASAP7_75t_L g2321 ( 
.A1(n_1965),
.A2(n_1975),
.B(n_1969),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2154),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2068),
.Y(n_2323)
);

INVx3_ASAP7_75t_L g2324 ( 
.A(n_2103),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2109),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_1923),
.B(n_1134),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1951),
.B(n_1204),
.Y(n_2327)
);

INVx3_ASAP7_75t_L g2328 ( 
.A(n_2111),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_1926),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1929),
.Y(n_2330)
);

INVx2_ASAP7_75t_SL g2331 ( 
.A(n_2128),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_1917),
.B(n_1139),
.Y(n_2332)
);

AOI21x1_ASAP7_75t_L g2333 ( 
.A1(n_1978),
.A2(n_1383),
.B(n_1379),
.Y(n_2333)
);

INVx2_ASAP7_75t_SL g2334 ( 
.A(n_2151),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1935),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_1925),
.B(n_1145),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2115),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_1938),
.Y(n_2338)
);

NAND3xp33_ASAP7_75t_L g2339 ( 
.A(n_1948),
.B(n_1155),
.C(n_1151),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_1939),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2003),
.B(n_1972),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2126),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1942),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_2134),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2140),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2142),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1903),
.Y(n_2347)
);

INVx1_ASAP7_75t_SL g2348 ( 
.A(n_1908),
.Y(n_2348)
);

INVx8_ASAP7_75t_L g2349 ( 
.A(n_2001),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_1904),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2155),
.B(n_2162),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_2159),
.Y(n_2352)
);

BUFx2_ASAP7_75t_L g2353 ( 
.A(n_2023),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1909),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1911),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_1918),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_2043),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_1898),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2161),
.Y(n_2359)
);

AO21x2_ASAP7_75t_L g2360 ( 
.A1(n_2011),
.A2(n_1393),
.B(n_1389),
.Y(n_2360)
);

AO21x2_ASAP7_75t_L g2361 ( 
.A1(n_1988),
.A2(n_1419),
.B(n_1396),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2019),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2020),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_1950),
.B(n_1161),
.Y(n_2364)
);

BUFx6f_ASAP7_75t_L g2365 ( 
.A(n_2054),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2021),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_1941),
.B(n_1207),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_1952),
.B(n_1208),
.Y(n_2368)
);

INVx3_ASAP7_75t_L g2369 ( 
.A(n_2164),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1990),
.B(n_1210),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2035),
.Y(n_2371)
);

INVxp33_ASAP7_75t_SL g2372 ( 
.A(n_1961),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2039),
.Y(n_2373)
);

NAND2xp33_ASAP7_75t_SL g2374 ( 
.A(n_1914),
.B(n_1660),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2042),
.Y(n_2375)
);

BUFx3_ASAP7_75t_L g2376 ( 
.A(n_1910),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2053),
.Y(n_2377)
);

NAND3xp33_ASAP7_75t_L g2378 ( 
.A(n_1997),
.B(n_1175),
.C(n_1162),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2062),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_SL g2380 ( 
.A(n_1928),
.B(n_1663),
.Y(n_2380)
);

INVx8_ASAP7_75t_L g2381 ( 
.A(n_2085),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1963),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2065),
.Y(n_2383)
);

INVx3_ASAP7_75t_L g2384 ( 
.A(n_1944),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1979),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1984),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_1936),
.B(n_1252),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2072),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2074),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2079),
.Y(n_2390)
);

INVxp67_ASAP7_75t_SL g2391 ( 
.A(n_1980),
.Y(n_2391)
);

INVxp67_ASAP7_75t_SL g2392 ( 
.A(n_1981),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2097),
.Y(n_2393)
);

HB1xp67_ASAP7_75t_L g2394 ( 
.A(n_2038),
.Y(n_2394)
);

AND3x2_ASAP7_75t_L g2395 ( 
.A(n_2040),
.B(n_1550),
.C(n_1548),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2052),
.A2(n_1298),
.B1(n_1371),
.B2(n_1280),
.Y(n_2396)
);

NAND2xp33_ASAP7_75t_L g2397 ( 
.A(n_2000),
.B(n_1403),
.Y(n_2397)
);

NOR2xp33_ASAP7_75t_L g2398 ( 
.A(n_2082),
.B(n_1178),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_2022),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2058),
.B(n_1211),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2099),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2116),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2117),
.Y(n_2403)
);

AOI21x1_ASAP7_75t_L g2404 ( 
.A1(n_1955),
.A2(n_1444),
.B(n_1442),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2121),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2133),
.Y(n_2406)
);

AND3x2_ASAP7_75t_L g2407 ( 
.A(n_2070),
.B(n_1677),
.C(n_1580),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2110),
.B(n_1252),
.Y(n_2408)
);

NAND2xp33_ASAP7_75t_SL g2409 ( 
.A(n_2168),
.B(n_1664),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2135),
.Y(n_2410)
);

AND2x2_ASAP7_75t_L g2411 ( 
.A(n_2174),
.B(n_2007),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2196),
.B(n_2184),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2173),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_L g2414 ( 
.A(n_2332),
.B(n_2095),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_2199),
.Y(n_2415)
);

XOR2xp5_ASAP7_75t_L g2416 ( 
.A(n_2372),
.B(n_2069),
.Y(n_2416)
);

NAND2xp33_ASAP7_75t_SL g2417 ( 
.A(n_2251),
.B(n_2008),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2181),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2193),
.B(n_2175),
.Y(n_2419)
);

XNOR2xp5_ASAP7_75t_L g2420 ( 
.A(n_2348),
.B(n_2150),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2351),
.B(n_2037),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2236),
.B(n_2055),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2192),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2297),
.B(n_2073),
.Y(n_2424)
);

AOI21x1_ASAP7_75t_L g2425 ( 
.A1(n_2404),
.A2(n_2157),
.B(n_2015),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2391),
.B(n_2392),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2336),
.B(n_2165),
.Y(n_2427)
);

INVx1_ASAP7_75t_SL g2428 ( 
.A(n_2189),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2205),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2206),
.Y(n_2430)
);

XNOR2xp5_ASAP7_75t_L g2431 ( 
.A(n_2274),
.B(n_2101),
.Y(n_2431)
);

INVx2_ASAP7_75t_SL g2432 ( 
.A(n_2306),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2331),
.B(n_2094),
.Y(n_2433)
);

AND2x4_ASAP7_75t_L g2434 ( 
.A(n_2186),
.B(n_2120),
.Y(n_2434)
);

XOR2xp5_ASAP7_75t_L g2435 ( 
.A(n_2353),
.B(n_1993),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2210),
.Y(n_2436)
);

INVxp67_ASAP7_75t_SL g2437 ( 
.A(n_2246),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2270),
.Y(n_2438)
);

CKINVDCx5p33_ASAP7_75t_R g2439 ( 
.A(n_2238),
.Y(n_2439)
);

CKINVDCx20_ASAP7_75t_R g2440 ( 
.A(n_2312),
.Y(n_2440)
);

XNOR2x2_ASAP7_75t_L g2441 ( 
.A(n_2396),
.B(n_1947),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2334),
.B(n_2144),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2242),
.B(n_1958),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2233),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2234),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_2255),
.B(n_1989),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2237),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2241),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2252),
.Y(n_2449)
);

XOR2xp5_ASAP7_75t_L g2450 ( 
.A(n_2240),
.B(n_1899),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2253),
.Y(n_2451)
);

XOR2xp5_ASAP7_75t_L g2452 ( 
.A(n_2295),
.B(n_1924),
.Y(n_2452)
);

XNOR2xp5_ASAP7_75t_L g2453 ( 
.A(n_2190),
.B(n_2028),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2256),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2264),
.B(n_2104),
.Y(n_2455)
);

INVx4_ASAP7_75t_SL g2456 ( 
.A(n_2209),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2257),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2269),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2387),
.B(n_2067),
.Y(n_2459)
);

INVxp33_ASAP7_75t_L g2460 ( 
.A(n_2305),
.Y(n_2460)
);

AND2x4_ASAP7_75t_L g2461 ( 
.A(n_2200),
.B(n_2137),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2273),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2298),
.B(n_1998),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2278),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2286),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2301),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2408),
.B(n_2124),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2307),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2308),
.Y(n_2469)
);

AND2x4_ASAP7_75t_L g2470 ( 
.A(n_2376),
.B(n_2138),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2310),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2265),
.B(n_1457),
.Y(n_2472)
);

NAND2xp33_ASAP7_75t_R g2473 ( 
.A(n_2341),
.B(n_1223),
.Y(n_2473)
);

CKINVDCx5p33_ASAP7_75t_R g2474 ( 
.A(n_2267),
.Y(n_2474)
);

BUFx6f_ASAP7_75t_L g2475 ( 
.A(n_2180),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2311),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2313),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2280),
.B(n_2141),
.Y(n_2478)
);

NAND2x1p5_ASAP7_75t_L g2479 ( 
.A(n_2223),
.B(n_2143),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2316),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_SL g2481 ( 
.A(n_2288),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2322),
.Y(n_2482)
);

CKINVDCx20_ASAP7_75t_R g2483 ( 
.A(n_2349),
.Y(n_2483)
);

CKINVDCx20_ASAP7_75t_R g2484 ( 
.A(n_2349),
.Y(n_2484)
);

NOR2xp33_ASAP7_75t_L g2485 ( 
.A(n_2290),
.B(n_2044),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_SL g2486 ( 
.A(n_2380),
.B(n_2046),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2329),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2275),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_2180),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2282),
.Y(n_2490)
);

XOR2xp5_ASAP7_75t_L g2491 ( 
.A(n_2394),
.B(n_2078),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2179),
.B(n_2131),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2326),
.B(n_2145),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_2381),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2283),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2330),
.Y(n_2496)
);

AND2x2_ASAP7_75t_L g2497 ( 
.A(n_2399),
.B(n_2148),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2285),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2289),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2291),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_2204),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2294),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2388),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2390),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2246),
.B(n_2152),
.Y(n_2505)
);

BUFx6f_ASAP7_75t_L g2506 ( 
.A(n_2204),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_2260),
.B(n_2384),
.Y(n_2507)
);

INVx1_ASAP7_75t_SL g2508 ( 
.A(n_2409),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2402),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2410),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2358),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2266),
.B(n_1458),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2362),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_2381),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2363),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2366),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2371),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_2208),
.B(n_1416),
.Y(n_2518)
);

BUFx2_ASAP7_75t_R g2519 ( 
.A(n_2228),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2268),
.B(n_1477),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2373),
.Y(n_2521)
);

INVx2_ASAP7_75t_SL g2522 ( 
.A(n_2170),
.Y(n_2522)
);

BUFx5_ASAP7_75t_L g2523 ( 
.A(n_2382),
.Y(n_2523)
);

INVx2_ASAP7_75t_SL g2524 ( 
.A(n_2172),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2335),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2375),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2377),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2227),
.B(n_1553),
.Y(n_2528)
);

INVxp67_ASAP7_75t_SL g2529 ( 
.A(n_2260),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2178),
.B(n_1228),
.Y(n_2530)
);

XOR2xp5_ASAP7_75t_L g2531 ( 
.A(n_2378),
.B(n_1676),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2379),
.Y(n_2532)
);

BUFx2_ASAP7_75t_L g2533 ( 
.A(n_2235),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2383),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2389),
.Y(n_2535)
);

XOR2xp5_ASAP7_75t_L g2536 ( 
.A(n_2339),
.B(n_1681),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2393),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2401),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2403),
.Y(n_2539)
);

INVx3_ASAP7_75t_R g2540 ( 
.A(n_2405),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2219),
.B(n_2153),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_L g2542 ( 
.A(n_2239),
.B(n_2254),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2324),
.B(n_2158),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2281),
.B(n_1480),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2406),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2338),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2340),
.Y(n_2547)
);

OAI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_2317),
.A2(n_2029),
.B(n_1484),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2343),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2302),
.B(n_1569),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2347),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_2370),
.B(n_2314),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2350),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2354),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_2304),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2328),
.B(n_2160),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2355),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2356),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2299),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2315),
.Y(n_2560)
);

INVx3_ASAP7_75t_R g2561 ( 
.A(n_2177),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2323),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2325),
.Y(n_2563)
);

AND2x2_ASAP7_75t_SL g2564 ( 
.A(n_2364),
.B(n_1714),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2337),
.Y(n_2565)
);

NAND2x1p5_ASAP7_75t_L g2566 ( 
.A(n_2245),
.B(n_2166),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2188),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_SL g2568 ( 
.A(n_2209),
.B(n_2027),
.Y(n_2568)
);

XOR2xp5_ASAP7_75t_L g2569 ( 
.A(n_2400),
.B(n_1725),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2342),
.Y(n_2570)
);

INVxp33_ASAP7_75t_L g2571 ( 
.A(n_2176),
.Y(n_2571)
);

INVxp67_ASAP7_75t_SL g2572 ( 
.A(n_2207),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2345),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2346),
.Y(n_2574)
);

AOI21xp5_ASAP7_75t_L g2575 ( 
.A1(n_2182),
.A2(n_1486),
.B(n_1483),
.Y(n_2575)
);

AOI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2185),
.A2(n_1491),
.B(n_1487),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2448),
.Y(n_2577)
);

OAI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_2443),
.A2(n_2319),
.B(n_2327),
.Y(n_2578)
);

INVx3_ASAP7_75t_L g2579 ( 
.A(n_2501),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2413),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2542),
.B(n_2398),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_L g2582 ( 
.A(n_2455),
.B(n_2183),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2426),
.B(n_2360),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2564),
.B(n_2232),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2414),
.B(n_2321),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2427),
.B(n_2225),
.Y(n_2586)
);

BUFx8_ASAP7_75t_L g2587 ( 
.A(n_2481),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_2412),
.B(n_2385),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2418),
.Y(n_2589)
);

BUFx5_ASAP7_75t_L g2590 ( 
.A(n_2423),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2419),
.B(n_2344),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2518),
.B(n_2213),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2428),
.B(n_2411),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2446),
.B(n_2187),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2449),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_2528),
.B(n_2386),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2475),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2550),
.B(n_2552),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2429),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2472),
.B(n_2243),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2467),
.B(n_2304),
.Y(n_2601)
);

INVx3_ASAP7_75t_L g2602 ( 
.A(n_2501),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2485),
.A2(n_2374),
.B1(n_2244),
.B2(n_2361),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2469),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_2415),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2421),
.B(n_2293),
.Y(n_2606)
);

HB1xp67_ASAP7_75t_L g2607 ( 
.A(n_2475),
.Y(n_2607)
);

AOI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2492),
.A2(n_2320),
.B1(n_2258),
.B2(n_2276),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_2571),
.B(n_2367),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2430),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_2463),
.B(n_2352),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2487),
.Y(n_2612)
);

BUFx6f_ASAP7_75t_L g2613 ( 
.A(n_2489),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2493),
.B(n_2272),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2486),
.B(n_2369),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2496),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2523),
.B(n_2279),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2523),
.B(n_2368),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2436),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_SL g2620 ( 
.A(n_2459),
.B(n_2271),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2432),
.B(n_2271),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2523),
.B(n_2296),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2438),
.Y(n_2623)
);

INVx2_ASAP7_75t_SL g2624 ( 
.A(n_2506),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_2417),
.B(n_2262),
.Y(n_2625)
);

NOR2xp33_ASAP7_75t_L g2626 ( 
.A(n_2460),
.B(n_2300),
.Y(n_2626)
);

AOI21xp5_ASAP7_75t_L g2627 ( 
.A1(n_2548),
.A2(n_2520),
.B(n_2512),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2523),
.B(n_2544),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2478),
.B(n_2303),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2503),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2525),
.Y(n_2631)
);

BUFx6f_ASAP7_75t_L g2632 ( 
.A(n_2489),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2504),
.B(n_2509),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2510),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2444),
.Y(n_2635)
);

INVx3_ASAP7_75t_L g2636 ( 
.A(n_2506),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2445),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2447),
.Y(n_2638)
);

AOI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2441),
.A2(n_2365),
.B1(n_2357),
.B2(n_1541),
.Y(n_2639)
);

O2A1O1Ixp5_ASAP7_75t_L g2640 ( 
.A1(n_2530),
.A2(n_2284),
.B(n_2333),
.C(n_2229),
.Y(n_2640)
);

INVx3_ASAP7_75t_L g2641 ( 
.A(n_2461),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_2508),
.B(n_2422),
.Y(n_2642)
);

OAI21xp5_ASAP7_75t_L g2643 ( 
.A1(n_2425),
.A2(n_2277),
.B(n_2249),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2451),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2454),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2457),
.B(n_2191),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2458),
.B(n_2194),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_L g2648 ( 
.A(n_2569),
.B(n_2235),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2462),
.B(n_2464),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2465),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2466),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_SL g2652 ( 
.A(n_2424),
.B(n_2207),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2468),
.Y(n_2653)
);

INVxp67_ASAP7_75t_L g2654 ( 
.A(n_2433),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_2452),
.B(n_2247),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2471),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2476),
.B(n_2195),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2477),
.B(n_2197),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2480),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2482),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2546),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2536),
.B(n_2453),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2547),
.B(n_2198),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2549),
.B(n_2201),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2551),
.B(n_2202),
.Y(n_2665)
);

NOR2xp67_ASAP7_75t_SL g2666 ( 
.A(n_2439),
.B(n_2474),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2553),
.B(n_2203),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2554),
.B(n_2211),
.Y(n_2668)
);

AOI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2557),
.A2(n_2365),
.B(n_2357),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2558),
.B(n_2212),
.Y(n_2670)
);

INVxp67_ASAP7_75t_SL g2671 ( 
.A(n_2507),
.Y(n_2671)
);

NOR3xp33_ASAP7_75t_L g2672 ( 
.A(n_2533),
.B(n_2250),
.C(n_2248),
.Y(n_2672)
);

AOI22xp33_ASAP7_75t_L g2673 ( 
.A1(n_2575),
.A2(n_1549),
.B1(n_1578),
.B2(n_1565),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2488),
.B(n_2214),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2490),
.B(n_2215),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2598),
.B(n_2495),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2613),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2580),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2581),
.B(n_2498),
.Y(n_2679)
);

AOI22xp33_ASAP7_75t_L g2680 ( 
.A1(n_2582),
.A2(n_2499),
.B1(n_2502),
.B2(n_2500),
.Y(n_2680)
);

BUFx2_ASAP7_75t_L g2681 ( 
.A(n_2593),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_L g2682 ( 
.A(n_2613),
.Y(n_2682)
);

HB1xp67_ASAP7_75t_L g2683 ( 
.A(n_2632),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2577),
.Y(n_2684)
);

AND2x4_ASAP7_75t_L g2685 ( 
.A(n_2591),
.B(n_2470),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2589),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2671),
.B(n_2434),
.Y(n_2687)
);

BUFx3_ASAP7_75t_L g2688 ( 
.A(n_2632),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2595),
.Y(n_2689)
);

BUFx3_ASAP7_75t_L g2690 ( 
.A(n_2579),
.Y(n_2690)
);

BUFx6f_ASAP7_75t_L g2691 ( 
.A(n_2624),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2599),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2610),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2619),
.Y(n_2694)
);

INVx3_ASAP7_75t_L g2695 ( 
.A(n_2602),
.Y(n_2695)
);

INVx2_ASAP7_75t_SL g2696 ( 
.A(n_2597),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2623),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2606),
.B(n_2437),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2630),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2634),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_2605),
.Y(n_2701)
);

NAND2x1p5_ASAP7_75t_L g2702 ( 
.A(n_2636),
.B(n_2442),
.Y(n_2702)
);

HB1xp67_ASAP7_75t_L g2703 ( 
.A(n_2607),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2586),
.B(n_2511),
.Y(n_2704)
);

BUFx2_ASAP7_75t_L g2705 ( 
.A(n_2601),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2633),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2649),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_2641),
.B(n_2529),
.Y(n_2708)
);

NOR3xp33_ASAP7_75t_SL g2709 ( 
.A(n_2648),
.B(n_2555),
.C(n_2473),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2637),
.Y(n_2710)
);

A2O1A1Ixp33_ASAP7_75t_L g2711 ( 
.A1(n_2594),
.A2(n_2576),
.B(n_2560),
.C(n_2562),
.Y(n_2711)
);

AOI22xp5_ASAP7_75t_L g2712 ( 
.A1(n_2609),
.A2(n_2497),
.B1(n_2515),
.B2(n_2513),
.Y(n_2712)
);

HB1xp67_ASAP7_75t_L g2713 ( 
.A(n_2654),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2672),
.B(n_2456),
.Y(n_2714)
);

CKINVDCx20_ASAP7_75t_R g2715 ( 
.A(n_2587),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2614),
.B(n_2531),
.Y(n_2716)
);

INVx5_ASAP7_75t_L g2717 ( 
.A(n_2635),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2638),
.Y(n_2718)
);

INVx3_ASAP7_75t_L g2719 ( 
.A(n_2661),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2604),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2644),
.Y(n_2721)
);

NOR2xp33_ASAP7_75t_L g2722 ( 
.A(n_2592),
.B(n_2420),
.Y(n_2722)
);

INVxp67_ASAP7_75t_SL g2723 ( 
.A(n_2590),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2600),
.B(n_2516),
.Y(n_2724)
);

BUFx3_ASAP7_75t_L g2725 ( 
.A(n_2655),
.Y(n_2725)
);

AOI22x1_ASAP7_75t_L g2726 ( 
.A1(n_2627),
.A2(n_2578),
.B1(n_2643),
.B2(n_2669),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2629),
.B(n_2517),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2612),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2603),
.B(n_2521),
.Y(n_2729)
);

NAND3xp33_ASAP7_75t_SL g2730 ( 
.A(n_2608),
.B(n_2568),
.C(n_2450),
.Y(n_2730)
);

HB1xp67_ASAP7_75t_L g2731 ( 
.A(n_2645),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2616),
.Y(n_2732)
);

AND2x4_ASAP7_75t_L g2733 ( 
.A(n_2652),
.B(n_2456),
.Y(n_2733)
);

O2A1O1Ixp5_ASAP7_75t_L g2734 ( 
.A1(n_2585),
.A2(n_2527),
.B(n_2532),
.C(n_2526),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2631),
.Y(n_2735)
);

NAND2x1p5_ASAP7_75t_L g2736 ( 
.A(n_2666),
.B(n_2218),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2590),
.B(n_2534),
.Y(n_2737)
);

AOI221xp5_ASAP7_75t_L g2738 ( 
.A1(n_2662),
.A2(n_2491),
.B1(n_1766),
.B2(n_1760),
.C(n_1739),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2621),
.B(n_2572),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2590),
.B(n_2535),
.Y(n_2740)
);

INVx2_ASAP7_75t_SL g2741 ( 
.A(n_2620),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2650),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2651),
.A2(n_2538),
.B1(n_2539),
.B2(n_2537),
.Y(n_2743)
);

BUFx6f_ASAP7_75t_L g2744 ( 
.A(n_2642),
.Y(n_2744)
);

BUFx2_ASAP7_75t_L g2745 ( 
.A(n_2653),
.Y(n_2745)
);

NAND2xp33_ASAP7_75t_L g2746 ( 
.A(n_2590),
.B(n_2494),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2656),
.A2(n_2545),
.B1(n_2563),
.B2(n_2559),
.Y(n_2747)
);

INVx3_ASAP7_75t_L g2748 ( 
.A(n_2659),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2660),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2674),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2596),
.B(n_2543),
.Y(n_2751)
);

AND2x6_ASAP7_75t_L g2752 ( 
.A(n_2617),
.B(n_2565),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2588),
.B(n_2570),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2675),
.Y(n_2754)
);

BUFx6f_ASAP7_75t_L g2755 ( 
.A(n_2615),
.Y(n_2755)
);

AND2x4_ASAP7_75t_L g2756 ( 
.A(n_2611),
.B(n_2573),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_R g2757 ( 
.A(n_2626),
.B(n_2514),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_2584),
.Y(n_2758)
);

NAND2xp33_ASAP7_75t_SL g2759 ( 
.A(n_2618),
.B(n_2540),
.Y(n_2759)
);

INVx4_ASAP7_75t_L g2760 ( 
.A(n_2677),
.Y(n_2760)
);

OAI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2729),
.A2(n_2734),
.B(n_2679),
.Y(n_2761)
);

OA22x2_ASAP7_75t_L g2762 ( 
.A1(n_2758),
.A2(n_2171),
.B1(n_2407),
.B2(n_2395),
.Y(n_2762)
);

OAI21xp33_ASAP7_75t_L g2763 ( 
.A1(n_2738),
.A2(n_2519),
.B(n_1736),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2690),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2678),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2749),
.Y(n_2766)
);

AOI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2726),
.A2(n_2628),
.B(n_2583),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2686),
.Y(n_2768)
);

AOI21xp5_ASAP7_75t_L g2769 ( 
.A1(n_2723),
.A2(n_2622),
.B(n_2704),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2724),
.A2(n_2639),
.B(n_2625),
.Y(n_2770)
);

OA21x2_ASAP7_75t_L g2771 ( 
.A1(n_2737),
.A2(n_2740),
.B(n_2711),
.Y(n_2771)
);

OR2x2_ASAP7_75t_L g2772 ( 
.A(n_2681),
.B(n_2416),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2676),
.A2(n_2640),
.B(n_2665),
.Y(n_2773)
);

BUFx6f_ASAP7_75t_L g2774 ( 
.A(n_2677),
.Y(n_2774)
);

INVx1_ASAP7_75t_SL g2775 ( 
.A(n_2725),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2688),
.Y(n_2776)
);

AOI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2727),
.A2(n_2706),
.B(n_2707),
.Y(n_2777)
);

BUFx12f_ASAP7_75t_L g2778 ( 
.A(n_2701),
.Y(n_2778)
);

AOI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_2746),
.A2(n_2668),
.B(n_2667),
.Y(n_2779)
);

AO31x2_ASAP7_75t_L g2780 ( 
.A1(n_2754),
.A2(n_2718),
.A3(n_2721),
.B(n_2710),
.Y(n_2780)
);

INVx3_ASAP7_75t_L g2781 ( 
.A(n_2717),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2692),
.Y(n_2782)
);

AOI21xp5_ASAP7_75t_L g2783 ( 
.A1(n_2751),
.A2(n_2670),
.B(n_2647),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2722),
.B(n_2556),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2750),
.B(n_2716),
.Y(n_2785)
);

NAND2x1p5_ASAP7_75t_L g2786 ( 
.A(n_2717),
.B(n_2522),
.Y(n_2786)
);

AOI21x1_ASAP7_75t_L g2787 ( 
.A1(n_2693),
.A2(n_2657),
.B(n_2646),
.Y(n_2787)
);

AOI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2680),
.A2(n_2663),
.B(n_2658),
.Y(n_2788)
);

OAI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2712),
.A2(n_2743),
.B(n_2747),
.Y(n_2789)
);

OAI21x1_ASAP7_75t_L g2790 ( 
.A1(n_2748),
.A2(n_2664),
.B(n_2574),
.Y(n_2790)
);

OAI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2694),
.A2(n_2479),
.B1(n_2567),
.B2(n_2524),
.Y(n_2791)
);

NAND3xp33_ASAP7_75t_L g2792 ( 
.A(n_2709),
.B(n_2071),
.C(n_2064),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2755),
.B(n_2505),
.Y(n_2793)
);

AO21x1_ASAP7_75t_L g2794 ( 
.A1(n_2759),
.A2(n_2756),
.B(n_2699),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2697),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2700),
.Y(n_2796)
);

OR2x2_ASAP7_75t_L g2797 ( 
.A(n_2705),
.B(n_2435),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2731),
.Y(n_2798)
);

OAI21x1_ASAP7_75t_L g2799 ( 
.A1(n_2684),
.A2(n_2566),
.B(n_2217),
.Y(n_2799)
);

CKINVDCx20_ASAP7_75t_R g2800 ( 
.A(n_2715),
.Y(n_2800)
);

OAI21xp5_ASAP7_75t_L g2801 ( 
.A1(n_2689),
.A2(n_2673),
.B(n_2541),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2720),
.Y(n_2802)
);

OAI21x1_ASAP7_75t_L g2803 ( 
.A1(n_2728),
.A2(n_2222),
.B(n_2216),
.Y(n_2803)
);

O2A1O1Ixp5_ASAP7_75t_L g2804 ( 
.A1(n_2753),
.A2(n_2224),
.B(n_2231),
.C(n_2230),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2732),
.Y(n_2805)
);

AO21x1_ASAP7_75t_L g2806 ( 
.A1(n_2735),
.A2(n_2292),
.B(n_1597),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2755),
.B(n_2719),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2742),
.B(n_2359),
.Y(n_2808)
);

OAI21x1_ASAP7_75t_L g2809 ( 
.A1(n_2702),
.A2(n_2261),
.B(n_2259),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2698),
.B(n_2431),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2730),
.B(n_2483),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2682),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2745),
.B(n_2741),
.Y(n_2813)
);

AND2x2_ASAP7_75t_SL g2814 ( 
.A(n_2714),
.B(n_2484),
.Y(n_2814)
);

OAI21x1_ASAP7_75t_L g2815 ( 
.A1(n_2736),
.A2(n_2263),
.B(n_2226),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2713),
.B(n_2090),
.Y(n_2816)
);

AOI21x1_ASAP7_75t_L g2817 ( 
.A1(n_2739),
.A2(n_2221),
.B(n_2167),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2687),
.A2(n_2397),
.B(n_1407),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2744),
.B(n_2220),
.Y(n_2819)
);

BUFx3_ASAP7_75t_L g2820 ( 
.A(n_2682),
.Y(n_2820)
);

OAI21xp5_ASAP7_75t_L g2821 ( 
.A1(n_2752),
.A2(n_1604),
.B(n_1593),
.Y(n_2821)
);

AOI21xp33_ASAP7_75t_L g2822 ( 
.A1(n_2744),
.A2(n_1752),
.B(n_1734),
.Y(n_2822)
);

BUFx2_ASAP7_75t_L g2823 ( 
.A(n_2703),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2708),
.B(n_2287),
.Y(n_2824)
);

OAI21x1_ASAP7_75t_L g2825 ( 
.A1(n_2790),
.A2(n_2318),
.B(n_2309),
.Y(n_2825)
);

INVx4_ASAP7_75t_L g2826 ( 
.A(n_2774),
.Y(n_2826)
);

INVx1_ASAP7_75t_SL g2827 ( 
.A(n_2775),
.Y(n_2827)
);

BUFx3_ASAP7_75t_L g2828 ( 
.A(n_2812),
.Y(n_2828)
);

OAI21x1_ASAP7_75t_L g2829 ( 
.A1(n_2767),
.A2(n_1619),
.B(n_1616),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2764),
.B(n_2685),
.Y(n_2830)
);

OAI21x1_ASAP7_75t_L g2831 ( 
.A1(n_2803),
.A2(n_1675),
.B(n_1634),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2777),
.B(n_2757),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2784),
.B(n_2696),
.Y(n_2833)
);

A2O1A1Ixp33_ASAP7_75t_L g2834 ( 
.A1(n_2789),
.A2(n_2733),
.B(n_1684),
.C(n_1701),
.Y(n_2834)
);

OAI22xp5_ASAP7_75t_L g2835 ( 
.A1(n_2785),
.A2(n_2763),
.B1(n_2813),
.B2(n_2793),
.Y(n_2835)
);

OAI21x1_ASAP7_75t_L g2836 ( 
.A1(n_2773),
.A2(n_1705),
.B(n_1680),
.Y(n_2836)
);

AO31x2_ASAP7_75t_L g2837 ( 
.A1(n_2806),
.A2(n_2794),
.A3(n_2769),
.B(n_2770),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2798),
.B(n_2683),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2761),
.A2(n_2752),
.B(n_1407),
.Y(n_2839)
);

OAI21x1_ASAP7_75t_L g2840 ( 
.A1(n_2799),
.A2(n_1712),
.B(n_1711),
.Y(n_2840)
);

OAI21x1_ASAP7_75t_L g2841 ( 
.A1(n_2787),
.A2(n_1719),
.B(n_1713),
.Y(n_2841)
);

AOI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2779),
.A2(n_2752),
.B(n_1407),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2772),
.B(n_2695),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2768),
.Y(n_2844)
);

AO31x2_ASAP7_75t_L g2845 ( 
.A1(n_2783),
.A2(n_1740),
.A3(n_1750),
.B(n_1724),
.Y(n_2845)
);

AO31x2_ASAP7_75t_L g2846 ( 
.A1(n_2788),
.A2(n_2818),
.A3(n_2791),
.B(n_2782),
.Y(n_2846)
);

OAI21x1_ASAP7_75t_L g2847 ( 
.A1(n_2771),
.A2(n_1220),
.B(n_1217),
.Y(n_2847)
);

OAI21x1_ASAP7_75t_L g2848 ( 
.A1(n_2817),
.A2(n_2815),
.B(n_2809),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_2778),
.Y(n_2849)
);

BUFx3_ASAP7_75t_L g2850 ( 
.A(n_2820),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2823),
.Y(n_2851)
);

AOI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2801),
.A2(n_2821),
.B(n_2796),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2766),
.B(n_2691),
.Y(n_2853)
);

AO21x1_ASAP7_75t_L g2854 ( 
.A1(n_2765),
.A2(n_1226),
.B(n_1222),
.Y(n_2854)
);

INVxp67_ASAP7_75t_SL g2855 ( 
.A(n_2795),
.Y(n_2855)
);

OAI21x1_ASAP7_75t_L g2856 ( 
.A1(n_2804),
.A2(n_1239),
.B(n_1230),
.Y(n_2856)
);

INVx3_ASAP7_75t_L g2857 ( 
.A(n_2760),
.Y(n_2857)
);

O2A1O1Ixp5_ASAP7_75t_L g2858 ( 
.A1(n_2811),
.A2(n_1254),
.B(n_1263),
.C(n_1250),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2807),
.B(n_2691),
.Y(n_2859)
);

AOI21xp5_ASAP7_75t_L g2860 ( 
.A1(n_2802),
.A2(n_1478),
.B(n_1403),
.Y(n_2860)
);

AOI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2805),
.A2(n_1478),
.B(n_1403),
.Y(n_2861)
);

OAI21xp5_ASAP7_75t_L g2862 ( 
.A1(n_2808),
.A2(n_2824),
.B(n_2819),
.Y(n_2862)
);

AO31x2_ASAP7_75t_L g2863 ( 
.A1(n_2780),
.A2(n_1773),
.A3(n_1753),
.B(n_1273),
.Y(n_2863)
);

AO31x2_ASAP7_75t_L g2864 ( 
.A1(n_2780),
.A2(n_1276),
.A3(n_1279),
.B(n_1272),
.Y(n_2864)
);

OAI21x1_ASAP7_75t_L g2865 ( 
.A1(n_2786),
.A2(n_1286),
.B(n_1282),
.Y(n_2865)
);

OAI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2797),
.A2(n_2440),
.B1(n_2218),
.B2(n_1183),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2781),
.Y(n_2867)
);

AO21x2_ASAP7_75t_L g2868 ( 
.A1(n_2792),
.A2(n_1303),
.B(n_1293),
.Y(n_2868)
);

OAI21xp33_ASAP7_75t_SL g2869 ( 
.A1(n_2762),
.A2(n_1318),
.B(n_1312),
.Y(n_2869)
);

A2O1A1Ixp33_ASAP7_75t_L g2870 ( 
.A1(n_2822),
.A2(n_1339),
.B(n_1340),
.C(n_1326),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2774),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2776),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2814),
.Y(n_2873)
);

INVx3_ASAP7_75t_SL g2874 ( 
.A(n_2800),
.Y(n_2874)
);

AO21x2_ASAP7_75t_L g2875 ( 
.A1(n_2810),
.A2(n_1352),
.B(n_1350),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2816),
.Y(n_2876)
);

A2O1A1Ixp33_ASAP7_75t_L g2877 ( 
.A1(n_2789),
.A2(n_1366),
.B(n_1369),
.C(n_1358),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2768),
.Y(n_2878)
);

OAI21x1_ASAP7_75t_L g2879 ( 
.A1(n_2790),
.A2(n_1380),
.B(n_1377),
.Y(n_2879)
);

OAI21xp5_ASAP7_75t_L g2880 ( 
.A1(n_2770),
.A2(n_1384),
.B(n_1381),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2768),
.Y(n_2881)
);

AO31x2_ASAP7_75t_L g2882 ( 
.A1(n_2767),
.A2(n_1386),
.A3(n_1426),
.B(n_1417),
.Y(n_2882)
);

OAI21x1_ASAP7_75t_L g2883 ( 
.A1(n_2790),
.A2(n_1443),
.B(n_1440),
.Y(n_2883)
);

AO31x2_ASAP7_75t_L g2884 ( 
.A1(n_2767),
.A2(n_1447),
.A3(n_1469),
.B(n_1462),
.Y(n_2884)
);

AOI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2767),
.A2(n_1529),
.B(n_1478),
.Y(n_2885)
);

INVx8_ASAP7_75t_L g2886 ( 
.A(n_2830),
.Y(n_2886)
);

OAI21xp5_ASAP7_75t_L g2887 ( 
.A1(n_2880),
.A2(n_1560),
.B(n_1539),
.Y(n_2887)
);

AOI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_2875),
.A2(n_1186),
.B1(n_1189),
.B2(n_1181),
.Y(n_2888)
);

BUFx4f_ASAP7_75t_SL g2889 ( 
.A(n_2874),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2835),
.B(n_1780),
.Y(n_2890)
);

AOI22xp33_ASAP7_75t_L g2891 ( 
.A1(n_2873),
.A2(n_1283),
.B1(n_1402),
.B2(n_1259),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2844),
.Y(n_2892)
);

INVx4_ASAP7_75t_L g2893 ( 
.A(n_2826),
.Y(n_2893)
);

AOI22xp5_ASAP7_75t_L g2894 ( 
.A1(n_2876),
.A2(n_1205),
.B1(n_1209),
.B2(n_1199),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2878),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2864),
.Y(n_2896)
);

CKINVDCx20_ASAP7_75t_R g2897 ( 
.A(n_2849),
.Y(n_2897)
);

OAI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2832),
.A2(n_1213),
.B1(n_1214),
.B2(n_1212),
.Y(n_2898)
);

INVx1_ASAP7_75t_SL g2899 ( 
.A(n_2827),
.Y(n_2899)
);

AOI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2869),
.A2(n_2868),
.B1(n_2866),
.B2(n_2843),
.Y(n_2900)
);

INVx6_ASAP7_75t_L g2901 ( 
.A(n_2828),
.Y(n_2901)
);

CKINVDCx5p33_ASAP7_75t_R g2902 ( 
.A(n_2850),
.Y(n_2902)
);

BUFx3_ASAP7_75t_L g2903 ( 
.A(n_2851),
.Y(n_2903)
);

AOI22xp5_ASAP7_75t_SL g2904 ( 
.A1(n_2872),
.A2(n_1488),
.B1(n_1489),
.B2(n_1474),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2855),
.B(n_1775),
.Y(n_2905)
);

INVx6_ASAP7_75t_L g2906 ( 
.A(n_2871),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2864),
.Y(n_2907)
);

AOI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2854),
.A2(n_1224),
.B1(n_1225),
.B2(n_1221),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2881),
.Y(n_2909)
);

BUFx3_ASAP7_75t_L g2910 ( 
.A(n_2859),
.Y(n_2910)
);

AOI22xp33_ASAP7_75t_L g2911 ( 
.A1(n_2833),
.A2(n_1283),
.B1(n_1402),
.B2(n_1259),
.Y(n_2911)
);

INVx3_ASAP7_75t_L g2912 ( 
.A(n_2857),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2853),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2852),
.A2(n_1470),
.B1(n_1653),
.B2(n_1372),
.Y(n_2914)
);

BUFx5_ASAP7_75t_L g2915 ( 
.A(n_2867),
.Y(n_2915)
);

BUFx8_ASAP7_75t_SL g2916 ( 
.A(n_2838),
.Y(n_2916)
);

OAI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2834),
.A2(n_1233),
.B1(n_1234),
.B2(n_1231),
.Y(n_2917)
);

INVx1_ASAP7_75t_SL g2918 ( 
.A(n_2862),
.Y(n_2918)
);

CKINVDCx11_ASAP7_75t_R g2919 ( 
.A(n_2870),
.Y(n_2919)
);

AOI22xp33_ASAP7_75t_SL g2920 ( 
.A1(n_2839),
.A2(n_1653),
.B1(n_1470),
.B2(n_1501),
.Y(n_2920)
);

AO22x1_ASAP7_75t_L g2921 ( 
.A1(n_2877),
.A2(n_1244),
.B1(n_1247),
.B2(n_1243),
.Y(n_2921)
);

INVx6_ASAP7_75t_L g2922 ( 
.A(n_2865),
.Y(n_2922)
);

INVx2_ASAP7_75t_SL g2923 ( 
.A(n_2863),
.Y(n_2923)
);

CKINVDCx5p33_ASAP7_75t_R g2924 ( 
.A(n_2860),
.Y(n_2924)
);

BUFx6f_ASAP7_75t_L g2925 ( 
.A(n_2856),
.Y(n_2925)
);

BUFx4f_ASAP7_75t_SL g2926 ( 
.A(n_2858),
.Y(n_2926)
);

AOI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2842),
.A2(n_1260),
.B1(n_1262),
.B2(n_1256),
.Y(n_2927)
);

OAI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2885),
.A2(n_1270),
.B1(n_1274),
.B2(n_1269),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2863),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2861),
.Y(n_2930)
);

AOI22xp33_ASAP7_75t_L g2931 ( 
.A1(n_2836),
.A2(n_1522),
.B1(n_1530),
.B2(n_1498),
.Y(n_2931)
);

OAI22xp5_ASAP7_75t_L g2932 ( 
.A1(n_2846),
.A2(n_1295),
.B1(n_1299),
.B2(n_1277),
.Y(n_2932)
);

BUFx3_ASAP7_75t_L g2933 ( 
.A(n_2846),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2882),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2884),
.Y(n_2935)
);

AOI22xp33_ASAP7_75t_L g2936 ( 
.A1(n_2879),
.A2(n_1543),
.B1(n_1566),
.B2(n_1534),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2883),
.A2(n_1598),
.B1(n_1611),
.B2(n_1585),
.Y(n_2937)
);

INVx4_ASAP7_75t_L g2938 ( 
.A(n_2845),
.Y(n_2938)
);

BUFx3_ASAP7_75t_L g2939 ( 
.A(n_2848),
.Y(n_2939)
);

AOI22xp33_ASAP7_75t_L g2940 ( 
.A1(n_2847),
.A2(n_1632),
.B1(n_1636),
.B2(n_1617),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2918),
.B(n_2837),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2909),
.Y(n_2942)
);

CKINVDCx20_ASAP7_75t_R g2943 ( 
.A(n_2897),
.Y(n_2943)
);

BUFx2_ASAP7_75t_L g2944 ( 
.A(n_2903),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2892),
.Y(n_2945)
);

OR2x6_ASAP7_75t_L g2946 ( 
.A(n_2886),
.B(n_2841),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2895),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2896),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2915),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2907),
.Y(n_2950)
);

CKINVDCx11_ASAP7_75t_R g2951 ( 
.A(n_2899),
.Y(n_2951)
);

AND2x4_ASAP7_75t_L g2952 ( 
.A(n_2910),
.B(n_2845),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2913),
.B(n_2890),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2915),
.B(n_2837),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_L g2955 ( 
.A1(n_2919),
.A2(n_1637),
.B1(n_1661),
.B2(n_1656),
.Y(n_2955)
);

CKINVDCx5p33_ASAP7_75t_R g2956 ( 
.A(n_2889),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2929),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2901),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2905),
.B(n_1300),
.Y(n_2959)
);

OR2x6_ASAP7_75t_L g2960 ( 
.A(n_2886),
.B(n_2840),
.Y(n_2960)
);

OAI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2887),
.A2(n_2829),
.B(n_2825),
.Y(n_2961)
);

OAI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2920),
.A2(n_2831),
.B(n_1670),
.Y(n_2962)
);

AOI21x1_ASAP7_75t_L g2963 ( 
.A1(n_2932),
.A2(n_1686),
.B(n_1669),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2934),
.Y(n_2964)
);

HB1xp67_ASAP7_75t_L g2965 ( 
.A(n_2935),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2940),
.A2(n_1703),
.B(n_1696),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2912),
.B(n_733),
.Y(n_2967)
);

BUFx2_ASAP7_75t_L g2968 ( 
.A(n_2915),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2923),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2933),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2904),
.B(n_1301),
.Y(n_2971)
);

INVx3_ASAP7_75t_L g2972 ( 
.A(n_2902),
.Y(n_2972)
);

OAI21x1_ASAP7_75t_L g2973 ( 
.A1(n_2931),
.A2(n_1731),
.B(n_1729),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2939),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2906),
.Y(n_2975)
);

AOI22xp33_ASAP7_75t_L g2976 ( 
.A1(n_2926),
.A2(n_1732),
.B1(n_1743),
.B2(n_1733),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2938),
.Y(n_2977)
);

OAI21x1_ASAP7_75t_L g2978 ( 
.A1(n_2936),
.A2(n_1761),
.B(n_1746),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2925),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2922),
.Y(n_2980)
);

OAI21x1_ASAP7_75t_L g2981 ( 
.A1(n_2937),
.A2(n_1765),
.B(n_2561),
.Y(n_2981)
);

HB1xp67_ASAP7_75t_L g2982 ( 
.A(n_2924),
.Y(n_2982)
);

INVx2_ASAP7_75t_SL g2983 ( 
.A(n_2893),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2925),
.Y(n_2984)
);

BUFx2_ASAP7_75t_L g2985 ( 
.A(n_2916),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2930),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2900),
.Y(n_2987)
);

INVx3_ASAP7_75t_L g2988 ( 
.A(n_2972),
.Y(n_2988)
);

OA21x2_ASAP7_75t_L g2989 ( 
.A1(n_2941),
.A2(n_2914),
.B(n_2888),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2947),
.Y(n_2990)
);

BUFx3_ASAP7_75t_L g2991 ( 
.A(n_2958),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2945),
.B(n_2898),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2942),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2987),
.B(n_2927),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2948),
.Y(n_2995)
);

BUFx2_ASAP7_75t_L g2996 ( 
.A(n_2944),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2949),
.Y(n_2997)
);

AO21x2_ASAP7_75t_L g2998 ( 
.A1(n_2964),
.A2(n_2908),
.B(n_2928),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2968),
.Y(n_2999)
);

OR2x2_ASAP7_75t_L g3000 ( 
.A(n_2965),
.B(n_2921),
.Y(n_3000)
);

OA21x2_ASAP7_75t_L g3001 ( 
.A1(n_2974),
.A2(n_2891),
.B(n_2911),
.Y(n_3001)
);

INVx2_ASAP7_75t_SL g3002 ( 
.A(n_2975),
.Y(n_3002)
);

OA21x2_ASAP7_75t_L g3003 ( 
.A1(n_2950),
.A2(n_2957),
.B(n_2977),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2970),
.Y(n_3004)
);

AO21x2_ASAP7_75t_L g3005 ( 
.A1(n_2979),
.A2(n_2917),
.B(n_2894),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2969),
.Y(n_3006)
);

HB1xp67_ASAP7_75t_L g3007 ( 
.A(n_2954),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2984),
.Y(n_3008)
);

HB1xp67_ASAP7_75t_L g3009 ( 
.A(n_2952),
.Y(n_3009)
);

INVxp67_ASAP7_75t_SL g3010 ( 
.A(n_2953),
.Y(n_3010)
);

AOI22xp33_ASAP7_75t_L g3011 ( 
.A1(n_2955),
.A2(n_1529),
.B1(n_1307),
.B2(n_1310),
.Y(n_3011)
);

BUFx3_ASAP7_75t_L g3012 ( 
.A(n_2956),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2980),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2986),
.Y(n_3014)
);

HB1xp67_ASAP7_75t_L g3015 ( 
.A(n_2982),
.Y(n_3015)
);

AND2x4_ASAP7_75t_L g3016 ( 
.A(n_2983),
.B(n_737),
.Y(n_3016)
);

OAI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_2976),
.A2(n_1311),
.B1(n_1325),
.B2(n_1304),
.Y(n_3017)
);

AO21x2_ASAP7_75t_L g3018 ( 
.A1(n_2961),
.A2(n_0),
.B(n_1),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2978),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2951),
.B(n_1529),
.Y(n_3020)
);

INVx3_ASAP7_75t_L g3021 ( 
.A(n_2985),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2973),
.Y(n_3022)
);

AO21x2_ASAP7_75t_L g3023 ( 
.A1(n_2963),
.A2(n_0),
.B(n_3),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2966),
.Y(n_3024)
);

BUFx2_ASAP7_75t_L g3025 ( 
.A(n_2960),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2946),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2946),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2959),
.B(n_1327),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2960),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2971),
.B(n_1328),
.Y(n_3030)
);

CKINVDCx5p33_ASAP7_75t_R g3031 ( 
.A(n_2943),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2967),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2981),
.Y(n_3033)
);

BUFx2_ASAP7_75t_L g3034 ( 
.A(n_2962),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2945),
.B(n_1331),
.Y(n_3035)
);

OR2x2_ASAP7_75t_L g3036 ( 
.A(n_2942),
.B(n_3),
.Y(n_3036)
);

BUFx6f_ASAP7_75t_L g3037 ( 
.A(n_2951),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2942),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2942),
.B(n_4),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2942),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2942),
.Y(n_3041)
);

OR2x2_ASAP7_75t_L g3042 ( 
.A(n_2942),
.B(n_4),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2947),
.Y(n_3043)
);

AND2x4_ASAP7_75t_L g3044 ( 
.A(n_2944),
.B(n_738),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2942),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2999),
.Y(n_3046)
);

BUFx2_ASAP7_75t_L g3047 ( 
.A(n_3025),
.Y(n_3047)
);

AOI22xp33_ASAP7_75t_L g3048 ( 
.A1(n_3034),
.A2(n_1782),
.B1(n_1334),
.B2(n_1362),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2993),
.Y(n_3049)
);

BUFx6f_ASAP7_75t_L g3050 ( 
.A(n_3037),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2996),
.B(n_5),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2997),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_3038),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_3045),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_3040),
.Y(n_3055)
);

INVx3_ASAP7_75t_L g3056 ( 
.A(n_2988),
.Y(n_3056)
);

AND2x2_ASAP7_75t_L g3057 ( 
.A(n_3015),
.B(n_3009),
.Y(n_3057)
);

HB1xp67_ASAP7_75t_L g3058 ( 
.A(n_3007),
.Y(n_3058)
);

INVx3_ASAP7_75t_L g3059 ( 
.A(n_3021),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_3041),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2995),
.Y(n_3061)
);

INVx1_ASAP7_75t_SL g3062 ( 
.A(n_3037),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2990),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_3004),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_3043),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_3010),
.B(n_5),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_3008),
.Y(n_3067)
);

HB1xp67_ASAP7_75t_L g3068 ( 
.A(n_3003),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_3027),
.B(n_6),
.Y(n_3069)
);

AND2x2_ASAP7_75t_L g3070 ( 
.A(n_3026),
.B(n_7),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_3006),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_3029),
.Y(n_3072)
);

AND2x4_ASAP7_75t_L g3073 ( 
.A(n_3014),
.B(n_7),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_3013),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_3000),
.B(n_1332),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3036),
.Y(n_3076)
);

OAI22xp33_ASAP7_75t_L g3077 ( 
.A1(n_2989),
.A2(n_1375),
.B1(n_1378),
.B2(n_1367),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_3002),
.B(n_8),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_3042),
.Y(n_3079)
);

HB1xp67_ASAP7_75t_L g3080 ( 
.A(n_3039),
.Y(n_3080)
);

HB1xp67_ASAP7_75t_L g3081 ( 
.A(n_3039),
.Y(n_3081)
);

INVx4_ASAP7_75t_L g3082 ( 
.A(n_3031),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_3035),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_3019),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2991),
.B(n_3032),
.Y(n_3085)
);

INVxp67_ASAP7_75t_L g3086 ( 
.A(n_3020),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_3022),
.Y(n_3087)
);

BUFx3_ASAP7_75t_L g3088 ( 
.A(n_3012),
.Y(n_3088)
);

BUFx3_ASAP7_75t_L g3089 ( 
.A(n_3044),
.Y(n_3089)
);

HB1xp67_ASAP7_75t_L g3090 ( 
.A(n_3024),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2992),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_3033),
.Y(n_3092)
);

AND2x2_ASAP7_75t_L g3093 ( 
.A(n_3018),
.B(n_8),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2998),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_3023),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2994),
.Y(n_3096)
);

AND2x2_ASAP7_75t_L g3097 ( 
.A(n_3005),
.B(n_9),
.Y(n_3097)
);

INVxp33_ASAP7_75t_L g3098 ( 
.A(n_3028),
.Y(n_3098)
);

OR2x2_ASAP7_75t_L g3099 ( 
.A(n_3001),
.B(n_9),
.Y(n_3099)
);

NAND3xp33_ASAP7_75t_L g3100 ( 
.A(n_3030),
.B(n_1390),
.C(n_1387),
.Y(n_3100)
);

AND2x4_ASAP7_75t_L g3101 ( 
.A(n_3016),
.B(n_10),
.Y(n_3101)
);

INVxp67_ASAP7_75t_L g3102 ( 
.A(n_3017),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_3096),
.B(n_3011),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_3047),
.Y(n_3104)
);

INVxp67_ASAP7_75t_SL g3105 ( 
.A(n_3068),
.Y(n_3105)
);

INVxp67_ASAP7_75t_SL g3106 ( 
.A(n_3094),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_3057),
.B(n_10),
.Y(n_3107)
);

AND2x2_ASAP7_75t_L g3108 ( 
.A(n_3059),
.B(n_11),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_3047),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_3091),
.B(n_1391),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_3067),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_3072),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_3080),
.B(n_3081),
.Y(n_3113)
);

INVx3_ASAP7_75t_SL g3114 ( 
.A(n_3050),
.Y(n_3114)
);

HB1xp67_ASAP7_75t_L g3115 ( 
.A(n_3058),
.Y(n_3115)
);

AND2x2_ASAP7_75t_L g3116 ( 
.A(n_3056),
.B(n_11),
.Y(n_3116)
);

BUFx2_ASAP7_75t_L g3117 ( 
.A(n_3086),
.Y(n_3117)
);

HB1xp67_ASAP7_75t_L g3118 ( 
.A(n_3090),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_3054),
.Y(n_3119)
);

INVx3_ASAP7_75t_L g3120 ( 
.A(n_3050),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_3055),
.Y(n_3121)
);

NOR2xp67_ASAP7_75t_L g3122 ( 
.A(n_3082),
.B(n_12),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_3049),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_SL g3124 ( 
.A(n_3077),
.B(n_1392),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3053),
.Y(n_3125)
);

OR2x2_ASAP7_75t_L g3126 ( 
.A(n_3076),
.B(n_12),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_3060),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_3085),
.B(n_13),
.Y(n_3128)
);

INVx2_ASAP7_75t_SL g3129 ( 
.A(n_3062),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_3064),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_3061),
.Y(n_3131)
);

BUFx3_ASAP7_75t_L g3132 ( 
.A(n_3088),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_3098),
.B(n_1397),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3084),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_3074),
.Y(n_3135)
);

AND2x2_ASAP7_75t_L g3136 ( 
.A(n_3079),
.B(n_13),
.Y(n_3136)
);

INVx4_ASAP7_75t_R g3137 ( 
.A(n_3089),
.Y(n_3137)
);

INVxp67_ASAP7_75t_SL g3138 ( 
.A(n_3099),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_3083),
.B(n_1400),
.Y(n_3139)
);

CKINVDCx20_ASAP7_75t_R g3140 ( 
.A(n_3102),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3087),
.Y(n_3141)
);

AND2x2_ASAP7_75t_L g3142 ( 
.A(n_3046),
.B(n_15),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3071),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_3063),
.B(n_1404),
.Y(n_3144)
);

AND2x4_ASAP7_75t_L g3145 ( 
.A(n_3065),
.B(n_3069),
.Y(n_3145)
);

INVx4_ASAP7_75t_L g3146 ( 
.A(n_3073),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_3052),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3092),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_3066),
.B(n_15),
.Y(n_3149)
);

BUFx6f_ASAP7_75t_L g3150 ( 
.A(n_3078),
.Y(n_3150)
);

NOR2x1_ASAP7_75t_L g3151 ( 
.A(n_3097),
.B(n_17),
.Y(n_3151)
);

OR2x2_ASAP7_75t_SL g3152 ( 
.A(n_3075),
.B(n_17),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3095),
.Y(n_3153)
);

AND2x2_ASAP7_75t_L g3154 ( 
.A(n_3051),
.B(n_18),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3070),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_3093),
.B(n_18),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_3101),
.B(n_19),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_3048),
.B(n_20),
.Y(n_3158)
);

INVx4_ASAP7_75t_L g3159 ( 
.A(n_3100),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3049),
.Y(n_3160)
);

HB1xp67_ASAP7_75t_L g3161 ( 
.A(n_3058),
.Y(n_3161)
);

OR2x2_ASAP7_75t_L g3162 ( 
.A(n_3080),
.B(n_21),
.Y(n_3162)
);

OR2x2_ASAP7_75t_L g3163 ( 
.A(n_3080),
.B(n_21),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_3047),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_3047),
.Y(n_3165)
);

CKINVDCx16_ASAP7_75t_R g3166 ( 
.A(n_3050),
.Y(n_3166)
);

OAI21xp5_ASAP7_75t_SL g3167 ( 
.A1(n_3077),
.A2(n_33),
.B(n_22),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_3049),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_3047),
.Y(n_3169)
);

BUFx6f_ASAP7_75t_L g3170 ( 
.A(n_3050),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3049),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3049),
.Y(n_3172)
);

BUFx2_ASAP7_75t_L g3173 ( 
.A(n_3047),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_3057),
.B(n_22),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3049),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_3096),
.B(n_1405),
.Y(n_3176)
);

OAI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_3099),
.A2(n_1415),
.B1(n_1420),
.B2(n_1412),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_3047),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3049),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_3047),
.Y(n_3180)
);

OAI221xp5_ASAP7_75t_L g3181 ( 
.A1(n_3048),
.A2(n_1428),
.B1(n_1431),
.B2(n_1424),
.C(n_1423),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3049),
.Y(n_3182)
);

AND2x2_ASAP7_75t_L g3183 ( 
.A(n_3057),
.B(n_23),
.Y(n_3183)
);

BUFx2_ASAP7_75t_L g3184 ( 
.A(n_3047),
.Y(n_3184)
);

NOR2x1_ASAP7_75t_SL g3185 ( 
.A(n_3094),
.B(n_23),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_3057),
.B(n_24),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_3057),
.B(n_24),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_3047),
.Y(n_3188)
);

OAI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_3099),
.A2(n_1436),
.B1(n_1441),
.B2(n_1433),
.Y(n_3189)
);

HB1xp67_ASAP7_75t_L g3190 ( 
.A(n_3058),
.Y(n_3190)
);

AND2x2_ASAP7_75t_L g3191 ( 
.A(n_3057),
.B(n_25),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3049),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_3047),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_3096),
.B(n_1445),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3096),
.B(n_1451),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_3057),
.B(n_28),
.Y(n_3196)
);

BUFx2_ASAP7_75t_L g3197 ( 
.A(n_3047),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3049),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3049),
.Y(n_3199)
);

AND2x2_ASAP7_75t_L g3200 ( 
.A(n_3057),
.B(n_28),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3049),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_3096),
.B(n_1456),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_3057),
.B(n_29),
.Y(n_3203)
);

OR2x2_ASAP7_75t_L g3204 ( 
.A(n_3080),
.B(n_30),
.Y(n_3204)
);

AND2x2_ASAP7_75t_L g3205 ( 
.A(n_3057),
.B(n_31),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_3057),
.B(n_31),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_3057),
.B(n_33),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3049),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_3057),
.B(n_34),
.Y(n_3209)
);

HB1xp67_ASAP7_75t_L g3210 ( 
.A(n_3058),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_3047),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_3057),
.B(n_34),
.Y(n_3212)
);

HB1xp67_ASAP7_75t_L g3213 ( 
.A(n_3058),
.Y(n_3213)
);

OR2x2_ASAP7_75t_L g3214 ( 
.A(n_3138),
.B(n_35),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3143),
.Y(n_3215)
);

OR2x2_ASAP7_75t_L g3216 ( 
.A(n_3115),
.B(n_35),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3123),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3125),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3127),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_3113),
.B(n_36),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_3173),
.B(n_36),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3184),
.B(n_37),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_3117),
.B(n_1460),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_3161),
.B(n_1463),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_3190),
.B(n_1464),
.Y(n_3225)
);

INVx2_ASAP7_75t_SL g3226 ( 
.A(n_3137),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3131),
.Y(n_3227)
);

HB1xp67_ASAP7_75t_L g3228 ( 
.A(n_3197),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_3104),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3160),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3168),
.Y(n_3231)
);

INVxp67_ASAP7_75t_SL g3232 ( 
.A(n_3185),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_3109),
.B(n_37),
.Y(n_3233)
);

INVx3_ASAP7_75t_L g3234 ( 
.A(n_3166),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_3164),
.B(n_38),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3171),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_3165),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_3129),
.B(n_39),
.Y(n_3238)
);

HB1xp67_ASAP7_75t_L g3239 ( 
.A(n_3210),
.Y(n_3239)
);

OR2x2_ASAP7_75t_L g3240 ( 
.A(n_3213),
.B(n_39),
.Y(n_3240)
);

OR2x2_ASAP7_75t_L g3241 ( 
.A(n_3169),
.B(n_40),
.Y(n_3241)
);

OR2x2_ASAP7_75t_L g3242 ( 
.A(n_3178),
.B(n_3180),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3172),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3103),
.B(n_1466),
.Y(n_3244)
);

AND2x2_ASAP7_75t_L g3245 ( 
.A(n_3188),
.B(n_40),
.Y(n_3245)
);

OR2x2_ASAP7_75t_L g3246 ( 
.A(n_3193),
.B(n_41),
.Y(n_3246)
);

NOR2xp67_ASAP7_75t_SL g3247 ( 
.A(n_3167),
.B(n_1479),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3175),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3211),
.B(n_3145),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3179),
.Y(n_3250)
);

OR2x2_ASAP7_75t_L g3251 ( 
.A(n_3112),
.B(n_41),
.Y(n_3251)
);

AND2x4_ASAP7_75t_SL g3252 ( 
.A(n_3170),
.B(n_42),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_3155),
.B(n_43),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_3150),
.B(n_44),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_3150),
.B(n_44),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3147),
.B(n_3212),
.Y(n_3256)
);

AND2x2_ASAP7_75t_L g3257 ( 
.A(n_3209),
.B(n_3196),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_3119),
.Y(n_3258)
);

AND2x2_ASAP7_75t_L g3259 ( 
.A(n_3107),
.B(n_45),
.Y(n_3259)
);

BUFx3_ASAP7_75t_L g3260 ( 
.A(n_3114),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3182),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_3174),
.B(n_45),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_3183),
.B(n_3203),
.Y(n_3263)
);

AND2x2_ASAP7_75t_L g3264 ( 
.A(n_3186),
.B(n_46),
.Y(n_3264)
);

OR2x2_ASAP7_75t_L g3265 ( 
.A(n_3121),
.B(n_47),
.Y(n_3265)
);

AND2x2_ASAP7_75t_L g3266 ( 
.A(n_3187),
.B(n_48),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_3135),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_3191),
.B(n_48),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3111),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3142),
.B(n_1482),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_3132),
.B(n_50),
.Y(n_3271)
);

OR2x2_ASAP7_75t_L g3272 ( 
.A(n_3130),
.B(n_52),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_3208),
.B(n_1485),
.Y(n_3273)
);

NOR2x1_ASAP7_75t_L g3274 ( 
.A(n_3151),
.B(n_53),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_3207),
.B(n_53),
.Y(n_3275)
);

AND2x4_ASAP7_75t_L g3276 ( 
.A(n_3120),
.B(n_54),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3192),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3200),
.B(n_56),
.Y(n_3278)
);

AND2x4_ASAP7_75t_L g3279 ( 
.A(n_3146),
.B(n_57),
.Y(n_3279)
);

HB1xp67_ASAP7_75t_L g3280 ( 
.A(n_3118),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_3153),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_3205),
.B(n_57),
.Y(n_3282)
);

AND2x2_ASAP7_75t_SL g3283 ( 
.A(n_3159),
.B(n_58),
.Y(n_3283)
);

NOR3xp33_ASAP7_75t_L g3284 ( 
.A(n_3124),
.B(n_1493),
.C(n_1490),
.Y(n_3284)
);

BUFx6f_ASAP7_75t_L g3285 ( 
.A(n_3170),
.Y(n_3285)
);

AND2x2_ASAP7_75t_L g3286 ( 
.A(n_3206),
.B(n_58),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_3105),
.B(n_59),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3198),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3199),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3201),
.B(n_1494),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3134),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3141),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_3122),
.B(n_3177),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3136),
.B(n_1495),
.Y(n_3294)
);

HB1xp67_ASAP7_75t_L g3295 ( 
.A(n_3148),
.Y(n_3295)
);

INVxp67_ASAP7_75t_L g3296 ( 
.A(n_3110),
.Y(n_3296)
);

INVx3_ASAP7_75t_L g3297 ( 
.A(n_3116),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_3128),
.B(n_3108),
.Y(n_3298)
);

HB1xp67_ASAP7_75t_L g3299 ( 
.A(n_3162),
.Y(n_3299)
);

INVx3_ASAP7_75t_L g3300 ( 
.A(n_3126),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3144),
.Y(n_3301)
);

AND2x2_ASAP7_75t_L g3302 ( 
.A(n_3106),
.B(n_59),
.Y(n_3302)
);

INVxp67_ASAP7_75t_SL g3303 ( 
.A(n_3140),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3163),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3204),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3189),
.B(n_1497),
.Y(n_3306)
);

INVx3_ASAP7_75t_L g3307 ( 
.A(n_3157),
.Y(n_3307)
);

OR2x2_ASAP7_75t_L g3308 ( 
.A(n_3156),
.B(n_60),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3176),
.Y(n_3309)
);

AND2x4_ASAP7_75t_L g3310 ( 
.A(n_3149),
.B(n_60),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3194),
.B(n_1502),
.Y(n_3311)
);

OR2x2_ASAP7_75t_L g3312 ( 
.A(n_3195),
.B(n_61),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3202),
.B(n_1505),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3139),
.B(n_1508),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3152),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_3154),
.Y(n_3316)
);

OR2x2_ASAP7_75t_L g3317 ( 
.A(n_3133),
.B(n_61),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3158),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3181),
.B(n_62),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3143),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3113),
.B(n_62),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3143),
.Y(n_3322)
);

HB1xp67_ASAP7_75t_L g3323 ( 
.A(n_3173),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3143),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_3138),
.B(n_1511),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3138),
.B(n_1513),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3143),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3138),
.B(n_1514),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3143),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3143),
.Y(n_3330)
);

OR2x2_ASAP7_75t_L g3331 ( 
.A(n_3138),
.B(n_63),
.Y(n_3331)
);

OR2x2_ASAP7_75t_L g3332 ( 
.A(n_3138),
.B(n_63),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3138),
.B(n_1517),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_3113),
.B(n_64),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_3113),
.B(n_64),
.Y(n_3335)
);

OR2x2_ASAP7_75t_L g3336 ( 
.A(n_3138),
.B(n_65),
.Y(n_3336)
);

AND2x2_ASAP7_75t_L g3337 ( 
.A(n_3113),
.B(n_65),
.Y(n_3337)
);

INVx2_ASAP7_75t_SL g3338 ( 
.A(n_3137),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_SL g3339 ( 
.A(n_3166),
.B(n_1528),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_3173),
.Y(n_3340)
);

OR2x2_ASAP7_75t_L g3341 ( 
.A(n_3138),
.B(n_66),
.Y(n_3341)
);

AND2x2_ASAP7_75t_L g3342 ( 
.A(n_3113),
.B(n_66),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_3113),
.B(n_67),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3143),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3113),
.B(n_67),
.Y(n_3345)
);

AND2x4_ASAP7_75t_L g3346 ( 
.A(n_3129),
.B(n_68),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3113),
.B(n_68),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3173),
.Y(n_3348)
);

AND2x4_ASAP7_75t_L g3349 ( 
.A(n_3129),
.B(n_69),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3173),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3138),
.B(n_1532),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3113),
.B(n_69),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3173),
.Y(n_3353)
);

OR2x2_ASAP7_75t_L g3354 ( 
.A(n_3138),
.B(n_70),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_3113),
.B(n_70),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3143),
.Y(n_3356)
);

HB1xp67_ASAP7_75t_L g3357 ( 
.A(n_3173),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3143),
.Y(n_3358)
);

INVx3_ASAP7_75t_L g3359 ( 
.A(n_3166),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3138),
.B(n_1535),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3113),
.B(n_71),
.Y(n_3361)
);

AOI22xp33_ASAP7_75t_L g3362 ( 
.A1(n_3159),
.A2(n_1538),
.B1(n_1540),
.B2(n_1537),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3138),
.B(n_1544),
.Y(n_3363)
);

INVx3_ASAP7_75t_L g3364 ( 
.A(n_3166),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3143),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3113),
.B(n_71),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3143),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3113),
.B(n_72),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_3234),
.B(n_73),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_3359),
.B(n_1756),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3364),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3232),
.B(n_1547),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3226),
.B(n_73),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3215),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3217),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3218),
.Y(n_3376)
);

OR2x2_ASAP7_75t_L g3377 ( 
.A(n_3242),
.B(n_3239),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3219),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3300),
.B(n_1551),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3227),
.Y(n_3380)
);

INVxp67_ASAP7_75t_L g3381 ( 
.A(n_3274),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3230),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3231),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3299),
.B(n_1552),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3305),
.B(n_1555),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3236),
.Y(n_3386)
);

NOR2xp33_ASAP7_75t_L g3387 ( 
.A(n_3260),
.B(n_1763),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3243),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3309),
.B(n_1557),
.Y(n_3389)
);

OR2x2_ASAP7_75t_L g3390 ( 
.A(n_3340),
.B(n_74),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3248),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3250),
.Y(n_3392)
);

HB1xp67_ASAP7_75t_L g3393 ( 
.A(n_3228),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3304),
.B(n_3301),
.Y(n_3394)
);

NAND2x1p5_ASAP7_75t_L g3395 ( 
.A(n_3338),
.B(n_74),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3261),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3318),
.B(n_1558),
.Y(n_3397)
);

OAI21xp33_ASAP7_75t_SL g3398 ( 
.A1(n_3323),
.A2(n_75),
.B(n_76),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3287),
.B(n_1561),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3249),
.B(n_75),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3348),
.B(n_76),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3285),
.Y(n_3402)
);

OR2x2_ASAP7_75t_L g3403 ( 
.A(n_3350),
.B(n_77),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3296),
.B(n_1563),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3277),
.Y(n_3405)
);

OR2x2_ASAP7_75t_SL g3406 ( 
.A(n_3315),
.B(n_77),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3288),
.Y(n_3407)
);

AO22x1_ASAP7_75t_L g3408 ( 
.A1(n_3303),
.A2(n_3302),
.B1(n_3222),
.B2(n_3221),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3316),
.B(n_1564),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3289),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3353),
.B(n_3357),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3291),
.Y(n_3412)
);

OR2x2_ASAP7_75t_L g3413 ( 
.A(n_3280),
.B(n_78),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_3256),
.B(n_78),
.Y(n_3414)
);

HB1xp67_ASAP7_75t_L g3415 ( 
.A(n_3295),
.Y(n_3415)
);

HB1xp67_ASAP7_75t_L g3416 ( 
.A(n_3258),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3220),
.B(n_1567),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3292),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3320),
.Y(n_3419)
);

OR2x2_ASAP7_75t_L g3420 ( 
.A(n_3229),
.B(n_79),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3322),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3321),
.B(n_1568),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3285),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3307),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3324),
.Y(n_3425)
);

INVxp67_ASAP7_75t_SL g3426 ( 
.A(n_3293),
.Y(n_3426)
);

OR2x2_ASAP7_75t_L g3427 ( 
.A(n_3237),
.B(n_80),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3334),
.B(n_1572),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3327),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_3297),
.B(n_80),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3298),
.B(n_81),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3329),
.Y(n_3432)
);

AND2x2_ASAP7_75t_L g3433 ( 
.A(n_3257),
.B(n_81),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3330),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3344),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3267),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_3263),
.B(n_82),
.Y(n_3437)
);

AND2x2_ASAP7_75t_L g3438 ( 
.A(n_3335),
.B(n_83),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3356),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3358),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3337),
.B(n_84),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_3269),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3265),
.Y(n_3443)
);

INVx2_ASAP7_75t_L g3444 ( 
.A(n_3272),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3342),
.B(n_85),
.Y(n_3445)
);

AND2x2_ASAP7_75t_L g3446 ( 
.A(n_3343),
.B(n_86),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3345),
.B(n_1575),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3347),
.B(n_1577),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3365),
.Y(n_3449)
);

AND2x2_ASAP7_75t_L g3450 ( 
.A(n_3352),
.B(n_86),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_3244),
.B(n_1581),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_3355),
.B(n_88),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_3251),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3367),
.Y(n_3454)
);

OAI22xp5_ASAP7_75t_L g3455 ( 
.A1(n_3283),
.A2(n_1606),
.B1(n_1633),
.B2(n_1592),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3281),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3361),
.B(n_88),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3366),
.B(n_90),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_3368),
.B(n_91),
.Y(n_3459)
);

OR2x2_ASAP7_75t_L g3460 ( 
.A(n_3241),
.B(n_3246),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_3253),
.B(n_92),
.Y(n_3461)
);

HB1xp67_ASAP7_75t_L g3462 ( 
.A(n_3214),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_3233),
.B(n_93),
.Y(n_3463)
);

INVx3_ASAP7_75t_L g3464 ( 
.A(n_3279),
.Y(n_3464)
);

AND2x2_ASAP7_75t_L g3465 ( 
.A(n_3235),
.B(n_94),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3245),
.Y(n_3466)
);

NAND2x1_ASAP7_75t_L g3467 ( 
.A(n_3238),
.B(n_95),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3331),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3332),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3336),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3341),
.B(n_96),
.Y(n_3471)
);

OAI21xp33_ASAP7_75t_L g3472 ( 
.A1(n_3362),
.A2(n_1588),
.B(n_1586),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3354),
.B(n_1590),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3254),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3216),
.Y(n_3475)
);

AND2x2_ASAP7_75t_L g3476 ( 
.A(n_3255),
.B(n_97),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3325),
.B(n_1596),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3240),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3346),
.B(n_97),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3273),
.Y(n_3480)
);

OR2x6_ASAP7_75t_L g3481 ( 
.A(n_3349),
.B(n_100),
.Y(n_3481)
);

BUFx3_ASAP7_75t_L g3482 ( 
.A(n_3271),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3326),
.B(n_1601),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3276),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3328),
.B(n_1602),
.Y(n_3485)
);

OR2x2_ASAP7_75t_L g3486 ( 
.A(n_3224),
.B(n_100),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3290),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3333),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_3225),
.B(n_101),
.Y(n_3489)
);

NAND2x2_ASAP7_75t_L g3490 ( 
.A(n_3312),
.B(n_101),
.Y(n_3490)
);

BUFx2_ASAP7_75t_L g3491 ( 
.A(n_3310),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3351),
.A2(n_1764),
.B(n_1758),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3360),
.Y(n_3493)
);

BUFx2_ASAP7_75t_L g3494 ( 
.A(n_3308),
.Y(n_3494)
);

INVxp67_ASAP7_75t_SL g3495 ( 
.A(n_3363),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3259),
.B(n_103),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3223),
.B(n_3262),
.Y(n_3497)
);

INVxp67_ASAP7_75t_L g3498 ( 
.A(n_3339),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3264),
.B(n_103),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3266),
.B(n_104),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3268),
.Y(n_3501)
);

INVx2_ASAP7_75t_SL g3502 ( 
.A(n_3252),
.Y(n_3502)
);

OR2x2_ASAP7_75t_L g3503 ( 
.A(n_3317),
.B(n_105),
.Y(n_3503)
);

OR2x2_ASAP7_75t_L g3504 ( 
.A(n_3270),
.B(n_105),
.Y(n_3504)
);

INVx3_ASAP7_75t_L g3505 ( 
.A(n_3275),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3278),
.B(n_1609),
.Y(n_3506)
);

AND2x4_ASAP7_75t_L g3507 ( 
.A(n_3282),
.B(n_107),
.Y(n_3507)
);

INVx3_ASAP7_75t_L g3508 ( 
.A(n_3286),
.Y(n_3508)
);

AOI32xp33_ASAP7_75t_L g3509 ( 
.A1(n_3319),
.A2(n_1613),
.A3(n_1618),
.B1(n_1612),
.B2(n_1610),
.Y(n_3509)
);

OR2x2_ASAP7_75t_L g3510 ( 
.A(n_3294),
.B(n_107),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3311),
.Y(n_3511)
);

NAND2x1p5_ASAP7_75t_L g3512 ( 
.A(n_3247),
.B(n_108),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3313),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3306),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3314),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3284),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3215),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3234),
.Y(n_3518)
);

OAI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_3274),
.A2(n_1623),
.B(n_1621),
.Y(n_3519)
);

OR2x2_ASAP7_75t_L g3520 ( 
.A(n_3242),
.B(n_109),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3215),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3232),
.B(n_1624),
.Y(n_3522)
);

OAI21xp5_ASAP7_75t_L g3523 ( 
.A1(n_3274),
.A2(n_1627),
.B(n_1626),
.Y(n_3523)
);

HB1xp67_ASAP7_75t_L g3524 ( 
.A(n_3228),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3232),
.B(n_1628),
.Y(n_3525)
);

NAND2x1_ASAP7_75t_L g3526 ( 
.A(n_3234),
.B(n_109),
.Y(n_3526)
);

OR2x6_ASAP7_75t_L g3527 ( 
.A(n_3226),
.B(n_110),
.Y(n_3527)
);

OR2x2_ASAP7_75t_L g3528 ( 
.A(n_3242),
.B(n_111),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3234),
.B(n_111),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3215),
.Y(n_3530)
);

INVx2_ASAP7_75t_L g3531 ( 
.A(n_3234),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3234),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3215),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3215),
.Y(n_3534)
);

OR2x2_ASAP7_75t_L g3535 ( 
.A(n_3242),
.B(n_112),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3232),
.B(n_1630),
.Y(n_3536)
);

NAND2x1_ASAP7_75t_L g3537 ( 
.A(n_3234),
.B(n_113),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3234),
.B(n_114),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3234),
.B(n_114),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3234),
.B(n_115),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3215),
.Y(n_3541)
);

AND2x2_ASAP7_75t_L g3542 ( 
.A(n_3234),
.B(n_115),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3234),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3232),
.B(n_1635),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3232),
.B(n_1640),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3232),
.B(n_1641),
.Y(n_3546)
);

BUFx2_ASAP7_75t_L g3547 ( 
.A(n_3234),
.Y(n_3547)
);

AOI22xp33_ASAP7_75t_L g3548 ( 
.A1(n_3247),
.A2(n_1643),
.B1(n_1646),
.B2(n_1642),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_3234),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3234),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3215),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3215),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3232),
.B(n_1651),
.Y(n_3553)
);

AND2x4_ASAP7_75t_L g3554 ( 
.A(n_3226),
.B(n_116),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_3234),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3234),
.B(n_116),
.Y(n_3556)
);

INVx1_ASAP7_75t_SL g3557 ( 
.A(n_3260),
.Y(n_3557)
);

NAND3xp33_ASAP7_75t_L g3558 ( 
.A(n_3274),
.B(n_1779),
.C(n_1654),
.Y(n_3558)
);

AND2x4_ASAP7_75t_SL g3559 ( 
.A(n_3527),
.B(n_117),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3381),
.B(n_1652),
.Y(n_3560)
);

OAI22xp33_ASAP7_75t_L g3561 ( 
.A1(n_3426),
.A2(n_1658),
.B1(n_1667),
.B2(n_1659),
.Y(n_3561)
);

AOI22xp5_ASAP7_75t_L g3562 ( 
.A1(n_3547),
.A2(n_1671),
.B1(n_1673),
.B2(n_1655),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3408),
.B(n_1674),
.Y(n_3563)
);

AO221x2_ASAP7_75t_L g3564 ( 
.A1(n_3398),
.A2(n_120),
.B1(n_117),
.B2(n_118),
.C(n_121),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3415),
.Y(n_3565)
);

AO221x2_ASAP7_75t_L g3566 ( 
.A1(n_3371),
.A2(n_122),
.B1(n_124),
.B2(n_121),
.C(n_123),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3464),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3505),
.B(n_3508),
.Y(n_3568)
);

AO221x2_ASAP7_75t_L g3569 ( 
.A1(n_3518),
.A2(n_123),
.B1(n_126),
.B2(n_122),
.C(n_125),
.Y(n_3569)
);

NAND2xp33_ASAP7_75t_SL g3570 ( 
.A(n_3526),
.B(n_1682),
.Y(n_3570)
);

OAI221xp5_ASAP7_75t_L g3571 ( 
.A1(n_3519),
.A2(n_3523),
.B1(n_3543),
.B2(n_3532),
.C(n_3531),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3474),
.B(n_1688),
.Y(n_3572)
);

NAND2xp33_ASAP7_75t_SL g3573 ( 
.A(n_3537),
.B(n_1689),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3494),
.B(n_1690),
.Y(n_3574)
);

INVx2_ASAP7_75t_SL g3575 ( 
.A(n_3482),
.Y(n_3575)
);

OR2x2_ASAP7_75t_L g3576 ( 
.A(n_3377),
.B(n_118),
.Y(n_3576)
);

NAND2xp33_ASAP7_75t_SL g3577 ( 
.A(n_3467),
.B(n_3491),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3501),
.B(n_1693),
.Y(n_3578)
);

NAND2x1_ASAP7_75t_L g3579 ( 
.A(n_3411),
.B(n_127),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3466),
.B(n_1697),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3393),
.B(n_1698),
.Y(n_3581)
);

OAI22xp33_ASAP7_75t_L g3582 ( 
.A1(n_3549),
.A2(n_1700),
.B1(n_1706),
.B2(n_1699),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_SL g3583 ( 
.A(n_3557),
.B(n_1707),
.Y(n_3583)
);

NAND2xp33_ASAP7_75t_SL g3584 ( 
.A(n_3462),
.B(n_1708),
.Y(n_3584)
);

AO221x2_ASAP7_75t_L g3585 ( 
.A1(n_3514),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3524),
.B(n_1715),
.Y(n_3586)
);

INVxp33_ASAP7_75t_SL g3587 ( 
.A(n_3455),
.Y(n_3587)
);

AO221x2_ASAP7_75t_L g3588 ( 
.A1(n_3550),
.A2(n_130),
.B1(n_132),
.B2(n_129),
.C(n_131),
.Y(n_3588)
);

OAI22xp33_ASAP7_75t_L g3589 ( 
.A1(n_3555),
.A2(n_1718),
.B1(n_1721),
.B2(n_1716),
.Y(n_3589)
);

OAI221xp5_ASAP7_75t_L g3590 ( 
.A1(n_3509),
.A2(n_1727),
.B1(n_1735),
.B2(n_1726),
.C(n_1722),
.Y(n_3590)
);

OAI221xp5_ASAP7_75t_L g3591 ( 
.A1(n_3558),
.A2(n_1745),
.B1(n_1747),
.B2(n_1741),
.C(n_1737),
.Y(n_3591)
);

OAI22xp33_ASAP7_75t_L g3592 ( 
.A1(n_3424),
.A2(n_1749),
.B1(n_1770),
.B2(n_1751),
.Y(n_3592)
);

NAND2xp33_ASAP7_75t_SL g3593 ( 
.A(n_3502),
.B(n_128),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_3495),
.A2(n_1235),
.B1(n_1258),
.B2(n_1232),
.Y(n_3594)
);

AO221x2_ASAP7_75t_L g3595 ( 
.A1(n_3488),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_3595)
);

OAI221xp5_ASAP7_75t_L g3596 ( 
.A1(n_3394),
.A2(n_1267),
.B1(n_1278),
.B2(n_1266),
.C(n_1264),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3468),
.B(n_134),
.Y(n_3597)
);

CKINVDCx20_ASAP7_75t_R g3598 ( 
.A(n_3406),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3374),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3469),
.B(n_136),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3470),
.B(n_136),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3475),
.B(n_137),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3478),
.B(n_138),
.Y(n_3603)
);

AOI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3480),
.A2(n_1288),
.B1(n_1289),
.B2(n_1287),
.Y(n_3604)
);

AO221x2_ASAP7_75t_L g3605 ( 
.A1(n_3493),
.A2(n_140),
.B1(n_142),
.B2(n_139),
.C(n_141),
.Y(n_3605)
);

CKINVDCx5p33_ASAP7_75t_R g3606 ( 
.A(n_3527),
.Y(n_3606)
);

NOR2x1_ASAP7_75t_L g3607 ( 
.A(n_3372),
.B(n_138),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_SL g3608 ( 
.A(n_3498),
.B(n_1291),
.Y(n_3608)
);

AND2x2_ASAP7_75t_L g3609 ( 
.A(n_3402),
.B(n_142),
.Y(n_3609)
);

NOR2xp67_ASAP7_75t_L g3610 ( 
.A(n_3460),
.B(n_143),
.Y(n_3610)
);

INVxp67_ASAP7_75t_L g3611 ( 
.A(n_3423),
.Y(n_3611)
);

OAI22xp33_ASAP7_75t_L g3612 ( 
.A1(n_3413),
.A2(n_1302),
.B1(n_1313),
.B2(n_1292),
.Y(n_3612)
);

AO221x2_ASAP7_75t_L g3613 ( 
.A1(n_3487),
.A2(n_148),
.B1(n_150),
.B2(n_145),
.C(n_149),
.Y(n_3613)
);

NAND2xp33_ASAP7_75t_SL g3614 ( 
.A(n_3484),
.B(n_144),
.Y(n_3614)
);

AO221x2_ASAP7_75t_L g3615 ( 
.A1(n_3497),
.A2(n_149),
.B1(n_144),
.B2(n_148),
.C(n_150),
.Y(n_3615)
);

INVxp33_ASAP7_75t_SL g3616 ( 
.A(n_3373),
.Y(n_3616)
);

INVxp67_ASAP7_75t_L g3617 ( 
.A(n_3522),
.Y(n_3617)
);

INVx2_ASAP7_75t_L g3618 ( 
.A(n_3420),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3443),
.B(n_151),
.Y(n_3619)
);

INVx2_ASAP7_75t_SL g3620 ( 
.A(n_3554),
.Y(n_3620)
);

NAND2xp33_ASAP7_75t_SL g3621 ( 
.A(n_3520),
.B(n_151),
.Y(n_3621)
);

AND2x4_ASAP7_75t_L g3622 ( 
.A(n_3444),
.B(n_152),
.Y(n_3622)
);

AND2x4_ASAP7_75t_L g3623 ( 
.A(n_3453),
.B(n_153),
.Y(n_3623)
);

INVx3_ASAP7_75t_L g3624 ( 
.A(n_3395),
.Y(n_3624)
);

OAI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3490),
.A2(n_1762),
.B1(n_1317),
.B2(n_1319),
.Y(n_3625)
);

INVxp33_ASAP7_75t_SL g3626 ( 
.A(n_3387),
.Y(n_3626)
);

INVxp67_ASAP7_75t_SL g3627 ( 
.A(n_3384),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3515),
.B(n_3511),
.Y(n_3628)
);

OAI22xp33_ASAP7_75t_L g3629 ( 
.A1(n_3528),
.A2(n_1769),
.B1(n_1321),
.B2(n_1323),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3525),
.B(n_153),
.Y(n_3630)
);

AO221x2_ASAP7_75t_L g3631 ( 
.A1(n_3513),
.A2(n_157),
.B1(n_154),
.B2(n_155),
.C(n_160),
.Y(n_3631)
);

OAI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3535),
.A2(n_1759),
.B1(n_1702),
.B2(n_1337),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_3536),
.B(n_154),
.Y(n_3633)
);

CKINVDCx5p33_ASAP7_75t_R g3634 ( 
.A(n_3481),
.Y(n_3634)
);

CKINVDCx5p33_ASAP7_75t_R g3635 ( 
.A(n_3481),
.Y(n_3635)
);

OAI22xp33_ASAP7_75t_L g3636 ( 
.A1(n_3416),
.A2(n_1781),
.B1(n_1738),
.B2(n_1342),
.Y(n_3636)
);

OAI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3512),
.A2(n_1744),
.B1(n_1344),
.B2(n_1347),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3544),
.B(n_157),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3375),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_3545),
.B(n_1316),
.Y(n_3640)
);

NOR4xp25_ASAP7_75t_SL g3641 ( 
.A(n_3376),
.B(n_1355),
.C(n_1359),
.D(n_1348),
.Y(n_3641)
);

NAND2xp33_ASAP7_75t_R g3642 ( 
.A(n_3546),
.B(n_163),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3553),
.B(n_161),
.Y(n_3643)
);

NAND2xp33_ASAP7_75t_SL g3644 ( 
.A(n_3369),
.B(n_163),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3400),
.B(n_164),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3401),
.B(n_164),
.Y(n_3646)
);

NAND2xp33_ASAP7_75t_SL g3647 ( 
.A(n_3529),
.B(n_165),
.Y(n_3647)
);

OAI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3390),
.A2(n_1768),
.B1(n_1691),
.B2(n_1361),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3538),
.B(n_166),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3378),
.Y(n_3650)
);

AND2x4_ASAP7_75t_L g3651 ( 
.A(n_3539),
.B(n_167),
.Y(n_3651)
);

CKINVDCx5p33_ASAP7_75t_R g3652 ( 
.A(n_3516),
.Y(n_3652)
);

INVxp67_ASAP7_75t_L g3653 ( 
.A(n_3403),
.Y(n_3653)
);

AND2x4_ASAP7_75t_SL g3654 ( 
.A(n_3507),
.B(n_168),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3540),
.B(n_168),
.Y(n_3655)
);

AO221x2_ASAP7_75t_L g3656 ( 
.A1(n_3417),
.A2(n_171),
.B1(n_174),
.B2(n_170),
.C(n_173),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3542),
.B(n_169),
.Y(n_3657)
);

CKINVDCx5p33_ASAP7_75t_R g3658 ( 
.A(n_3556),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3414),
.B(n_169),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3433),
.B(n_170),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3437),
.B(n_173),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3431),
.B(n_175),
.Y(n_3662)
);

INVxp67_ASAP7_75t_L g3663 ( 
.A(n_3427),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3380),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3436),
.B(n_176),
.Y(n_3665)
);

NAND2xp33_ASAP7_75t_SL g3666 ( 
.A(n_3430),
.B(n_176),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3471),
.B(n_177),
.Y(n_3667)
);

NAND2xp33_ASAP7_75t_SL g3668 ( 
.A(n_3503),
.B(n_177),
.Y(n_3668)
);

NAND2xp33_ASAP7_75t_SL g3669 ( 
.A(n_3438),
.B(n_178),
.Y(n_3669)
);

NOR2xp33_ASAP7_75t_L g3670 ( 
.A(n_3486),
.B(n_180),
.Y(n_3670)
);

NAND2xp33_ASAP7_75t_SL g3671 ( 
.A(n_3441),
.B(n_181),
.Y(n_3671)
);

AO221x2_ASAP7_75t_L g3672 ( 
.A1(n_3389),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.C(n_184),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3385),
.B(n_182),
.Y(n_3673)
);

NAND2xp33_ASAP7_75t_SL g3674 ( 
.A(n_3445),
.B(n_183),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3382),
.Y(n_3675)
);

NOR2x1p5_ASAP7_75t_L g3676 ( 
.A(n_3489),
.B(n_1360),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3442),
.B(n_185),
.Y(n_3677)
);

AOI22xp5_ASAP7_75t_L g3678 ( 
.A1(n_3456),
.A2(n_1365),
.B1(n_1368),
.B2(n_1364),
.Y(n_3678)
);

OAI221xp5_ASAP7_75t_L g3679 ( 
.A1(n_3451),
.A2(n_3492),
.B1(n_3485),
.B2(n_3483),
.C(n_3477),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3397),
.B(n_185),
.Y(n_3680)
);

NAND2xp33_ASAP7_75t_SL g3681 ( 
.A(n_3446),
.B(n_187),
.Y(n_3681)
);

NOR2xp33_ASAP7_75t_SL g3682 ( 
.A(n_3370),
.B(n_1370),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3409),
.B(n_188),
.Y(n_3683)
);

AO221x2_ASAP7_75t_L g3684 ( 
.A1(n_3422),
.A2(n_3447),
.B1(n_3448),
.B2(n_3428),
.C(n_3399),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3379),
.B(n_188),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3383),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3463),
.B(n_189),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3386),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3465),
.B(n_190),
.Y(n_3689)
);

NOR2x1_ASAP7_75t_L g3690 ( 
.A(n_3510),
.B(n_191),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3461),
.B(n_192),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_R g3692 ( 
.A(n_3450),
.B(n_192),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3620),
.B(n_3610),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_3642),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3575),
.B(n_3624),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3565),
.Y(n_3696)
);

AND2x2_ASAP7_75t_L g3697 ( 
.A(n_3567),
.B(n_3476),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3628),
.Y(n_3698)
);

AOI22xp5_ASAP7_75t_L g3699 ( 
.A1(n_3598),
.A2(n_3391),
.B1(n_3392),
.B2(n_3388),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3606),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_SL g3701 ( 
.A(n_3577),
.B(n_3473),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3579),
.Y(n_3702)
);

OR2x2_ASAP7_75t_L g3703 ( 
.A(n_3618),
.B(n_3396),
.Y(n_3703)
);

INVx2_ASAP7_75t_SL g3704 ( 
.A(n_3559),
.Y(n_3704)
);

O2A1O1Ixp33_ASAP7_75t_L g3705 ( 
.A1(n_3563),
.A2(n_3504),
.B(n_3404),
.C(n_3407),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3658),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3616),
.B(n_3634),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3677),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3635),
.B(n_3405),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3652),
.B(n_3410),
.Y(n_3710)
);

O2A1O1Ixp33_ASAP7_75t_L g3711 ( 
.A1(n_3561),
.A2(n_3418),
.B(n_3419),
.C(n_3412),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3665),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3686),
.Y(n_3713)
);

AND2x4_ASAP7_75t_L g3714 ( 
.A(n_3611),
.B(n_3496),
.Y(n_3714)
);

INVxp67_ASAP7_75t_L g3715 ( 
.A(n_3570),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3676),
.B(n_3653),
.Y(n_3716)
);

OR2x2_ASAP7_75t_L g3717 ( 
.A(n_3663),
.B(n_3576),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3599),
.Y(n_3718)
);

HB1xp67_ASAP7_75t_L g3719 ( 
.A(n_3690),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3639),
.Y(n_3720)
);

AND2x4_ASAP7_75t_L g3721 ( 
.A(n_3568),
.B(n_3499),
.Y(n_3721)
);

NAND2x1_ASAP7_75t_L g3722 ( 
.A(n_3622),
.B(n_3623),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3627),
.B(n_3452),
.Y(n_3723)
);

NOR2xp33_ASAP7_75t_L g3724 ( 
.A(n_3626),
.B(n_3506),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3650),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3664),
.Y(n_3726)
);

INVx1_ASAP7_75t_SL g3727 ( 
.A(n_3573),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3564),
.B(n_3421),
.Y(n_3728)
);

AOI21xp33_ASAP7_75t_SL g3729 ( 
.A1(n_3587),
.A2(n_3458),
.B(n_3457),
.Y(n_3729)
);

NOR2xp67_ASAP7_75t_L g3730 ( 
.A(n_3571),
.B(n_3425),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3675),
.Y(n_3731)
);

OR2x2_ASAP7_75t_L g3732 ( 
.A(n_3619),
.B(n_3429),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3688),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3609),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3602),
.Y(n_3735)
);

AND2x4_ASAP7_75t_L g3736 ( 
.A(n_3607),
.B(n_3500),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3564),
.B(n_3432),
.Y(n_3737)
);

AOI21xp33_ASAP7_75t_SL g3738 ( 
.A1(n_3625),
.A2(n_3637),
.B(n_3617),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3684),
.B(n_3434),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3651),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3603),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3584),
.A2(n_3668),
.B(n_3621),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3597),
.B(n_3435),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3654),
.Y(n_3744)
);

NOR2xp67_ASAP7_75t_L g3745 ( 
.A(n_3562),
.B(n_3581),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3600),
.Y(n_3746)
);

XOR2x2_ASAP7_75t_L g3747 ( 
.A(n_3679),
.B(n_3459),
.Y(n_3747)
);

AOI222xp33_ASAP7_75t_L g3748 ( 
.A1(n_3669),
.A2(n_3472),
.B1(n_3454),
.B2(n_3440),
.C1(n_3449),
.C2(n_3439),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3670),
.B(n_3692),
.Y(n_3749)
);

INVx1_ASAP7_75t_SL g3750 ( 
.A(n_3593),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3629),
.B(n_3517),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3632),
.B(n_3521),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3615),
.B(n_3530),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3601),
.B(n_3479),
.Y(n_3754)
);

INVxp67_ASAP7_75t_L g3755 ( 
.A(n_3644),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3667),
.B(n_3533),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3580),
.Y(n_3757)
);

INVx1_ASAP7_75t_SL g3758 ( 
.A(n_3647),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3572),
.Y(n_3759)
);

AOI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_3566),
.A2(n_3541),
.B1(n_3551),
.B2(n_3534),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3645),
.B(n_3552),
.Y(n_3761)
);

AND2x4_ASAP7_75t_L g3762 ( 
.A(n_3649),
.B(n_3548),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3578),
.Y(n_3763)
);

OR2x2_ASAP7_75t_L g3764 ( 
.A(n_3574),
.B(n_193),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3687),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3615),
.B(n_193),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3691),
.B(n_194),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3582),
.B(n_3589),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3689),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3569),
.B(n_194),
.Y(n_3770)
);

NOR2x1_ASAP7_75t_L g3771 ( 
.A(n_3586),
.B(n_3560),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3659),
.B(n_195),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3660),
.B(n_195),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3646),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3588),
.B(n_197),
.Y(n_3775)
);

INVx2_ASAP7_75t_SL g3776 ( 
.A(n_3631),
.Y(n_3776)
);

NAND2x1p5_ASAP7_75t_L g3777 ( 
.A(n_3583),
.B(n_200),
.Y(n_3777)
);

INVxp67_ASAP7_75t_L g3778 ( 
.A(n_3671),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3661),
.B(n_199),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3613),
.B(n_3605),
.Y(n_3780)
);

OR2x2_ASAP7_75t_L g3781 ( 
.A(n_3655),
.B(n_199),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3742),
.A2(n_3701),
.B(n_3719),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3717),
.Y(n_3783)
);

OAI332xp33_ASAP7_75t_L g3784 ( 
.A1(n_3776),
.A2(n_3630),
.A3(n_3638),
.B1(n_3643),
.B2(n_3673),
.B3(n_3633),
.C1(n_3685),
.C2(n_3683),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3695),
.B(n_3662),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3704),
.Y(n_3786)
);

NOR2x1p5_ASAP7_75t_L g3787 ( 
.A(n_3722),
.B(n_3657),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3758),
.B(n_3631),
.Y(n_3788)
);

INVxp67_ASAP7_75t_L g3789 ( 
.A(n_3736),
.Y(n_3789)
);

AND2x2_ASAP7_75t_L g3790 ( 
.A(n_3750),
.B(n_3640),
.Y(n_3790)
);

AOI32xp33_ASAP7_75t_L g3791 ( 
.A1(n_3780),
.A2(n_3674),
.A3(n_3681),
.B1(n_3666),
.B2(n_3614),
.Y(n_3791)
);

NOR2x1_ASAP7_75t_L g3792 ( 
.A(n_3707),
.B(n_3766),
.Y(n_3792)
);

OAI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3694),
.A2(n_3699),
.B1(n_3730),
.B2(n_3778),
.Y(n_3793)
);

OAI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_3755),
.A2(n_3594),
.B(n_3636),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3723),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3744),
.B(n_3595),
.Y(n_3796)
);

INVx2_ASAP7_75t_SL g3797 ( 
.A(n_3702),
.Y(n_3797)
);

OAI22xp33_ASAP7_75t_L g3798 ( 
.A1(n_3753),
.A2(n_3608),
.B1(n_3682),
.B2(n_3596),
.Y(n_3798)
);

AOI21xp33_ASAP7_75t_L g3799 ( 
.A1(n_3693),
.A2(n_3648),
.B(n_3592),
.Y(n_3799)
);

OAI222xp33_ASAP7_75t_L g3800 ( 
.A1(n_3728),
.A2(n_3680),
.B1(n_3678),
.B2(n_3656),
.C1(n_3672),
.C2(n_3585),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3700),
.B(n_3672),
.Y(n_3801)
);

XNOR2x1_ASAP7_75t_L g3802 ( 
.A(n_3747),
.B(n_3612),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3697),
.B(n_3595),
.Y(n_3803)
);

INVxp67_ASAP7_75t_L g3804 ( 
.A(n_3749),
.Y(n_3804)
);

INVx2_ASAP7_75t_SL g3805 ( 
.A(n_3714),
.Y(n_3805)
);

AOI221xp5_ASAP7_75t_L g3806 ( 
.A1(n_3739),
.A2(n_3737),
.B1(n_3696),
.B2(n_3729),
.C(n_3711),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3703),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3781),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3756),
.Y(n_3809)
);

AOI221xp5_ASAP7_75t_L g3810 ( 
.A1(n_3698),
.A2(n_3590),
.B1(n_3591),
.B2(n_3604),
.C(n_3585),
.Y(n_3810)
);

OAI221xp5_ASAP7_75t_L g3811 ( 
.A1(n_3760),
.A2(n_3709),
.B1(n_3710),
.B2(n_3706),
.C(n_3751),
.Y(n_3811)
);

OAI221xp5_ASAP7_75t_L g3812 ( 
.A1(n_3752),
.A2(n_3641),
.B1(n_1454),
.B2(n_1527),
.C(n_1418),
.Y(n_3812)
);

BUFx2_ASAP7_75t_L g3813 ( 
.A(n_3715),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3761),
.Y(n_3814)
);

AOI221xp5_ASAP7_75t_L g3815 ( 
.A1(n_3735),
.A2(n_1385),
.B1(n_1394),
.B2(n_1376),
.C(n_1373),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3727),
.B(n_200),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3740),
.B(n_201),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3768),
.A2(n_1409),
.B(n_1395),
.Y(n_3818)
);

AOI21xp33_ASAP7_75t_L g3819 ( 
.A1(n_3705),
.A2(n_201),
.B(n_204),
.Y(n_3819)
);

INVx1_ASAP7_75t_SL g3820 ( 
.A(n_3716),
.Y(n_3820)
);

NOR3xp33_ASAP7_75t_L g3821 ( 
.A(n_3708),
.B(n_3746),
.C(n_3741),
.Y(n_3821)
);

AND2x4_ASAP7_75t_L g3822 ( 
.A(n_3721),
.B(n_205),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3712),
.Y(n_3823)
);

OAI221xp5_ASAP7_75t_L g3824 ( 
.A1(n_3734),
.A2(n_1425),
.B1(n_1576),
.B2(n_1545),
.C(n_1473),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3754),
.B(n_204),
.Y(n_3825)
);

AOI22xp5_ASAP7_75t_L g3826 ( 
.A1(n_3724),
.A2(n_1411),
.B1(n_1427),
.B2(n_1410),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3743),
.B(n_205),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3762),
.B(n_206),
.Y(n_3828)
);

AOI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3745),
.A2(n_1438),
.B1(n_1439),
.B2(n_1435),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3767),
.Y(n_3830)
);

HB1xp67_ASAP7_75t_L g3831 ( 
.A(n_3777),
.Y(n_3831)
);

O2A1O1Ixp5_ASAP7_75t_L g3832 ( 
.A1(n_3713),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_3832)
);

INVx1_ASAP7_75t_SL g3833 ( 
.A(n_3770),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3774),
.B(n_207),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3775),
.A2(n_1449),
.B(n_1448),
.Y(n_3835)
);

OR2x2_ASAP7_75t_L g3836 ( 
.A(n_3788),
.B(n_3732),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3795),
.Y(n_3837)
);

AOI221xp5_ASAP7_75t_L g3838 ( 
.A1(n_3806),
.A2(n_3738),
.B1(n_3725),
.B2(n_3726),
.C(n_3720),
.Y(n_3838)
);

AND2x2_ASAP7_75t_L g3839 ( 
.A(n_3786),
.B(n_3789),
.Y(n_3839)
);

INVx1_ASAP7_75t_SL g3840 ( 
.A(n_3820),
.Y(n_3840)
);

OAI22xp5_ASAP7_75t_L g3841 ( 
.A1(n_3802),
.A2(n_3765),
.B1(n_3769),
.B2(n_3771),
.Y(n_3841)
);

AOI22xp5_ASAP7_75t_L g3842 ( 
.A1(n_3793),
.A2(n_3757),
.B1(n_3759),
.B2(n_3763),
.Y(n_3842)
);

O2A1O1Ixp5_ASAP7_75t_L g3843 ( 
.A1(n_3782),
.A2(n_3731),
.B(n_3733),
.C(n_3718),
.Y(n_3843)
);

INVx2_ASAP7_75t_SL g3844 ( 
.A(n_3787),
.Y(n_3844)
);

AOI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3805),
.A2(n_3748),
.B1(n_3773),
.B2(n_3772),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3816),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_SL g3847 ( 
.A(n_3791),
.B(n_3779),
.Y(n_3847)
);

A2O1A1Ixp33_ASAP7_75t_L g3848 ( 
.A1(n_3832),
.A2(n_3764),
.B(n_1476),
.C(n_1481),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3803),
.B(n_209),
.Y(n_3849)
);

INVxp67_ASAP7_75t_L g3850 ( 
.A(n_3796),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_3813),
.B(n_1455),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3801),
.B(n_210),
.Y(n_3852)
);

OAI22xp33_ASAP7_75t_L g3853 ( 
.A1(n_3811),
.A2(n_1503),
.B1(n_1507),
.B2(n_1499),
.Y(n_3853)
);

AOI221xp5_ASAP7_75t_L g3854 ( 
.A1(n_3800),
.A2(n_1771),
.B1(n_1546),
.B2(n_1554),
.C(n_1542),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3797),
.B(n_211),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3785),
.B(n_211),
.Y(n_3856)
);

INVx1_ASAP7_75t_SL g3857 ( 
.A(n_3822),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3804),
.Y(n_3858)
);

OR2x2_ASAP7_75t_L g3859 ( 
.A(n_3833),
.B(n_212),
.Y(n_3859)
);

OR2x2_ASAP7_75t_L g3860 ( 
.A(n_3783),
.B(n_3807),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3825),
.Y(n_3861)
);

INVxp33_ASAP7_75t_L g3862 ( 
.A(n_3792),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3831),
.B(n_212),
.Y(n_3863)
);

OAI31xp33_ASAP7_75t_L g3864 ( 
.A1(n_3798),
.A2(n_215),
.A3(n_213),
.B(n_214),
.Y(n_3864)
);

NOR2xp33_ASAP7_75t_L g3865 ( 
.A(n_3784),
.B(n_214),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3817),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3790),
.B(n_3830),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3822),
.B(n_216),
.Y(n_3868)
);

AOI22xp33_ASAP7_75t_L g3869 ( 
.A1(n_3809),
.A2(n_3814),
.B1(n_3808),
.B2(n_3821),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3823),
.B(n_216),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3827),
.B(n_218),
.Y(n_3871)
);

NAND2x1_ASAP7_75t_L g3872 ( 
.A(n_3834),
.B(n_218),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3828),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3829),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3794),
.B(n_219),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3857),
.B(n_3840),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3867),
.Y(n_3877)
);

AOI221xp5_ASAP7_75t_L g3878 ( 
.A1(n_3862),
.A2(n_3819),
.B1(n_3799),
.B2(n_3810),
.C(n_3818),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3839),
.B(n_3835),
.Y(n_3879)
);

CKINVDCx16_ASAP7_75t_R g3880 ( 
.A(n_3841),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3856),
.Y(n_3881)
);

O2A1O1Ixp5_ASAP7_75t_L g3882 ( 
.A1(n_3847),
.A2(n_3812),
.B(n_3824),
.C(n_3815),
.Y(n_3882)
);

OAI21x1_ASAP7_75t_SL g3883 ( 
.A1(n_3844),
.A2(n_3826),
.B(n_219),
.Y(n_3883)
);

AOI221xp5_ASAP7_75t_L g3884 ( 
.A1(n_3838),
.A2(n_1559),
.B1(n_1562),
.B2(n_1556),
.C(n_1536),
.Y(n_3884)
);

AOI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3865),
.A2(n_1574),
.B(n_1571),
.Y(n_3885)
);

OAI322xp33_ASAP7_75t_SL g3886 ( 
.A1(n_3858),
.A2(n_225),
.A3(n_224),
.B1(n_222),
.B2(n_220),
.C1(n_221),
.C2(n_223),
.Y(n_3886)
);

AOI22xp5_ASAP7_75t_L g3887 ( 
.A1(n_3875),
.A2(n_1591),
.B1(n_1594),
.B2(n_1583),
.Y(n_3887)
);

INVx1_ASAP7_75t_SL g3888 ( 
.A(n_3872),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3863),
.Y(n_3889)
);

INVx3_ASAP7_75t_L g3890 ( 
.A(n_3860),
.Y(n_3890)
);

AO221x1_ASAP7_75t_L g3891 ( 
.A1(n_3853),
.A2(n_223),
.B1(n_220),
.B2(n_222),
.C(n_224),
.Y(n_3891)
);

OAI22xp5_ASAP7_75t_L g3892 ( 
.A1(n_3845),
.A2(n_1599),
.B1(n_1603),
.B2(n_1595),
.Y(n_3892)
);

OAI21xp5_ASAP7_75t_SL g3893 ( 
.A1(n_3850),
.A2(n_225),
.B(n_226),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3846),
.Y(n_3894)
);

OAI211xp5_ASAP7_75t_SL g3895 ( 
.A1(n_3842),
.A2(n_228),
.B(n_226),
.C(n_227),
.Y(n_3895)
);

AOI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_3849),
.A2(n_1615),
.B(n_1614),
.Y(n_3896)
);

AOI221x1_ASAP7_75t_L g3897 ( 
.A1(n_3837),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.C(n_232),
.Y(n_3897)
);

INVx2_ASAP7_75t_SL g3898 ( 
.A(n_3870),
.Y(n_3898)
);

OAI21xp33_ASAP7_75t_L g3899 ( 
.A1(n_3869),
.A2(n_1639),
.B(n_1620),
.Y(n_3899)
);

AND2x2_ASAP7_75t_L g3900 ( 
.A(n_3852),
.B(n_229),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3871),
.Y(n_3901)
);

OR2x2_ASAP7_75t_L g3902 ( 
.A(n_3836),
.B(n_230),
.Y(n_3902)
);

AOI222xp33_ASAP7_75t_L g3903 ( 
.A1(n_3861),
.A2(n_1657),
.B1(n_1648),
.B2(n_1665),
.C1(n_1650),
.C2(n_1644),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3859),
.Y(n_3904)
);

OR2x2_ASAP7_75t_L g3905 ( 
.A(n_3855),
.B(n_233),
.Y(n_3905)
);

AND2x2_ASAP7_75t_L g3906 ( 
.A(n_3873),
.B(n_234),
.Y(n_3906)
);

AOI22xp5_ASAP7_75t_L g3907 ( 
.A1(n_3874),
.A2(n_1687),
.B1(n_1695),
.B2(n_1683),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3848),
.A2(n_1728),
.B(n_1710),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3868),
.Y(n_3909)
);

O2A1O1Ixp5_ASAP7_75t_L g3910 ( 
.A1(n_3843),
.A2(n_3866),
.B(n_3851),
.C(n_3864),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3854),
.A2(n_1754),
.B1(n_1755),
.B2(n_1742),
.Y(n_3911)
);

AOI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3865),
.A2(n_1767),
.B1(n_236),
.B2(n_234),
.Y(n_3912)
);

XNOR2x1_ASAP7_75t_L g3913 ( 
.A(n_3840),
.B(n_235),
.Y(n_3913)
);

OAI222xp33_ASAP7_75t_L g3914 ( 
.A1(n_3840),
.A2(n_237),
.B1(n_240),
.B2(n_235),
.C1(n_236),
.C2(n_238),
.Y(n_3914)
);

AOI211xp5_ASAP7_75t_SL g3915 ( 
.A1(n_3853),
.A2(n_249),
.B(n_259),
.C(n_237),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3857),
.B(n_240),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3890),
.Y(n_3917)
);

INVxp33_ASAP7_75t_SL g3918 ( 
.A(n_3876),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3890),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3877),
.Y(n_3920)
);

NOR2xp33_ASAP7_75t_L g3921 ( 
.A(n_3888),
.B(n_243),
.Y(n_3921)
);

NOR2xp33_ASAP7_75t_L g3922 ( 
.A(n_3880),
.B(n_244),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3900),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3916),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3889),
.Y(n_3925)
);

HB1xp67_ASAP7_75t_L g3926 ( 
.A(n_3913),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3881),
.Y(n_3927)
);

BUFx2_ASAP7_75t_L g3928 ( 
.A(n_3898),
.Y(n_3928)
);

NOR2xp33_ASAP7_75t_L g3929 ( 
.A(n_3893),
.B(n_245),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3902),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3906),
.Y(n_3931)
);

HB1xp67_ASAP7_75t_L g3932 ( 
.A(n_3904),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3905),
.Y(n_3933)
);

INVx8_ASAP7_75t_L g3934 ( 
.A(n_3894),
.Y(n_3934)
);

INVx1_ASAP7_75t_SL g3935 ( 
.A(n_3901),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3909),
.Y(n_3936)
);

INVx1_ASAP7_75t_SL g3937 ( 
.A(n_3879),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3897),
.Y(n_3938)
);

INVxp67_ASAP7_75t_L g3939 ( 
.A(n_3883),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3891),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3910),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3895),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3907),
.Y(n_3943)
);

INVxp33_ASAP7_75t_L g3944 ( 
.A(n_3878),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3912),
.Y(n_3945)
);

INVx2_ASAP7_75t_L g3946 ( 
.A(n_3882),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3915),
.B(n_245),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3887),
.Y(n_3948)
);

CKINVDCx5p33_ASAP7_75t_R g3949 ( 
.A(n_3892),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3899),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3896),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3885),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3911),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3903),
.Y(n_3954)
);

CKINVDCx5p33_ASAP7_75t_R g3955 ( 
.A(n_3886),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3914),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3908),
.Y(n_3957)
);

BUFx4_ASAP7_75t_SL g3958 ( 
.A(n_3884),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3890),
.Y(n_3959)
);

INVx3_ASAP7_75t_L g3960 ( 
.A(n_3890),
.Y(n_3960)
);

BUFx2_ASAP7_75t_L g3961 ( 
.A(n_3890),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3890),
.Y(n_3962)
);

BUFx2_ASAP7_75t_L g3963 ( 
.A(n_3890),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3890),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3890),
.Y(n_3965)
);

INVxp33_ASAP7_75t_L g3966 ( 
.A(n_3913),
.Y(n_3966)
);

NOR2xp67_ASAP7_75t_L g3967 ( 
.A(n_3960),
.B(n_246),
.Y(n_3967)
);

NAND4xp25_ASAP7_75t_L g3968 ( 
.A(n_3918),
.B(n_248),
.C(n_246),
.D(n_247),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3961),
.B(n_3963),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3926),
.B(n_247),
.Y(n_3970)
);

NOR2xp33_ASAP7_75t_L g3971 ( 
.A(n_3966),
.B(n_250),
.Y(n_3971)
);

NOR3xp33_ASAP7_75t_L g3972 ( 
.A(n_3941),
.B(n_260),
.C(n_250),
.Y(n_3972)
);

NAND5xp2_ASAP7_75t_L g3973 ( 
.A(n_3944),
.B(n_254),
.C(n_251),
.D(n_252),
.E(n_256),
.Y(n_3973)
);

OR2x2_ASAP7_75t_L g3974 ( 
.A(n_3956),
.B(n_251),
.Y(n_3974)
);

NOR2x1_ASAP7_75t_L g3975 ( 
.A(n_3917),
.B(n_252),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3928),
.B(n_256),
.Y(n_3976)
);

NOR3xp33_ASAP7_75t_L g3977 ( 
.A(n_3939),
.B(n_266),
.C(n_257),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_3922),
.A2(n_3935),
.B(n_3919),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3959),
.B(n_3962),
.Y(n_3979)
);

AOI21xp5_ASAP7_75t_L g3980 ( 
.A1(n_3964),
.A2(n_257),
.B(n_258),
.Y(n_3980)
);

OAI211xp5_ASAP7_75t_SL g3981 ( 
.A1(n_3937),
.A2(n_261),
.B(n_258),
.C(n_259),
.Y(n_3981)
);

OAI21xp33_ASAP7_75t_L g3982 ( 
.A1(n_3955),
.A2(n_270),
.B(n_261),
.Y(n_3982)
);

NOR2x1_ASAP7_75t_L g3983 ( 
.A(n_3965),
.B(n_262),
.Y(n_3983)
);

NOR2xp33_ASAP7_75t_L g3984 ( 
.A(n_3938),
.B(n_262),
.Y(n_3984)
);

NOR2x1_ASAP7_75t_L g3985 ( 
.A(n_3946),
.B(n_263),
.Y(n_3985)
);

NOR2xp33_ASAP7_75t_L g3986 ( 
.A(n_3942),
.B(n_3940),
.Y(n_3986)
);

NAND4xp25_ASAP7_75t_L g3987 ( 
.A(n_3945),
.B(n_265),
.C(n_263),
.D(n_264),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3934),
.B(n_266),
.Y(n_3988)
);

OAI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_3921),
.A2(n_268),
.B(n_269),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3934),
.B(n_268),
.Y(n_3990)
);

NOR2xp33_ASAP7_75t_SL g3991 ( 
.A(n_3932),
.B(n_269),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_L g3992 ( 
.A(n_3923),
.B(n_270),
.Y(n_3992)
);

INVx1_ASAP7_75t_SL g3993 ( 
.A(n_3947),
.Y(n_3993)
);

AOI211x1_ASAP7_75t_L g3994 ( 
.A1(n_3920),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_3994)
);

AOI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3930),
.A2(n_271),
.B(n_272),
.Y(n_3995)
);

NOR2xp33_ASAP7_75t_L g3996 ( 
.A(n_3931),
.B(n_273),
.Y(n_3996)
);

OA22x2_ASAP7_75t_L g3997 ( 
.A1(n_3927),
.A2(n_276),
.B1(n_277),
.B2(n_275),
.Y(n_3997)
);

NOR2xp33_ASAP7_75t_L g3998 ( 
.A(n_3925),
.B(n_274),
.Y(n_3998)
);

NOR2xp33_ASAP7_75t_L g3999 ( 
.A(n_3929),
.B(n_276),
.Y(n_3999)
);

NAND4xp25_ASAP7_75t_L g4000 ( 
.A(n_3924),
.B(n_280),
.C(n_277),
.D(n_279),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3933),
.B(n_279),
.Y(n_4001)
);

XNOR2x2_ASAP7_75t_L g4002 ( 
.A(n_3936),
.B(n_281),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3954),
.B(n_281),
.Y(n_4003)
);

NOR3xp33_ASAP7_75t_SL g4004 ( 
.A(n_3949),
.B(n_283),
.C(n_284),
.Y(n_4004)
);

OAI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3952),
.A2(n_283),
.B(n_284),
.Y(n_4005)
);

OAI322xp33_ASAP7_75t_L g4006 ( 
.A1(n_3957),
.A2(n_290),
.A3(n_289),
.B1(n_287),
.B2(n_285),
.C1(n_286),
.C2(n_288),
.Y(n_4006)
);

NOR2xp33_ASAP7_75t_L g4007 ( 
.A(n_3951),
.B(n_285),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3950),
.Y(n_4008)
);

NOR2x1p5_ASAP7_75t_SL g4009 ( 
.A(n_3953),
.B(n_286),
.Y(n_4009)
);

NOR2x1_ASAP7_75t_L g4010 ( 
.A(n_3943),
.B(n_289),
.Y(n_4010)
);

AOI211xp5_ASAP7_75t_L g4011 ( 
.A1(n_3948),
.A2(n_293),
.B(n_291),
.C(n_292),
.Y(n_4011)
);

HB1xp67_ASAP7_75t_L g4012 ( 
.A(n_3958),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3961),
.Y(n_4013)
);

NOR2x1_ASAP7_75t_L g4014 ( 
.A(n_3961),
.B(n_293),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3961),
.Y(n_4015)
);

NOR3xp33_ASAP7_75t_L g4016 ( 
.A(n_3960),
.B(n_305),
.C(n_294),
.Y(n_4016)
);

INVx2_ASAP7_75t_SL g4017 ( 
.A(n_3961),
.Y(n_4017)
);

NOR2x1_ASAP7_75t_L g4018 ( 
.A(n_3961),
.B(n_295),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3961),
.Y(n_4019)
);

NAND3xp33_ASAP7_75t_L g4020 ( 
.A(n_3941),
.B(n_295),
.C(n_296),
.Y(n_4020)
);

NOR2xp33_ASAP7_75t_L g4021 ( 
.A(n_3966),
.B(n_296),
.Y(n_4021)
);

AND4x1_ASAP7_75t_L g4022 ( 
.A(n_3922),
.B(n_301),
.C(n_298),
.D(n_299),
.Y(n_4022)
);

NOR3xp33_ASAP7_75t_L g4023 ( 
.A(n_3960),
.B(n_312),
.C(n_299),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3961),
.B(n_302),
.Y(n_4024)
);

NOR2x1p5_ASAP7_75t_L g4025 ( 
.A(n_3960),
.B(n_305),
.Y(n_4025)
);

NOR3xp33_ASAP7_75t_L g4026 ( 
.A(n_3960),
.B(n_316),
.C(n_304),
.Y(n_4026)
);

NOR2x1_ASAP7_75t_L g4027 ( 
.A(n_3961),
.B(n_306),
.Y(n_4027)
);

NOR3xp33_ASAP7_75t_L g4028 ( 
.A(n_3960),
.B(n_317),
.C(n_306),
.Y(n_4028)
);

NOR2xp67_ASAP7_75t_SL g4029 ( 
.A(n_3960),
.B(n_308),
.Y(n_4029)
);

NOR3x1_ASAP7_75t_L g4030 ( 
.A(n_3961),
.B(n_310),
.C(n_311),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3961),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3961),
.B(n_310),
.Y(n_4032)
);

NOR2xp33_ASAP7_75t_L g4033 ( 
.A(n_3966),
.B(n_311),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3941),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_4034)
);

NOR3xp33_ASAP7_75t_L g4035 ( 
.A(n_3960),
.B(n_323),
.C(n_314),
.Y(n_4035)
);

NOR2xp33_ASAP7_75t_L g4036 ( 
.A(n_3966),
.B(n_316),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3961),
.B(n_317),
.Y(n_4037)
);

OAI21xp33_ASAP7_75t_L g4038 ( 
.A1(n_3966),
.A2(n_327),
.B(n_318),
.Y(n_4038)
);

NOR2xp33_ASAP7_75t_L g4039 ( 
.A(n_3966),
.B(n_318),
.Y(n_4039)
);

NOR2x1_ASAP7_75t_L g4040 ( 
.A(n_3961),
.B(n_319),
.Y(n_4040)
);

NOR3xp33_ASAP7_75t_L g4041 ( 
.A(n_3960),
.B(n_329),
.C(n_320),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3961),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3961),
.B(n_321),
.Y(n_4043)
);

NOR2x1_ASAP7_75t_SL g4044 ( 
.A(n_3917),
.B(n_322),
.Y(n_4044)
);

NOR3xp33_ASAP7_75t_SL g4045 ( 
.A(n_3955),
.B(n_322),
.C(n_324),
.Y(n_4045)
);

NOR2xp67_ASAP7_75t_L g4046 ( 
.A(n_3960),
.B(n_324),
.Y(n_4046)
);

AOI21xp5_ASAP7_75t_L g4047 ( 
.A1(n_3918),
.A2(n_325),
.B(n_326),
.Y(n_4047)
);

BUFx2_ASAP7_75t_L g4048 ( 
.A(n_3961),
.Y(n_4048)
);

NOR3xp33_ASAP7_75t_L g4049 ( 
.A(n_3960),
.B(n_336),
.C(n_326),
.Y(n_4049)
);

OAI211xp5_ASAP7_75t_SL g4050 ( 
.A1(n_3978),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_4050)
);

OAI221xp5_ASAP7_75t_L g4051 ( 
.A1(n_4017),
.A2(n_331),
.B1(n_328),
.B2(n_330),
.C(n_332),
.Y(n_4051)
);

OA211x2_ASAP7_75t_L g4052 ( 
.A1(n_3991),
.A2(n_334),
.B(n_331),
.C(n_332),
.Y(n_4052)
);

NOR2x1_ASAP7_75t_L g4053 ( 
.A(n_4048),
.B(n_337),
.Y(n_4053)
);

AOI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_3986),
.A2(n_341),
.B1(n_338),
.B2(n_339),
.Y(n_4054)
);

NAND4xp25_ASAP7_75t_SL g4055 ( 
.A(n_3969),
.B(n_342),
.C(n_338),
.D(n_339),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_4044),
.Y(n_4056)
);

AOI211xp5_ASAP7_75t_L g4057 ( 
.A1(n_4015),
.A2(n_345),
.B(n_343),
.C(n_344),
.Y(n_4057)
);

AOI221xp5_ASAP7_75t_L g4058 ( 
.A1(n_3984),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.C(n_347),
.Y(n_4058)
);

OAI21xp5_ASAP7_75t_SL g4059 ( 
.A1(n_4019),
.A2(n_347),
.B(n_348),
.Y(n_4059)
);

NOR4xp75_ASAP7_75t_SL g4060 ( 
.A(n_4034),
.B(n_351),
.C(n_349),
.D(n_350),
.Y(n_4060)
);

NAND4xp25_ASAP7_75t_L g4061 ( 
.A(n_3974),
.B(n_353),
.C(n_350),
.D(n_352),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_4014),
.Y(n_4062)
);

AOI221xp5_ASAP7_75t_L g4063 ( 
.A1(n_3972),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.C(n_355),
.Y(n_4063)
);

AND2x4_ASAP7_75t_L g4064 ( 
.A(n_3967),
.B(n_354),
.Y(n_4064)
);

AOI221xp5_ASAP7_75t_L g4065 ( 
.A1(n_4031),
.A2(n_358),
.B1(n_355),
.B2(n_356),
.C(n_359),
.Y(n_4065)
);

AO22x2_ASAP7_75t_L g4066 ( 
.A1(n_3994),
.A2(n_360),
.B1(n_356),
.B2(n_359),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_4046),
.B(n_360),
.Y(n_4067)
);

AOI221xp5_ASAP7_75t_SL g4068 ( 
.A1(n_4042),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.C(n_364),
.Y(n_4068)
);

OAI211xp5_ASAP7_75t_L g4069 ( 
.A1(n_3985),
.A2(n_370),
.B(n_381),
.C(n_361),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_4018),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_4029),
.B(n_3976),
.Y(n_4071)
);

NOR3xp33_ASAP7_75t_L g4072 ( 
.A(n_3971),
.B(n_362),
.C(n_364),
.Y(n_4072)
);

NAND3xp33_ASAP7_75t_SL g4073 ( 
.A(n_4013),
.B(n_365),
.C(n_366),
.Y(n_4073)
);

AOI211xp5_ASAP7_75t_L g4074 ( 
.A1(n_4020),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_4074)
);

NAND4xp25_ASAP7_75t_L g4075 ( 
.A(n_4008),
.B(n_369),
.C(n_367),
.D(n_368),
.Y(n_4075)
);

NAND4xp25_ASAP7_75t_L g4076 ( 
.A(n_3993),
.B(n_374),
.C(n_370),
.D(n_371),
.Y(n_4076)
);

NOR2xp33_ASAP7_75t_L g4077 ( 
.A(n_4022),
.B(n_371),
.Y(n_4077)
);

NAND4xp25_ASAP7_75t_L g4078 ( 
.A(n_3979),
.B(n_377),
.C(n_374),
.D(n_376),
.Y(n_4078)
);

NOR2x1_ASAP7_75t_L g4079 ( 
.A(n_4027),
.B(n_376),
.Y(n_4079)
);

NAND4xp25_ASAP7_75t_L g4080 ( 
.A(n_4021),
.B(n_380),
.C(n_378),
.D(n_379),
.Y(n_4080)
);

NAND3xp33_ASAP7_75t_SL g4081 ( 
.A(n_3977),
.B(n_379),
.C(n_380),
.Y(n_4081)
);

BUFx12f_ASAP7_75t_L g4082 ( 
.A(n_3970),
.Y(n_4082)
);

O2A1O1Ixp5_ASAP7_75t_L g4083 ( 
.A1(n_4024),
.A2(n_383),
.B(n_381),
.C(n_382),
.Y(n_4083)
);

OAI222xp33_ASAP7_75t_R g4084 ( 
.A1(n_4012),
.A2(n_384),
.B1(n_386),
.B2(n_382),
.C1(n_383),
.C2(n_385),
.Y(n_4084)
);

NOR2xp33_ASAP7_75t_L g4085 ( 
.A(n_3973),
.B(n_384),
.Y(n_4085)
);

NOR3xp33_ASAP7_75t_SL g4086 ( 
.A(n_3982),
.B(n_387),
.C(n_388),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_L g4087 ( 
.A(n_3968),
.B(n_387),
.Y(n_4087)
);

NOR3xp33_ASAP7_75t_L g4088 ( 
.A(n_4033),
.B(n_388),
.C(n_390),
.Y(n_4088)
);

OAI211xp5_ASAP7_75t_SL g4089 ( 
.A1(n_4045),
.A2(n_4004),
.B(n_4039),
.C(n_4036),
.Y(n_4089)
);

NAND3xp33_ASAP7_75t_L g4090 ( 
.A(n_4040),
.B(n_391),
.C(n_392),
.Y(n_4090)
);

NAND4xp25_ASAP7_75t_L g4091 ( 
.A(n_4003),
.B(n_393),
.C(n_391),
.D(n_392),
.Y(n_4091)
);

NOR2x1_ASAP7_75t_L g4092 ( 
.A(n_3975),
.B(n_393),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_4009),
.Y(n_4093)
);

OAI211xp5_ASAP7_75t_SL g4094 ( 
.A1(n_4032),
.A2(n_396),
.B(n_394),
.C(n_395),
.Y(n_4094)
);

AOI221xp5_ASAP7_75t_L g4095 ( 
.A1(n_3981),
.A2(n_397),
.B1(n_394),
.B2(n_395),
.C(n_398),
.Y(n_4095)
);

NOR2xp33_ASAP7_75t_L g4096 ( 
.A(n_3987),
.B(n_397),
.Y(n_4096)
);

OAI211xp5_ASAP7_75t_L g4097 ( 
.A1(n_4037),
.A2(n_410),
.B(n_418),
.C(n_399),
.Y(n_4097)
);

A2O1A1Ixp33_ASAP7_75t_L g4098 ( 
.A1(n_3998),
.A2(n_402),
.B(n_399),
.C(n_401),
.Y(n_4098)
);

OAI211xp5_ASAP7_75t_L g4099 ( 
.A1(n_4043),
.A2(n_413),
.B(n_421),
.C(n_401),
.Y(n_4099)
);

NAND4xp25_ASAP7_75t_L g4100 ( 
.A(n_4030),
.B(n_406),
.C(n_404),
.D(n_405),
.Y(n_4100)
);

AOI211xp5_ASAP7_75t_L g4101 ( 
.A1(n_4038),
.A2(n_406),
.B(n_404),
.C(n_405),
.Y(n_4101)
);

NAND3xp33_ASAP7_75t_SL g4102 ( 
.A(n_3988),
.B(n_407),
.C(n_408),
.Y(n_4102)
);

NAND3xp33_ASAP7_75t_SL g4103 ( 
.A(n_3990),
.B(n_407),
.C(n_411),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_4025),
.B(n_412),
.Y(n_4104)
);

OAI211xp5_ASAP7_75t_L g4105 ( 
.A1(n_4010),
.A2(n_423),
.B(n_431),
.C(n_414),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3983),
.Y(n_4106)
);

AOI22xp5_ASAP7_75t_L g4107 ( 
.A1(n_3999),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_4107)
);

NAND4xp25_ASAP7_75t_SL g4108 ( 
.A(n_3992),
.B(n_418),
.C(n_415),
.D(n_417),
.Y(n_4108)
);

AOI211x1_ASAP7_75t_L g4109 ( 
.A1(n_4047),
.A2(n_422),
.B(n_419),
.C(n_420),
.Y(n_4109)
);

NOR2x1_ASAP7_75t_L g4110 ( 
.A(n_4000),
.B(n_419),
.Y(n_4110)
);

NAND3xp33_ASAP7_75t_L g4111 ( 
.A(n_4011),
.B(n_420),
.C(n_423),
.Y(n_4111)
);

OAI211xp5_ASAP7_75t_L g4112 ( 
.A1(n_4001),
.A2(n_432),
.B(n_440),
.C(n_424),
.Y(n_4112)
);

OAI221xp5_ASAP7_75t_L g4113 ( 
.A1(n_3989),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.C(n_427),
.Y(n_4113)
);

NOR2xp67_ASAP7_75t_L g4114 ( 
.A(n_3980),
.B(n_425),
.Y(n_4114)
);

AOI211xp5_ASAP7_75t_L g4115 ( 
.A1(n_4006),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3995),
.B(n_4016),
.Y(n_4116)
);

AOI33xp33_ASAP7_75t_L g4117 ( 
.A1(n_4002),
.A2(n_431),
.A3(n_434),
.B1(n_429),
.B2(n_430),
.B3(n_433),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3997),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3996),
.Y(n_4119)
);

AOI211x1_ASAP7_75t_SL g4120 ( 
.A1(n_4005),
.A2(n_434),
.B(n_429),
.C(n_430),
.Y(n_4120)
);

NOR2x1_ASAP7_75t_L g4121 ( 
.A(n_4007),
.B(n_435),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4023),
.Y(n_4122)
);

NAND2x1p5_ASAP7_75t_L g4123 ( 
.A(n_4026),
.B(n_436),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_4028),
.B(n_435),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_4035),
.B(n_436),
.Y(n_4125)
);

NOR3xp33_ASAP7_75t_L g4126 ( 
.A(n_4041),
.B(n_4049),
.C(n_437),
.Y(n_4126)
);

NOR3x1_ASAP7_75t_L g4127 ( 
.A(n_4048),
.B(n_439),
.C(n_438),
.Y(n_4127)
);

NOR4xp25_ASAP7_75t_SL g4128 ( 
.A(n_4048),
.B(n_440),
.C(n_437),
.D(n_438),
.Y(n_4128)
);

NAND2x1p5_ASAP7_75t_L g4129 ( 
.A(n_4048),
.B(n_442),
.Y(n_4129)
);

NOR3xp33_ASAP7_75t_L g4130 ( 
.A(n_3969),
.B(n_441),
.C(n_443),
.Y(n_4130)
);

OAI221xp5_ASAP7_75t_L g4131 ( 
.A1(n_4017),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.C(n_447),
.Y(n_4131)
);

NOR3xp33_ASAP7_75t_SL g4132 ( 
.A(n_3969),
.B(n_444),
.C(n_445),
.Y(n_4132)
);

NOR2xp33_ASAP7_75t_L g4133 ( 
.A(n_4056),
.B(n_446),
.Y(n_4133)
);

OR2x2_ASAP7_75t_L g4134 ( 
.A(n_4093),
.B(n_448),
.Y(n_4134)
);

AOI211xp5_ASAP7_75t_L g4135 ( 
.A1(n_4089),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_4135)
);

NOR2x1_ASAP7_75t_L g4136 ( 
.A(n_4079),
.B(n_449),
.Y(n_4136)
);

AOI221xp5_ASAP7_75t_L g4137 ( 
.A1(n_4118),
.A2(n_453),
.B1(n_450),
.B2(n_451),
.C(n_454),
.Y(n_4137)
);

NOR2x1_ASAP7_75t_L g4138 ( 
.A(n_4053),
.B(n_455),
.Y(n_4138)
);

NOR5xp2_ASAP7_75t_L g4139 ( 
.A(n_4050),
.B(n_457),
.C(n_455),
.D(n_456),
.E(n_458),
.Y(n_4139)
);

OAI211xp5_ASAP7_75t_SL g4140 ( 
.A1(n_4071),
.A2(n_459),
.B(n_456),
.C(n_457),
.Y(n_4140)
);

NOR2x2_ASAP7_75t_L g4141 ( 
.A(n_4119),
.B(n_459),
.Y(n_4141)
);

NOR3xp33_ASAP7_75t_L g4142 ( 
.A(n_4081),
.B(n_462),
.C(n_461),
.Y(n_4142)
);

AOI221xp5_ASAP7_75t_L g4143 ( 
.A1(n_4062),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.C(n_463),
.Y(n_4143)
);

AOI221xp5_ASAP7_75t_SL g4144 ( 
.A1(n_4070),
.A2(n_4106),
.B1(n_4115),
.B2(n_4122),
.C(n_4116),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4064),
.Y(n_4145)
);

AND4x1_ASAP7_75t_L g4146 ( 
.A(n_4127),
.B(n_4117),
.C(n_4132),
.D(n_4077),
.Y(n_4146)
);

NAND4xp25_ASAP7_75t_SL g4147 ( 
.A(n_4126),
.B(n_464),
.C(n_460),
.D(n_463),
.Y(n_4147)
);

OAI221xp5_ASAP7_75t_L g4148 ( 
.A1(n_4059),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.C(n_467),
.Y(n_4148)
);

NOR2xp33_ASAP7_75t_L g4149 ( 
.A(n_4100),
.B(n_465),
.Y(n_4149)
);

NOR4xp25_ASAP7_75t_L g4150 ( 
.A(n_4069),
.B(n_469),
.C(n_466),
.D(n_468),
.Y(n_4150)
);

NOR2xp33_ASAP7_75t_L g4151 ( 
.A(n_4061),
.B(n_468),
.Y(n_4151)
);

NAND3xp33_ASAP7_75t_SL g4152 ( 
.A(n_4128),
.B(n_469),
.C(n_472),
.Y(n_4152)
);

AOI211xp5_ASAP7_75t_L g4153 ( 
.A1(n_4111),
.A2(n_474),
.B(n_472),
.C(n_473),
.Y(n_4153)
);

AOI211xp5_ASAP7_75t_L g4154 ( 
.A1(n_4114),
.A2(n_475),
.B(n_473),
.C(n_474),
.Y(n_4154)
);

OAI221xp5_ASAP7_75t_L g4155 ( 
.A1(n_4129),
.A2(n_479),
.B1(n_475),
.B2(n_477),
.C(n_480),
.Y(n_4155)
);

OAI321xp33_ASAP7_75t_L g4156 ( 
.A1(n_4123),
.A2(n_480),
.A3(n_483),
.B1(n_477),
.B2(n_479),
.C(n_482),
.Y(n_4156)
);

NOR3xp33_ASAP7_75t_L g4157 ( 
.A(n_4073),
.B(n_485),
.C(n_484),
.Y(n_4157)
);

NOR3xp33_ASAP7_75t_SL g4158 ( 
.A(n_4102),
.B(n_4103),
.C(n_4113),
.Y(n_4158)
);

NAND5xp2_ASAP7_75t_L g4159 ( 
.A(n_4095),
.B(n_486),
.C(n_482),
.D(n_485),
.E(n_487),
.Y(n_4159)
);

OAI211xp5_ASAP7_75t_SL g4160 ( 
.A1(n_4110),
.A2(n_489),
.B(n_486),
.C(n_488),
.Y(n_4160)
);

OAI321xp33_ASAP7_75t_L g4161 ( 
.A1(n_4094),
.A2(n_491),
.A3(n_494),
.B1(n_488),
.B2(n_490),
.C(n_492),
.Y(n_4161)
);

NAND3xp33_ASAP7_75t_SL g4162 ( 
.A(n_4120),
.B(n_4074),
.C(n_4130),
.Y(n_4162)
);

NAND4xp25_ASAP7_75t_L g4163 ( 
.A(n_4085),
.B(n_497),
.C(n_490),
.D(n_496),
.Y(n_4163)
);

NOR2xp33_ASAP7_75t_L g4164 ( 
.A(n_4091),
.B(n_496),
.Y(n_4164)
);

OAI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_4092),
.A2(n_502),
.B(n_499),
.Y(n_4165)
);

AOI211x1_ASAP7_75t_L g4166 ( 
.A1(n_4105),
.A2(n_503),
.B(n_498),
.C(n_499),
.Y(n_4166)
);

NOR2x1_ASAP7_75t_L g4167 ( 
.A(n_4090),
.B(n_503),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_4064),
.B(n_504),
.Y(n_4168)
);

NOR2x1_ASAP7_75t_L g4169 ( 
.A(n_4055),
.B(n_504),
.Y(n_4169)
);

AOI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_4082),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.Y(n_4170)
);

NOR5xp2_ASAP7_75t_L g4171 ( 
.A(n_4051),
.B(n_508),
.C(n_506),
.D(n_507),
.E(n_509),
.Y(n_4171)
);

AOI221xp5_ASAP7_75t_L g4172 ( 
.A1(n_4066),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.C(n_512),
.Y(n_4172)
);

NOR2xp33_ASAP7_75t_L g4173 ( 
.A(n_4078),
.B(n_514),
.Y(n_4173)
);

NOR2xp33_ASAP7_75t_L g4174 ( 
.A(n_4080),
.B(n_515),
.Y(n_4174)
);

NAND3xp33_ASAP7_75t_SL g4175 ( 
.A(n_4083),
.B(n_515),
.C(n_516),
.Y(n_4175)
);

AOI221xp5_ASAP7_75t_SL g4176 ( 
.A1(n_4063),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.C(n_519),
.Y(n_4176)
);

NAND2x1_ASAP7_75t_SL g4177 ( 
.A(n_4121),
.B(n_517),
.Y(n_4177)
);

NOR3xp33_ASAP7_75t_L g4178 ( 
.A(n_4096),
.B(n_520),
.C(n_519),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_SL g4179 ( 
.A(n_4060),
.B(n_518),
.Y(n_4179)
);

AOI211x1_ASAP7_75t_SL g4180 ( 
.A1(n_4068),
.A2(n_522),
.B(n_520),
.C(n_521),
.Y(n_4180)
);

OAI211xp5_ASAP7_75t_SL g4181 ( 
.A1(n_4086),
.A2(n_526),
.B(n_523),
.C(n_524),
.Y(n_4181)
);

NAND5xp2_ASAP7_75t_L g4182 ( 
.A(n_4101),
.B(n_526),
.C(n_523),
.D(n_524),
.E(n_527),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_SL g4183 ( 
.A(n_4067),
.B(n_527),
.Y(n_4183)
);

NOR2xp33_ASAP7_75t_L g4184 ( 
.A(n_4075),
.B(n_529),
.Y(n_4184)
);

NAND4xp25_ASAP7_75t_L g4185 ( 
.A(n_4109),
.B(n_531),
.C(n_529),
.D(n_530),
.Y(n_4185)
);

AOI211xp5_ASAP7_75t_SL g4186 ( 
.A1(n_4112),
.A2(n_534),
.B(n_530),
.C(n_533),
.Y(n_4186)
);

AOI221xp5_ASAP7_75t_L g4187 ( 
.A1(n_4066),
.A2(n_536),
.B1(n_533),
.B2(n_535),
.C(n_537),
.Y(n_4187)
);

NAND4xp25_ASAP7_75t_L g4188 ( 
.A(n_4087),
.B(n_539),
.C(n_537),
.D(n_538),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_L g4189 ( 
.A(n_4076),
.B(n_539),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_SL g4190 ( 
.A(n_4057),
.B(n_541),
.Y(n_4190)
);

AOI211xp5_ASAP7_75t_L g4191 ( 
.A1(n_4131),
.A2(n_544),
.B(n_542),
.C(n_543),
.Y(n_4191)
);

AOI321xp33_ASAP7_75t_L g4192 ( 
.A1(n_4072),
.A2(n_545),
.A3(n_547),
.B1(n_542),
.B2(n_543),
.C(n_546),
.Y(n_4192)
);

AOI211x1_ASAP7_75t_L g4193 ( 
.A1(n_4097),
.A2(n_548),
.B(n_546),
.C(n_547),
.Y(n_4193)
);

NOR3xp33_ASAP7_75t_L g4194 ( 
.A(n_4124),
.B(n_552),
.C(n_551),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_SL g4195 ( 
.A(n_4104),
.B(n_549),
.Y(n_4195)
);

NOR2x1p5_ASAP7_75t_L g4196 ( 
.A(n_4125),
.B(n_549),
.Y(n_4196)
);

NOR2x1_ASAP7_75t_L g4197 ( 
.A(n_4108),
.B(n_551),
.Y(n_4197)
);

OAI21xp5_ASAP7_75t_L g4198 ( 
.A1(n_4099),
.A2(n_555),
.B(n_554),
.Y(n_4198)
);

NAND3xp33_ASAP7_75t_SL g4199 ( 
.A(n_4088),
.B(n_4058),
.C(n_4065),
.Y(n_4199)
);

NAND3xp33_ASAP7_75t_SL g4200 ( 
.A(n_4054),
.B(n_4098),
.C(n_4107),
.Y(n_4200)
);

NOR4xp25_ASAP7_75t_L g4201 ( 
.A(n_4084),
.B(n_556),
.C(n_552),
.D(n_555),
.Y(n_4201)
);

CKINVDCx14_ASAP7_75t_R g4202 ( 
.A(n_4052),
.Y(n_4202)
);

NOR3xp33_ASAP7_75t_L g4203 ( 
.A(n_4089),
.B(n_558),
.C(n_557),
.Y(n_4203)
);

AND2x2_ASAP7_75t_L g4204 ( 
.A(n_4118),
.B(n_556),
.Y(n_4204)
);

NOR4xp25_ASAP7_75t_L g4205 ( 
.A(n_4089),
.B(n_560),
.C(n_558),
.D(n_559),
.Y(n_4205)
);

NOR3xp33_ASAP7_75t_L g4206 ( 
.A(n_4089),
.B(n_562),
.C(n_561),
.Y(n_4206)
);

NAND5xp2_ASAP7_75t_L g4207 ( 
.A(n_4118),
.B(n_562),
.C(n_560),
.D(n_561),
.E(n_563),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4064),
.B(n_563),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4064),
.B(n_564),
.Y(n_4209)
);

NOR5xp2_ASAP7_75t_L g4210 ( 
.A(n_4089),
.B(n_567),
.C(n_564),
.D(n_565),
.E(n_568),
.Y(n_4210)
);

A2O1A1Ixp33_ASAP7_75t_L g4211 ( 
.A1(n_4085),
.A2(n_571),
.B(n_569),
.C(n_570),
.Y(n_4211)
);

NAND4xp25_ASAP7_75t_L g4212 ( 
.A(n_4089),
.B(n_572),
.C(n_569),
.D(n_570),
.Y(n_4212)
);

OAI21xp33_ASAP7_75t_L g4213 ( 
.A1(n_4118),
.A2(n_573),
.B(n_574),
.Y(n_4213)
);

AOI22xp33_ASAP7_75t_L g4214 ( 
.A1(n_4082),
.A2(n_575),
.B1(n_573),
.B2(n_574),
.Y(n_4214)
);

OAI211xp5_ASAP7_75t_L g4215 ( 
.A1(n_4115),
.A2(n_578),
.B(n_576),
.C(n_577),
.Y(n_4215)
);

AND2x4_ASAP7_75t_L g4216 ( 
.A(n_4056),
.B(n_577),
.Y(n_4216)
);

OAI221xp5_ASAP7_75t_L g4217 ( 
.A1(n_4056),
.A2(n_580),
.B1(n_576),
.B2(n_579),
.C(n_581),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_4204),
.B(n_579),
.Y(n_4218)
);

NAND3xp33_ASAP7_75t_L g4219 ( 
.A(n_4186),
.B(n_581),
.C(n_582),
.Y(n_4219)
);

NOR2x1_ASAP7_75t_L g4220 ( 
.A(n_4138),
.B(n_4136),
.Y(n_4220)
);

OAI322xp33_ASAP7_75t_L g4221 ( 
.A1(n_4202),
.A2(n_4145),
.A3(n_4190),
.B1(n_4134),
.B2(n_4179),
.C1(n_4149),
.C2(n_4133),
.Y(n_4221)
);

NOR4xp25_ASAP7_75t_L g4222 ( 
.A(n_4215),
.B(n_584),
.C(n_582),
.D(n_583),
.Y(n_4222)
);

NOR3x1_ASAP7_75t_L g4223 ( 
.A(n_4152),
.B(n_584),
.C(n_585),
.Y(n_4223)
);

NAND3xp33_ASAP7_75t_L g4224 ( 
.A(n_4172),
.B(n_585),
.C(n_586),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4177),
.Y(n_4225)
);

INVxp33_ASAP7_75t_L g4226 ( 
.A(n_4169),
.Y(n_4226)
);

NOR2x1_ASAP7_75t_L g4227 ( 
.A(n_4163),
.B(n_588),
.Y(n_4227)
);

HB1xp67_ASAP7_75t_L g4228 ( 
.A(n_4216),
.Y(n_4228)
);

NAND3xp33_ASAP7_75t_SL g4229 ( 
.A(n_4187),
.B(n_588),
.C(n_589),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4216),
.Y(n_4230)
);

INVx1_ASAP7_75t_SL g4231 ( 
.A(n_4141),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4201),
.B(n_589),
.Y(n_4232)
);

AOI322xp5_ASAP7_75t_L g4233 ( 
.A1(n_4162),
.A2(n_595),
.A3(n_594),
.B1(n_592),
.B2(n_590),
.C1(n_591),
.C2(n_593),
.Y(n_4233)
);

AOI22xp33_ASAP7_75t_L g4234 ( 
.A1(n_4142),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.Y(n_4234)
);

NAND2x1p5_ASAP7_75t_L g4235 ( 
.A(n_4197),
.B(n_4167),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_SL g4236 ( 
.A(n_4205),
.B(n_595),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_SL g4237 ( 
.A(n_4150),
.B(n_596),
.Y(n_4237)
);

AND2x4_ASAP7_75t_L g4238 ( 
.A(n_4165),
.B(n_596),
.Y(n_4238)
);

NAND4xp75_ASAP7_75t_L g4239 ( 
.A(n_4144),
.B(n_599),
.C(n_597),
.D(n_598),
.Y(n_4239)
);

INVx1_ASAP7_75t_SL g4240 ( 
.A(n_4168),
.Y(n_4240)
);

NAND3xp33_ASAP7_75t_SL g4241 ( 
.A(n_4171),
.B(n_598),
.C(n_599),
.Y(n_4241)
);

NAND3xp33_ASAP7_75t_SL g4242 ( 
.A(n_4139),
.B(n_601),
.C(n_602),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4208),
.Y(n_4243)
);

AOI22xp33_ASAP7_75t_L g4244 ( 
.A1(n_4157),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_4244)
);

AND2x4_ASAP7_75t_L g4245 ( 
.A(n_4196),
.B(n_603),
.Y(n_4245)
);

NOR2x1_ASAP7_75t_L g4246 ( 
.A(n_4212),
.B(n_605),
.Y(n_4246)
);

OR2x2_ASAP7_75t_L g4247 ( 
.A(n_4182),
.B(n_606),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4209),
.Y(n_4248)
);

NOR2xp67_ASAP7_75t_L g4249 ( 
.A(n_4175),
.B(n_606),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4146),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4166),
.Y(n_4251)
);

NOR2x1_ASAP7_75t_L g4252 ( 
.A(n_4207),
.B(n_4188),
.Y(n_4252)
);

INVxp67_ASAP7_75t_L g4253 ( 
.A(n_4159),
.Y(n_4253)
);

NOR3xp33_ASAP7_75t_L g4254 ( 
.A(n_4147),
.B(n_607),
.C(n_608),
.Y(n_4254)
);

INVx2_ASAP7_75t_SL g4255 ( 
.A(n_4183),
.Y(n_4255)
);

AOI221xp5_ASAP7_75t_SL g4256 ( 
.A1(n_4198),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.C(n_611),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4193),
.B(n_609),
.Y(n_4257)
);

NAND4xp75_ASAP7_75t_L g4258 ( 
.A(n_4176),
.B(n_612),
.C(n_610),
.D(n_611),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4192),
.Y(n_4259)
);

NAND3xp33_ASAP7_75t_L g4260 ( 
.A(n_4153),
.B(n_4191),
.C(n_4154),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4213),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4151),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4164),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_4158),
.B(n_612),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4184),
.Y(n_4265)
);

NOR3xp33_ASAP7_75t_L g4266 ( 
.A(n_4199),
.B(n_613),
.C(n_614),
.Y(n_4266)
);

NOR2x1_ASAP7_75t_L g4267 ( 
.A(n_4160),
.B(n_613),
.Y(n_4267)
);

AND2x4_ASAP7_75t_L g4268 ( 
.A(n_4178),
.B(n_615),
.Y(n_4268)
);

NOR2xp67_ASAP7_75t_L g4269 ( 
.A(n_4156),
.B(n_616),
.Y(n_4269)
);

NAND3xp33_ASAP7_75t_SL g4270 ( 
.A(n_4180),
.B(n_4210),
.C(n_4135),
.Y(n_4270)
);

NOR3xp33_ASAP7_75t_L g4271 ( 
.A(n_4195),
.B(n_617),
.C(n_618),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4189),
.B(n_620),
.Y(n_4272)
);

NOR2x1_ASAP7_75t_L g4273 ( 
.A(n_4155),
.B(n_621),
.Y(n_4273)
);

AND2x4_ASAP7_75t_L g4274 ( 
.A(n_4194),
.B(n_621),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4173),
.Y(n_4275)
);

NAND4xp25_ASAP7_75t_L g4276 ( 
.A(n_4200),
.B(n_624),
.C(n_622),
.D(n_623),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_4203),
.B(n_622),
.Y(n_4277)
);

NOR2xp67_ASAP7_75t_SL g4278 ( 
.A(n_4217),
.B(n_4148),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4170),
.Y(n_4279)
);

AOI22xp33_ASAP7_75t_L g4280 ( 
.A1(n_4181),
.A2(n_626),
.B1(n_623),
.B2(n_625),
.Y(n_4280)
);

AOI21xp5_ASAP7_75t_L g4281 ( 
.A1(n_4211),
.A2(n_4161),
.B(n_4140),
.Y(n_4281)
);

NOR2x1_ASAP7_75t_L g4282 ( 
.A(n_4185),
.B(n_626),
.Y(n_4282)
);

NOR2xp33_ASAP7_75t_L g4283 ( 
.A(n_4174),
.B(n_627),
.Y(n_4283)
);

OR2x2_ASAP7_75t_L g4284 ( 
.A(n_4206),
.B(n_628),
.Y(n_4284)
);

AND2x4_ASAP7_75t_L g4285 ( 
.A(n_4214),
.B(n_628),
.Y(n_4285)
);

NAND5xp2_ASAP7_75t_L g4286 ( 
.A(n_4137),
.B(n_631),
.C(n_629),
.D(n_630),
.E(n_632),
.Y(n_4286)
);

NOR2x1_ASAP7_75t_L g4287 ( 
.A(n_4143),
.B(n_630),
.Y(n_4287)
);

NAND4xp25_ASAP7_75t_L g4288 ( 
.A(n_4144),
.B(n_634),
.C(n_632),
.D(n_633),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4177),
.Y(n_4289)
);

INVxp67_ASAP7_75t_SL g4290 ( 
.A(n_4210),
.Y(n_4290)
);

NOR2x1_ASAP7_75t_L g4291 ( 
.A(n_4138),
.B(n_635),
.Y(n_4291)
);

NOR2xp33_ASAP7_75t_L g4292 ( 
.A(n_4152),
.B(n_635),
.Y(n_4292)
);

AOI22xp5_ASAP7_75t_L g4293 ( 
.A1(n_4202),
.A2(n_638),
.B1(n_636),
.B2(n_637),
.Y(n_4293)
);

CKINVDCx20_ASAP7_75t_R g4294 ( 
.A(n_4253),
.Y(n_4294)
);

OR3x2_ASAP7_75t_L g4295 ( 
.A(n_4288),
.B(n_636),
.C(n_637),
.Y(n_4295)
);

INVxp67_ASAP7_75t_SL g4296 ( 
.A(n_4228),
.Y(n_4296)
);

XNOR2xp5_ASAP7_75t_L g4297 ( 
.A(n_4252),
.B(n_639),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4291),
.Y(n_4298)
);

NOR2x1_ASAP7_75t_L g4299 ( 
.A(n_4220),
.B(n_639),
.Y(n_4299)
);

OR2x2_ASAP7_75t_L g4300 ( 
.A(n_4241),
.B(n_640),
.Y(n_4300)
);

NOR3xp33_ASAP7_75t_L g4301 ( 
.A(n_4221),
.B(n_651),
.C(n_641),
.Y(n_4301)
);

NOR3xp33_ASAP7_75t_SL g4302 ( 
.A(n_4229),
.B(n_642),
.C(n_643),
.Y(n_4302)
);

INVxp33_ASAP7_75t_L g4303 ( 
.A(n_4267),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4218),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_4231),
.B(n_642),
.Y(n_4305)
);

NAND4xp25_ASAP7_75t_L g4306 ( 
.A(n_4223),
.B(n_646),
.C(n_643),
.D(n_645),
.Y(n_4306)
);

AND2x2_ASAP7_75t_SL g4307 ( 
.A(n_4222),
.B(n_645),
.Y(n_4307)
);

NOR3xp33_ASAP7_75t_L g4308 ( 
.A(n_4250),
.B(n_648),
.C(n_649),
.Y(n_4308)
);

NOR3xp33_ASAP7_75t_L g4309 ( 
.A(n_4232),
.B(n_4292),
.C(n_4283),
.Y(n_4309)
);

OAI211xp5_ASAP7_75t_L g4310 ( 
.A1(n_4290),
.A2(n_651),
.B(n_648),
.C(n_650),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4230),
.Y(n_4311)
);

AND4x1_ASAP7_75t_L g4312 ( 
.A(n_4266),
.B(n_653),
.C(n_650),
.D(n_652),
.Y(n_4312)
);

XNOR2x1_ASAP7_75t_L g4313 ( 
.A(n_4239),
.B(n_654),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4235),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4247),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4257),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4251),
.B(n_4245),
.Y(n_4317)
);

NAND3x1_ASAP7_75t_SL g4318 ( 
.A(n_4227),
.B(n_654),
.C(n_655),
.Y(n_4318)
);

INVx1_ASAP7_75t_SL g4319 ( 
.A(n_4245),
.Y(n_4319)
);

INVx2_ASAP7_75t_SL g4320 ( 
.A(n_4225),
.Y(n_4320)
);

HB1xp67_ASAP7_75t_L g4321 ( 
.A(n_4249),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4264),
.Y(n_4322)
);

NAND3xp33_ASAP7_75t_SL g4323 ( 
.A(n_4226),
.B(n_655),
.C(n_656),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4233),
.B(n_657),
.Y(n_4324)
);

NOR2x1_ASAP7_75t_L g4325 ( 
.A(n_4289),
.B(n_657),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_4282),
.B(n_658),
.Y(n_4326)
);

OR2x6_ASAP7_75t_L g4327 ( 
.A(n_4255),
.B(n_659),
.Y(n_4327)
);

XNOR2x1_ASAP7_75t_L g4328 ( 
.A(n_4258),
.B(n_660),
.Y(n_4328)
);

NOR3x1_ASAP7_75t_L g4329 ( 
.A(n_4219),
.B(n_660),
.C(n_661),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4293),
.B(n_661),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4238),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4238),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4284),
.Y(n_4333)
);

INVx2_ASAP7_75t_L g4334 ( 
.A(n_4272),
.Y(n_4334)
);

NOR2xp33_ASAP7_75t_L g4335 ( 
.A(n_4276),
.B(n_662),
.Y(n_4335)
);

NAND4xp75_ASAP7_75t_L g4336 ( 
.A(n_4287),
.B(n_665),
.C(n_663),
.D(n_664),
.Y(n_4336)
);

NAND2x1p5_ASAP7_75t_SL g4337 ( 
.A(n_4279),
.B(n_4246),
.Y(n_4337)
);

AND2x4_ASAP7_75t_L g4338 ( 
.A(n_4261),
.B(n_663),
.Y(n_4338)
);

HB1xp67_ASAP7_75t_L g4339 ( 
.A(n_4269),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_SL g4340 ( 
.A(n_4256),
.B(n_4274),
.Y(n_4340)
);

INVxp67_ASAP7_75t_L g4341 ( 
.A(n_4286),
.Y(n_4341)
);

OAI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_4281),
.A2(n_664),
.B(n_665),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_4274),
.Y(n_4343)
);

AND2x4_ASAP7_75t_L g4344 ( 
.A(n_4243),
.B(n_666),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4259),
.B(n_666),
.Y(n_4345)
);

NOR4xp25_ASAP7_75t_L g4346 ( 
.A(n_4237),
.B(n_4236),
.C(n_4270),
.D(n_4240),
.Y(n_4346)
);

NAND4xp25_ASAP7_75t_L g4347 ( 
.A(n_4260),
.B(n_669),
.C(n_667),
.D(n_668),
.Y(n_4347)
);

NAND4xp75_ASAP7_75t_L g4348 ( 
.A(n_4273),
.B(n_4277),
.C(n_4275),
.D(n_4265),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4327),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4327),
.Y(n_4350)
);

CKINVDCx20_ASAP7_75t_R g4351 ( 
.A(n_4294),
.Y(n_4351)
);

INVx1_ASAP7_75t_SL g4352 ( 
.A(n_4307),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_4296),
.B(n_4280),
.Y(n_4353)
);

HB1xp67_ASAP7_75t_L g4354 ( 
.A(n_4299),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_4338),
.B(n_4254),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4300),
.Y(n_4356)
);

OA22x2_ASAP7_75t_L g4357 ( 
.A1(n_4342),
.A2(n_4285),
.B1(n_4268),
.B2(n_4248),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4325),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_4319),
.B(n_4244),
.Y(n_4359)
);

AOI22xp5_ASAP7_75t_L g4360 ( 
.A1(n_4311),
.A2(n_4242),
.B1(n_4271),
.B2(n_4278),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_4345),
.B(n_4234),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_SL g4362 ( 
.A(n_4298),
.B(n_4224),
.Y(n_4362)
);

AND3x1_ASAP7_75t_L g4363 ( 
.A(n_4346),
.B(n_4262),
.C(n_4263),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_4344),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4297),
.Y(n_4365)
);

AOI22xp5_ASAP7_75t_SL g4366 ( 
.A1(n_4303),
.A2(n_670),
.B1(n_667),
.B2(n_669),
.Y(n_4366)
);

HB1xp67_ASAP7_75t_L g4367 ( 
.A(n_4313),
.Y(n_4367)
);

OAI21xp5_ASAP7_75t_SL g4368 ( 
.A1(n_4328),
.A2(n_670),
.B(n_671),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4295),
.Y(n_4369)
);

AND3x4_ASAP7_75t_L g4370 ( 
.A(n_4302),
.B(n_671),
.C(n_672),
.Y(n_4370)
);

OAI211xp5_ASAP7_75t_SL g4371 ( 
.A1(n_4341),
.A2(n_676),
.B(n_672),
.C(n_674),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4305),
.Y(n_4372)
);

NOR2xp33_ASAP7_75t_L g4373 ( 
.A(n_4306),
.B(n_674),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4317),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4318),
.Y(n_4375)
);

AOI22xp33_ASAP7_75t_L g4376 ( 
.A1(n_4301),
.A2(n_4320),
.B1(n_4314),
.B2(n_4339),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4326),
.Y(n_4377)
);

INVx1_ASAP7_75t_SL g4378 ( 
.A(n_4336),
.Y(n_4378)
);

BUFx2_ASAP7_75t_L g4379 ( 
.A(n_4321),
.Y(n_4379)
);

INVxp33_ASAP7_75t_SL g4380 ( 
.A(n_4329),
.Y(n_4380)
);

BUFx2_ASAP7_75t_L g4381 ( 
.A(n_4337),
.Y(n_4381)
);

AOI221xp5_ASAP7_75t_SL g4382 ( 
.A1(n_4340),
.A2(n_679),
.B1(n_677),
.B2(n_678),
.C(n_680),
.Y(n_4382)
);

AO22x2_ASAP7_75t_L g4383 ( 
.A1(n_4370),
.A2(n_4348),
.B1(n_4310),
.B2(n_4323),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4354),
.Y(n_4384)
);

AO22x2_ASAP7_75t_L g4385 ( 
.A1(n_4352),
.A2(n_4304),
.B1(n_4332),
.B2(n_4331),
.Y(n_4385)
);

OAI22x1_ASAP7_75t_L g4386 ( 
.A1(n_4360),
.A2(n_4312),
.B1(n_4334),
.B2(n_4343),
.Y(n_4386)
);

NOR2x1_ASAP7_75t_L g4387 ( 
.A(n_4358),
.B(n_4347),
.Y(n_4387)
);

AO22x2_ASAP7_75t_L g4388 ( 
.A1(n_4375),
.A2(n_4315),
.B1(n_4322),
.B2(n_4316),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4351),
.Y(n_4389)
);

INVx1_ASAP7_75t_SL g4390 ( 
.A(n_4366),
.Y(n_4390)
);

AO22x2_ASAP7_75t_L g4391 ( 
.A1(n_4378),
.A2(n_4368),
.B1(n_4349),
.B2(n_4350),
.Y(n_4391)
);

OAI22xp5_ASAP7_75t_L g4392 ( 
.A1(n_4376),
.A2(n_4324),
.B1(n_4330),
.B2(n_4335),
.Y(n_4392)
);

AOI22xp33_ASAP7_75t_L g4393 ( 
.A1(n_4381),
.A2(n_4309),
.B1(n_4333),
.B2(n_4308),
.Y(n_4393)
);

OAI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_4374),
.A2(n_679),
.B1(n_677),
.B2(n_678),
.Y(n_4394)
);

OAI22x1_ASAP7_75t_L g4395 ( 
.A1(n_4379),
.A2(n_682),
.B1(n_680),
.B2(n_681),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4353),
.Y(n_4396)
);

OAI22x1_ASAP7_75t_L g4397 ( 
.A1(n_4369),
.A2(n_683),
.B1(n_681),
.B2(n_682),
.Y(n_4397)
);

OAI22xp5_ASAP7_75t_L g4398 ( 
.A1(n_4363),
.A2(n_685),
.B1(n_683),
.B2(n_684),
.Y(n_4398)
);

BUFx2_ASAP7_75t_L g4399 ( 
.A(n_4364),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4385),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4389),
.B(n_4356),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4398),
.Y(n_4402)
);

INVxp33_ASAP7_75t_SL g4403 ( 
.A(n_4386),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4399),
.Y(n_4404)
);

OAI22x1_ASAP7_75t_L g4405 ( 
.A1(n_4390),
.A2(n_4373),
.B1(n_4377),
.B2(n_4365),
.Y(n_4405)
);

OAI22x1_ASAP7_75t_L g4406 ( 
.A1(n_4384),
.A2(n_4367),
.B1(n_4362),
.B2(n_4372),
.Y(n_4406)
);

AOI22xp5_ASAP7_75t_L g4407 ( 
.A1(n_4383),
.A2(n_4380),
.B1(n_4371),
.B2(n_4357),
.Y(n_4407)
);

OAI21x1_ASAP7_75t_L g4408 ( 
.A1(n_4387),
.A2(n_4355),
.B(n_4359),
.Y(n_4408)
);

XNOR2xp5_ASAP7_75t_L g4409 ( 
.A(n_4391),
.B(n_4361),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4388),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4400),
.Y(n_4411)
);

AOI22xp5_ASAP7_75t_L g4412 ( 
.A1(n_4403),
.A2(n_4396),
.B1(n_4382),
.B2(n_4392),
.Y(n_4412)
);

OA21x2_ASAP7_75t_L g4413 ( 
.A1(n_4410),
.A2(n_4393),
.B(n_4394),
.Y(n_4413)
);

NOR3x2_ASAP7_75t_L g4414 ( 
.A(n_4409),
.B(n_4406),
.C(n_4405),
.Y(n_4414)
);

OAI21xp5_ASAP7_75t_L g4415 ( 
.A1(n_4404),
.A2(n_4395),
.B(n_4397),
.Y(n_4415)
);

INVxp67_ASAP7_75t_L g4416 ( 
.A(n_4401),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4402),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4414),
.Y(n_4418)
);

AOI22xp33_ASAP7_75t_L g4419 ( 
.A1(n_4411),
.A2(n_4408),
.B1(n_4407),
.B2(n_686),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4416),
.Y(n_4420)
);

AOI221xp5_ASAP7_75t_R g4421 ( 
.A1(n_4412),
.A2(n_686),
.B1(n_684),
.B2(n_685),
.C(n_688),
.Y(n_4421)
);

INVx1_ASAP7_75t_SL g4422 ( 
.A(n_4413),
.Y(n_4422)
);

AOI222xp33_ASAP7_75t_L g4423 ( 
.A1(n_4422),
.A2(n_4417),
.B1(n_4415),
.B2(n_692),
.C1(n_694),
.C2(n_689),
.Y(n_4423)
);

AOI21xp33_ASAP7_75t_L g4424 ( 
.A1(n_4418),
.A2(n_689),
.B(n_690),
.Y(n_4424)
);

AOI22xp5_ASAP7_75t_L g4425 ( 
.A1(n_4423),
.A2(n_4420),
.B1(n_4419),
.B2(n_4421),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_4425),
.B(n_4424),
.Y(n_4426)
);

OR2x6_ASAP7_75t_L g4427 ( 
.A(n_4426),
.B(n_693),
.Y(n_4427)
);

OAI22xp33_ASAP7_75t_L g4428 ( 
.A1(n_4427),
.A2(n_698),
.B1(n_694),
.B2(n_695),
.Y(n_4428)
);

AOI211xp5_ASAP7_75t_L g4429 ( 
.A1(n_4428),
.A2(n_704),
.B(n_702),
.C(n_703),
.Y(n_4429)
);


endmodule