module fake_jpeg_29864_n_71 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_67;
wire n_66;

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_35),
.B(n_37),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_38),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

A2O1A1O1Ixp25_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_25),
.B(n_26),
.C(n_20),
.D(n_13),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_24),
.B(n_22),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_46),
.B(n_3),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_26),
.C(n_19),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_30),
.C(n_2),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_30),
.B1(n_31),
.B2(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_53),
.C(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_54),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_52),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_2),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_11),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_59),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.C(n_52),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_4),
.C(n_5),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_41),
.B1(n_17),
.B2(n_16),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_61),
.B(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_57),
.Y(n_69)
);

A2O1A1O1Ixp25_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_67),
.B(n_15),
.C(n_12),
.D(n_7),
.Y(n_70)
);

AOI321xp33_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_71)
);


endmodule