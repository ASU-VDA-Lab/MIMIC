module fake_jpeg_11698_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_32),
.B(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_4),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_72),
.Y(n_74)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_46),
.B1(n_61),
.B2(n_50),
.Y(n_79)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_3),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_81),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_80),
.B(n_63),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_48),
.B1(n_50),
.B2(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_52),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_43),
.Y(n_88)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_98),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_13),
.C(n_14),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_80),
.B1(n_73),
.B2(n_48),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_93),
.B1(n_15),
.B2(n_40),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_51),
.B1(n_55),
.B2(n_60),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_51),
.B1(n_55),
.B2(n_49),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_53),
.B(n_58),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_95),
.C(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_101),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_58),
.B(n_56),
.C(n_24),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_58),
.B1(n_56),
.B2(n_23),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_106),
.C(n_21),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_82),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_56),
.B1(n_6),
.B2(n_7),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_27),
.C(n_38),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_109),
.C(n_112),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_106),
.B(n_10),
.C(n_11),
.Y(n_109)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_10),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_118),
.B(n_119),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_28),
.C(n_37),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_26),
.C(n_35),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_89),
.B(n_15),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_123),
.B(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_16),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_110),
.B1(n_117),
.B2(n_121),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_136),
.B1(n_130),
.B2(n_128),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_30),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_133),
.Y(n_140)
);

INVxp33_ASAP7_75t_SL g134 ( 
.A(n_107),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_34),
.B(n_119),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_111),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_138),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_125),
.B1(n_135),
.B2(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_139),
.B(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_137),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_131),
.C(n_138),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_145),
.B(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_142),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_142),
.Y(n_151)
);


endmodule