module real_jpeg_23782_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_1),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_2),
.A2(n_33),
.B1(n_65),
.B2(n_66),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_2),
.A2(n_33),
.B1(n_59),
.B2(n_60),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g58 ( 
.A(n_4),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_5),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_121),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_121),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_121),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_81),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_81),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_81),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_7),
.A2(n_66),
.B1(n_161),
.B2(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_161),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_161),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_8),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_8),
.B(n_74),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_8),
.B(n_28),
.C(n_40),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_165),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_8),
.B(n_87),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_8),
.A2(n_25),
.B1(n_238),
.B2(n_241),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_10),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_169),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_169),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_169),
.Y(n_238)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_13),
.A2(n_49),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_13),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_14),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_151)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_15),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_142),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_20),
.B(n_123),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_97),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_21),
.A2(n_76),
.B1(n_77),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_21),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_50),
.B2(n_75),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_22),
.A2(n_51),
.B(n_53),
.Y(n_140)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_24),
.A2(n_34),
.B1(n_51),
.B2(n_302),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_32),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_25),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_25),
.A2(n_102),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_25),
.A2(n_154),
.B1(n_231),
.B2(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_25),
.A2(n_32),
.B(n_152),
.Y(n_256)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_26),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_26),
.A2(n_151),
.B1(n_153),
.B2(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_26),
.A2(n_103),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_27),
.B(n_243),
.Y(n_242)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_29),
.Y(n_241)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_30),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_30),
.B(n_165),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_32),
.Y(n_105)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_34),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_43),
.B(n_46),
.Y(n_34)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_35),
.A2(n_42),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_35),
.A2(n_42),
.B1(n_217),
.B2(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_35),
.A2(n_90),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_37),
.A2(n_38),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_37),
.A2(n_85),
.B(n_252),
.C(n_254),
.Y(n_251)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_38),
.B(n_213),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_L g254 ( 
.A(n_38),
.B(n_59),
.C(n_84),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_42),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_42),
.A2(n_93),
.B(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_42),
.B(n_165),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_44),
.A2(n_92),
.B1(n_94),
.B2(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_47),
.A2(n_91),
.B(n_94),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_68),
.B(n_70),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_119),
.B(n_122),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_54),
.A2(n_56),
.B1(n_168),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_71),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_55),
.A2(n_74),
.B1(n_164),
.B2(n_167),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_55),
.A2(n_74),
.B1(n_120),
.B2(n_175),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_56),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_57),
.A2(n_60),
.B(n_166),
.C(n_188),
.Y(n_187)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_60),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_59),
.B(n_62),
.C(n_65),
.Y(n_188)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g253 ( 
.A(n_60),
.B(n_165),
.CON(n_253),
.SN(n_253)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_65),
.B(n_165),
.Y(n_166)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_67),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_69),
.B(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_89),
.B(n_96),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_86),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_88),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_82),
.A2(n_87),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_82),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_82),
.A2(n_87),
.B1(n_203),
.B2(n_253),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_82),
.A2(n_137),
.B(n_181),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_116),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_86),
.A2(n_179),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_87),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_91),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_92),
.A2(n_94),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_92),
.A2(n_94),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_125),
.B1(n_138),
.B2(n_139),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_96),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_97),
.A2(n_98),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.C(n_117),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_99),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_108),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_100),
.A2(n_101),
.B1(n_108),
.B2(n_109),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_106),
.A2(n_186),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_107),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_304)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_140),
.Y(n_123)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_309),
.B(n_315),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_297),
.B(n_308),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_205),
.B(n_285),
.C(n_296),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_190),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_146),
.B(n_190),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_170),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_157),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_148),
.B(n_157),
.C(n_170),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_149),
.B(n_156),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.C(n_163),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_192),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_182),
.B2(n_189),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_173),
.B(n_177),
.C(n_189),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B(n_180),
.Y(n_177)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_195),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_191),
.B(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_193),
.B(n_195),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_196),
.A2(n_199),
.B1(n_200),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_201),
.B(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_284),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_279),
.B(n_283),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_264),
.B(n_278),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_247),
.B(n_263),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_227),
.B(n_246),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_214),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_222),
.C(n_225),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_220),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_226),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_234),
.B(n_245),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_239),
.B(n_244),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_262),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_262),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_257),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_258),
.C(n_259),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_255),
.B2(n_256),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_266),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_271),
.B2(n_272),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_274),
.C(n_276),
.Y(n_282)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_273),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_290),
.C(n_295),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_293),
.C(n_294),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_307),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_303),
.B1(n_305),
.B2(n_306),
.Y(n_300)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_306),
.C(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);


endmodule