module fake_jpeg_10153_n_78 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_38),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.C(n_1),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_2),
.C(n_3),
.Y(n_58)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_9),
.B1(n_20),
.B2(n_19),
.Y(n_49)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_2),
.Y(n_55)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_13),
.B1(n_24),
.B2(n_22),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_10),
.B(n_21),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_28),
.B(n_33),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_46),
.B(n_49),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_57),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.C(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_3),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_4),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_4),
.C(n_5),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_6),
.Y(n_70)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_68),
.C(n_47),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_62),
.B(n_61),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_65),
.B(n_59),
.C(n_53),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_45),
.B1(n_66),
.B2(n_11),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_7),
.Y(n_78)
);


endmodule