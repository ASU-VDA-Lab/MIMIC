module fake_jpeg_27276_n_31 (n_3, n_2, n_1, n_0, n_4, n_5, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_5),
.Y(n_6)
);

BUFx4f_ASAP7_75t_SL g7 ( 
.A(n_2),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_0),
.Y(n_12)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_15),
.B(n_7),
.C(n_8),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_14),
.B1(n_7),
.B2(n_10),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_6),
.B(n_3),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_15),
.A2(n_7),
.B(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_17),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_3),
.C(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_21),
.B(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_11),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_11),
.C(n_10),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI211xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_25),
.B(n_28),
.C(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_11),
.Y(n_31)
);


endmodule