module fake_jpeg_7282_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_23),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_18),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_50),
.B(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_25),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_32),
.B1(n_28),
.B2(n_25),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_38),
.Y(n_69)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_35),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_75),
.B1(n_81),
.B2(n_60),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_88),
.Y(n_112)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_18),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_29),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_98),
.B1(n_38),
.B2(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_67),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_36),
.B1(n_39),
.B2(n_26),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_114),
.B1(n_125),
.B2(n_38),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_39),
.C(n_42),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_115),
.C(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_105),
.B(n_110),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_123),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_39),
.Y(n_109)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_111),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_26),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_36),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_118),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_41),
.B1(n_38),
.B2(n_55),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_97),
.B1(n_75),
.B2(n_46),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_54),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_76),
.A2(n_41),
.B1(n_67),
.B2(n_38),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_135),
.B1(n_139),
.B2(n_84),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_76),
.B1(n_120),
.B2(n_113),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_132),
.B1(n_149),
.B2(n_57),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_91),
.B1(n_79),
.B2(n_96),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_150),
.B1(n_151),
.B2(n_124),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_102),
.B1(n_101),
.B2(n_100),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_104),
.C(n_99),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_137),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_87),
.B1(n_84),
.B2(n_95),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_136),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_35),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_144),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_141),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_49),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_33),
.B1(n_25),
.B2(n_34),
.Y(n_181)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_147),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_57),
.B1(n_46),
.B2(n_85),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_46),
.B1(n_57),
.B2(n_85),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_109),
.B1(n_110),
.B2(n_99),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_35),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_88),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_78),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_42),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_166),
.B1(n_170),
.B2(n_181),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_171),
.C(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_169),
.B1(n_185),
.B2(n_144),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_116),
.B(n_111),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_168),
.B(n_178),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_111),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_119),
.B1(n_125),
.B2(n_111),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_116),
.B1(n_33),
.B2(n_25),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_49),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_40),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_175),
.B(n_180),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_34),
.B(n_20),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_0),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_0),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_86),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_34),
.B(n_20),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_43),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_42),
.C(n_40),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_184),
.C(n_189),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_40),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_130),
.A2(n_58),
.B1(n_78),
.B2(n_33),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_31),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_134),
.A2(n_95),
.B(n_30),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_129),
.B(n_42),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_40),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_43),
.C(n_19),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_127),
.A2(n_58),
.B1(n_33),
.B2(n_30),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_31),
.B1(n_19),
.B2(n_17),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_148),
.B1(n_127),
.B2(n_140),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_191),
.B(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_198),
.Y(n_223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_127),
.B(n_155),
.C(n_148),
.D(n_147),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_190),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_204),
.B1(n_208),
.B2(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_201),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_159),
.B(n_172),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_215),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_128),
.B1(n_136),
.B2(n_141),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_164),
.B1(n_186),
.B2(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_141),
.B1(n_19),
.B2(n_17),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_17),
.Y(n_209)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_216),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_1),
.C(n_2),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_17),
.B1(n_19),
.B2(n_43),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_9),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_218),
.A2(n_176),
.B1(n_11),
.B2(n_12),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_173),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_222),
.A2(n_205),
.B(n_214),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_171),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_227),
.B(n_233),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_202),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_162),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_241),
.C(n_246),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_186),
.B1(n_176),
.B2(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_236),
.A2(n_242),
.B1(n_192),
.B2(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_212),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_168),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_211),
.A2(n_168),
.B1(n_86),
.B2(n_72),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_209),
.C(n_219),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_224),
.C(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_257),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_216),
.B(n_210),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_SL g280 ( 
.A1(n_256),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_229),
.B(n_218),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_200),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_264),
.B1(n_232),
.B2(n_240),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_222),
.A2(n_9),
.B(n_14),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_6),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_242),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_271),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_241),
.A3(n_233),
.B1(n_225),
.B2(n_244),
.C1(n_238),
.C2(n_245),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_256),
.B(n_265),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_246),
.C(n_10),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_8),
.C(n_14),
.Y(n_279)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_7),
.C(n_13),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.C(n_284),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_7),
.C(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_1),
.C(n_3),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_273),
.B(n_249),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_270),
.C(n_274),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_295),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_252),
.Y(n_294)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_276),
.B(n_263),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_266),
.C(n_254),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_261),
.C(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_264),
.Y(n_300)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_303),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_261),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_287),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_262),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_296),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_6),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_280),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_310),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_280),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_317),
.C(n_306),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_285),
.B(n_287),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_299),
.B(n_304),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_280),
.B1(n_288),
.B2(n_3),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

INVx11_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_6),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_12),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_320),
.B(n_324),
.CI(n_314),
.CON(n_327),
.SN(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_321),
.A2(n_323),
.B(n_315),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_302),
.B(n_11),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_15),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_316),
.B(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_327),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_328),
.B1(n_322),
.B2(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_312),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_15),
.Y(n_332)
);

OAI321xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_4),
.A3(n_15),
.B1(n_323),
.B2(n_326),
.C(n_256),
.Y(n_333)
);


endmodule