module real_jpeg_18028_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_286;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_398),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_1),
.B(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_2),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_3),
.Y(n_182)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_3),
.Y(n_322)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_4),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_4),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_4),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_5),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_5),
.B(n_49),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_5),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_5),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_5),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_6),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_6),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_6),
.B(n_178),
.Y(n_177)
);

AND2x4_ASAP7_75t_SL g181 ( 
.A(n_6),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_6),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_6),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g255 ( 
.A(n_6),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_6),
.B(n_288),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_8),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_9),
.Y(n_399)
);

NAND2x1_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_10),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

AND2x4_ASAP7_75t_SL g75 ( 
.A(n_10),
.B(n_76),
.Y(n_75)
);

NAND2x1p5_ASAP7_75t_L g82 ( 
.A(n_10),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_10),
.B(n_123),
.Y(n_122)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_10),
.B(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_11),
.Y(n_164)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_11),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_12),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_12),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_12),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_12),
.B(n_202),
.Y(n_201)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_13),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_145),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_144),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NOR2xp67_ASAP7_75t_SL g144 ( 
.A(n_19),
.B(n_127),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_95),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_20),
.B(n_70),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_45),
.B1(n_46),
.B2(n_69),
.Y(n_20)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_32),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_22),
.B(n_34),
.C(n_38),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_25),
.C(n_28),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_23),
.B(n_121),
.C(n_125),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_23),
.A2(n_72),
.B1(n_73),
.B2(n_119),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_23),
.B(n_53),
.C(n_66),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_23),
.A2(n_119),
.B1(n_125),
.B2(n_141),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_104),
.C(n_107),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_25),
.A2(n_65),
.B1(n_66),
.B2(n_118),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_25),
.A2(n_66),
.B(n_155),
.C(n_205),
.Y(n_250)
);

AO22x1_ASAP7_75t_L g309 ( 
.A1(n_25),
.A2(n_107),
.B1(n_108),
.B2(n_118),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_38),
.B2(n_44),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_65),
.C(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_38),
.A2(n_44),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_38),
.A2(n_265),
.B(n_267),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_38),
.B(n_265),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_39),
.B(n_106),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_39),
.B(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_43),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_43),
.Y(n_229)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_58),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_47),
.B(n_58),
.C(n_69),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_48),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_48),
.A2(n_122),
.B(n_201),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_48),
.B(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_52),
.A2(n_53),
.B1(n_181),
.B2(n_185),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_52),
.A2(n_53),
.B1(n_139),
.B2(n_140),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_61),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_65),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_53),
.B(n_55),
.C(n_135),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_53),
.A2(n_181),
.B(n_200),
.C(n_205),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_53),
.B(n_181),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_55),
.A2(n_56),
.B1(n_104),
.B2(n_105),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_55),
.B(n_105),
.C(n_159),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_55),
.A2(n_56),
.B1(n_255),
.B2(n_259),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_56),
.B(n_60),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_56),
.B(n_86),
.C(n_255),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_56),
.A2(n_59),
.B(n_68),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_65),
.B(n_68),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_61),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_66),
.B1(n_75),
.B2(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_65),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_65),
.B(n_212),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.C(n_79),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_71),
.B(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_74),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_75),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_75),
.A2(n_122),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_75),
.B(n_122),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_75),
.A2(n_102),
.B1(n_165),
.B2(n_166),
.Y(n_241)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_77),
.Y(n_202)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.C(n_88),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_82),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_81),
.A2(n_82),
.B1(n_226),
.B2(n_230),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_81),
.A2(n_82),
.B1(n_183),
.B2(n_186),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_102),
.C(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_82),
.B(n_184),
.C(n_226),
.Y(n_268)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_86),
.A2(n_114),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_86),
.B(n_125),
.C(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_96),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_115),
.C(n_120),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2x2_ASAP7_75t_L g385 ( 
.A(n_98),
.B(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_111),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_99),
.B(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_102),
.B(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_103),
.B(n_111),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_104),
.A2(n_105),
.B1(n_226),
.B2(n_230),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_104),
.B(n_230),
.C(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_105),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_114),
.B(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_115),
.B(n_120),
.Y(n_386)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_121),
.B(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_122),
.A2(n_162),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_122),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_122),
.B(n_201),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_122),
.A2(n_171),
.B1(n_201),
.B2(n_203),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_123),
.Y(n_266)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_125),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_125),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_125),
.A2(n_141),
.B1(n_319),
.B2(n_323),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_125),
.B(n_317),
.C(n_319),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_125),
.B(n_286),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_143),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_137),
.B2(n_138),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_136),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_141),
.B(n_286),
.C(n_329),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_390),
.B(n_395),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_379),
.Y(n_146)
);

OAI321xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_300),
.A3(n_366),
.B1(n_372),
.B2(n_377),
.C(n_378),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_270),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_243),
.B(n_269),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_220),
.B(n_242),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_197),
.B(n_219),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_173),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_153),
.B(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_161),
.C(n_169),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_155),
.A2(n_159),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_169),
.B1(n_170),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_161),
.A2(n_162),
.B(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_165),
.A2(n_166),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_166),
.B(n_287),
.C(n_291),
.Y(n_317)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_187),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_188),
.C(n_196),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_211),
.B(n_213),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_176),
.A2(n_181),
.B(n_186),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_195),
.B2(n_196),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_192),
.A2(n_239),
.B1(n_254),
.B2(n_260),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_209),
.B(n_218),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_206),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_201),
.A2(n_203),
.B1(n_255),
.B2(n_259),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_201),
.B(n_239),
.C(n_255),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_215),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_214),
.B(n_217),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_222),
.Y(n_242)
);

XOR2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_231),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_231),
.C(n_232),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_226),
.Y(n_230)
);

OR2x6_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_237),
.C(n_241),
.Y(n_247)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_245),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_261),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_248),
.C(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.C(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_252),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_268),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_264),
.C(n_268),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_267),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_271),
.B(n_272),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_283),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_273),
.B(n_284),
.C(n_299),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_281),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_299),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_295),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_297),
.C(n_298),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_353),
.Y(n_300)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_301),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_342),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_302),
.B(n_342),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.C(n_324),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_325),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_304),
.B(n_306),
.C(n_308),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.C(n_314),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_313),
.A2(n_315),
.B1(n_316),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_335),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_333),
.B2(n_334),
.Y(n_326)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_334),
.C(n_335),
.Y(n_343)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.C(n_340),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_345),
.C(n_347),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_348),
.B(n_350),
.C(n_352),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

AOI31xp67_ASAP7_75t_L g372 ( 
.A1(n_353),
.A2(n_367),
.A3(n_373),
.B(n_376),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_356),
.Y(n_353)
);

NOR2x1_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_356),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_361),
.C(n_362),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_357),
.A2(n_358),
.B1(n_362),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_362),
.Y(n_370)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_368),
.B(n_371),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_380),
.Y(n_379)
);

AND2x4_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_382),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_385),
.C(n_387),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_396),
.B(n_397),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_394),
.Y(n_397)
);


endmodule