module fake_jpeg_11000_n_540 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_540);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_20),
.B(n_9),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_54),
.B(n_60),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_56),
.Y(n_159)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_10),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_25),
.B(n_8),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_25),
.B(n_8),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_103),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_101),
.B(n_102),
.Y(n_152)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_24),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_26),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_124),
.B(n_34),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_30),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_126),
.B(n_127),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_30),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_35),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_129),
.B(n_142),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_61),
.A2(n_32),
.B1(n_52),
.B2(n_39),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_138),
.B1(n_156),
.B2(n_45),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_32),
.B1(n_51),
.B2(n_35),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_51),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_52),
.B1(n_36),
.B2(n_46),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_143),
.A2(n_24),
.B1(n_34),
.B2(n_49),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_83),
.A2(n_39),
.B1(n_46),
.B2(n_36),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_153),
.B1(n_24),
.B2(n_56),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_73),
.B(n_48),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_146),
.B(n_154),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_84),
.A2(n_39),
.B1(n_47),
.B2(n_46),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_48),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_67),
.B(n_26),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_161),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_32),
.B1(n_45),
.B2(n_44),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_90),
.B(n_44),
.Y(n_161)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_113),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_175),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_170),
.Y(n_258)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_171),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g273 ( 
.A(n_172),
.B(n_185),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_116),
.A2(n_72),
.B1(n_53),
.B2(n_59),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_173),
.A2(n_199),
.B1(n_58),
.B2(n_80),
.Y(n_255)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_174),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_117),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_177),
.B(n_191),
.Y(n_252)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_119),
.B(n_40),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_180),
.B(n_181),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_24),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_116),
.A2(n_11),
.B(n_18),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_189),
.Y(n_264)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_114),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_132),
.A2(n_87),
.B1(n_86),
.B2(n_47),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_192),
.A2(n_194),
.B1(n_202),
.B2(n_212),
.Y(n_242)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_132),
.A2(n_47),
.B1(n_34),
.B2(n_49),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_197),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_198),
.B(n_201),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_79),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_150),
.C(n_79),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_120),
.A2(n_34),
.B1(n_49),
.B2(n_38),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_106),
.B(n_38),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_204),
.B(n_211),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_106),
.B(n_148),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g257 ( 
.A(n_205),
.B(n_128),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_209),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

BUFx2_ASAP7_75t_SL g212 ( 
.A(n_135),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_38),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_218),
.Y(n_247)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_115),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_220),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_150),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_222),
.B1(n_163),
.B2(n_141),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

OAI22x1_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_130),
.B1(n_141),
.B2(n_144),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_255),
.B1(n_262),
.B2(n_265),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_176),
.B(n_137),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_236),
.B(n_253),
.C(n_269),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_175),
.B1(n_144),
.B2(n_163),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_237),
.A2(n_241),
.B1(n_243),
.B2(n_270),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_195),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_149),
.B1(n_111),
.B2(n_118),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_133),
.B1(n_134),
.B2(n_111),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_101),
.C(n_95),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_257),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_183),
.A2(n_149),
.B1(n_75),
.B2(n_64),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_179),
.B(n_159),
.CI(n_139),
.CON(n_263),
.SN(n_263)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_186),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_167),
.A2(n_82),
.B1(n_63),
.B2(n_118),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_159),
.C(n_128),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_205),
.A2(n_134),
.B1(n_133),
.B2(n_151),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_205),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_288),
.Y(n_335)
);

O2A1O1Ixp33_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_185),
.B(n_208),
.C(n_188),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_276),
.A2(n_320),
.B(n_272),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_247),
.B(n_213),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_280),
.B(n_285),
.Y(n_338)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_282),
.Y(n_357)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_229),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_136),
.B1(n_151),
.B2(n_187),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_289),
.B1(n_307),
.B2(n_309),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_164),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_306),
.C(n_224),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_230),
.A2(n_178),
.B1(n_184),
.B2(n_168),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_318),
.B1(n_319),
.B2(n_227),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_231),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_258),
.A2(n_266),
.B1(n_242),
.B2(n_253),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_290),
.A2(n_293),
.B(n_298),
.Y(n_346)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_209),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_292),
.B(n_301),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_258),
.A2(n_189),
.B1(n_220),
.B2(n_193),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_294),
.Y(n_333)
);

BUFx24_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_257),
.A2(n_171),
.B(n_218),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_315),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_267),
.B(n_206),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_300),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_221),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_238),
.Y(n_302)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_234),
.B(n_215),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_303),
.B(n_304),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_252),
.B(n_197),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_260),
.B(n_136),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_305),
.B(n_232),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_239),
.B(n_182),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_241),
.A2(n_166),
.B1(n_49),
.B2(n_34),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_235),
.Y(n_308)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_270),
.A2(n_49),
.B1(n_41),
.B2(n_2),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_269),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_268),
.B1(n_232),
.B2(n_227),
.Y(n_324)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_263),
.A2(n_8),
.B(n_17),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_312),
.A2(n_316),
.B(n_317),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_263),
.A2(n_262),
.B1(n_250),
.B2(n_259),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_313),
.A2(n_12),
.B(n_16),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_18),
.B(n_7),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_226),
.B(n_240),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_0),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_259),
.A2(n_7),
.B(n_17),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_225),
.A2(n_0),
.B(n_1),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_265),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_225),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_248),
.A2(n_0),
.B(n_2),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_248),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_321),
.B(n_324),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_325),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_284),
.A2(n_223),
.B1(n_226),
.B2(n_251),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_327),
.A2(n_349),
.B(n_358),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_305),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_224),
.C(n_268),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_345),
.C(n_350),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_278),
.A2(n_261),
.B1(n_246),
.B2(n_256),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_344),
.B1(n_347),
.B2(n_277),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_334),
.B(n_298),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_261),
.B1(n_246),
.B2(n_251),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_336),
.A2(n_352),
.B1(n_354),
.B2(n_320),
.Y(n_377)
);

AO21x1_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_283),
.B(n_309),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_313),
.A2(n_244),
.B1(n_249),
.B2(n_245),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_228),
.C(n_244),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_278),
.A2(n_264),
.B1(n_228),
.B2(n_240),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_348),
.A2(n_298),
.B(n_355),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_312),
.A2(n_295),
.B(n_276),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_249),
.C(n_245),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_254),
.B1(n_240),
.B2(n_5),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_299),
.B(n_306),
.C(n_281),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_359),
.C(n_280),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_294),
.A2(n_254),
.B1(n_4),
.B2(n_3),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_293),
.A2(n_254),
.B(n_13),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_355),
.A2(n_316),
.B(n_314),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_276),
.A2(n_12),
.B(n_16),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_3),
.C(n_4),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_362),
.A2(n_317),
.B(n_310),
.Y(n_384)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_364),
.A2(n_397),
.B(n_326),
.Y(n_424)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_366),
.A2(n_378),
.B(n_389),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_338),
.B(n_303),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_367),
.B(n_369),
.Y(n_414)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_297),
.Y(n_370)
);

NAND3xp33_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_371),
.C(n_387),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_297),
.Y(n_371)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_335),
.A2(n_292),
.A3(n_275),
.B1(n_304),
.B2(n_288),
.Y(n_372)
);

XOR2x2_ASAP7_75t_SL g416 ( 
.A(n_372),
.B(n_346),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_323),
.A2(n_287),
.B1(n_274),
.B2(n_318),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_377),
.B1(n_391),
.B2(n_398),
.Y(n_427)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_375),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_361),
.A2(n_298),
.B(n_301),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_379),
.A2(n_394),
.B1(n_390),
.B2(n_324),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_356),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_388),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_392),
.C(n_396),
.Y(n_402)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_322),
.Y(n_383)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_383),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_384),
.A2(n_364),
.B1(n_373),
.B2(n_395),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_385),
.B(n_334),
.Y(n_407)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_322),
.Y(n_386)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_386),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_333),
.B(n_297),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_333),
.B(n_315),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_323),
.A2(n_274),
.B1(n_277),
.B2(n_283),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_291),
.C(n_302),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_282),
.Y(n_393)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_393),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_344),
.A2(n_307),
.B1(n_274),
.B2(n_279),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_360),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_398),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_345),
.B(n_350),
.C(n_328),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_342),
.A2(n_361),
.B(n_349),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_341),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_389),
.A2(n_335),
.B1(n_336),
.B2(n_356),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_400),
.A2(n_401),
.B1(n_426),
.B2(n_429),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_407),
.B(n_385),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_329),
.C(n_330),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_422),
.C(n_397),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_360),
.Y(n_411)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_411),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_380),
.B(n_382),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_418),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_427),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_390),
.A2(n_358),
.B1(n_321),
.B2(n_348),
.Y(n_417)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_417),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_330),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_351),
.Y(n_420)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_346),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_428),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_351),
.C(n_362),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_371),
.B(n_359),
.Y(n_423)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_423),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_424),
.A2(n_366),
.B(n_387),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_389),
.A2(n_352),
.B1(n_354),
.B2(n_326),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_369),
.B(n_385),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_430),
.B(n_411),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_432),
.B(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_376),
.C(n_378),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_451),
.C(n_455),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g436 ( 
.A(n_420),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_453),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_SL g437 ( 
.A(n_421),
.B(n_402),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_437),
.B(n_449),
.Y(n_471)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_438),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_376),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_408),
.B(n_388),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_445),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_373),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_368),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_399),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_419),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_414),
.B(n_367),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_372),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_424),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_383),
.C(n_375),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_452),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_412),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_405),
.A2(n_384),
.B(n_391),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_405),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_386),
.C(n_393),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_459),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_434),
.A2(n_427),
.B1(n_454),
.B2(n_440),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_460),
.A2(n_450),
.B1(n_435),
.B2(n_448),
.Y(n_478)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_431),
.Y(n_463)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_463),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_477),
.Y(n_481)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_466),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_416),
.C(n_404),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_468),
.Y(n_485)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_438),
.A2(n_434),
.B1(n_379),
.B2(n_442),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_470),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_425),
.C(n_400),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_473),
.C(n_475),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_425),
.C(n_399),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_444),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_426),
.C(n_403),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_447),
.A2(n_374),
.B1(n_377),
.B2(n_403),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_476),
.A2(n_455),
.B1(n_451),
.B2(n_394),
.Y(n_479)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_478),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_479),
.A2(n_456),
.B1(n_474),
.B2(n_471),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_461),
.A2(n_419),
.B1(n_409),
.B2(n_410),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_480),
.B(n_494),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_483),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_458),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_460),
.A2(n_462),
.B1(n_459),
.B2(n_473),
.Y(n_486)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_486),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_477),
.A2(n_439),
.B1(n_441),
.B2(n_413),
.Y(n_490)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_490),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_445),
.C(n_446),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_493),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_430),
.C(n_365),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_464),
.B(n_363),
.C(n_410),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_457),
.C(n_464),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_495),
.B(n_497),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_457),
.C(n_475),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_472),
.C(n_467),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_501),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_476),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_503),
.A2(n_508),
.B1(n_478),
.B2(n_490),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_413),
.C(n_409),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_506),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_339),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_479),
.A2(n_339),
.B1(n_357),
.B2(n_340),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_481),
.A2(n_340),
.B(n_357),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_509),
.A2(n_481),
.B(n_491),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_SL g525 ( 
.A1(n_512),
.A2(n_509),
.B(n_503),
.C(n_500),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_508),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_487),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_514),
.A2(n_519),
.B1(n_496),
.B2(n_498),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_502),
.B(n_481),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_515),
.A2(n_516),
.B(n_520),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_SL g516 ( 
.A(n_507),
.B(n_489),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_504),
.B(n_493),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_511),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_488),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_495),
.A2(n_488),
.B(n_357),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_523),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_518),
.B(n_497),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_524),
.B(n_525),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_319),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_527),
.B(n_510),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_528),
.B(n_531),
.C(n_6),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_522),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_6),
.B1(n_7),
.B2(n_14),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_SL g532 ( 
.A1(n_529),
.A2(n_515),
.B(n_514),
.C(n_525),
.Y(n_532)
);

O2A1O1Ixp33_ASAP7_75t_SL g536 ( 
.A1(n_532),
.A2(n_6),
.B(n_15),
.C(n_18),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_533),
.B(n_534),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_536),
.A2(n_532),
.B1(n_15),
.B2(n_4),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_537),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_535),
.C(n_3),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_4),
.Y(n_540)
);


endmodule