module fake_aes_158_n_650 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_650);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_650;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_195;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_20), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_52), .Y(n_78) );
INVxp67_ASAP7_75t_L g79 ( .A(n_63), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_44), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_3), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_13), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_29), .Y(n_83) );
INVx1_ASAP7_75t_SL g84 ( .A(n_32), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_2), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_1), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_68), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_25), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_35), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_64), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_13), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_51), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_14), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_4), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_47), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_1), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_18), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_41), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_8), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_6), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_17), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_39), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_7), .Y(n_103) );
BUFx2_ASAP7_75t_SL g104 ( .A(n_69), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_60), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_19), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_34), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_70), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_45), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_7), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_12), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_26), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_24), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_12), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_59), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_42), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_16), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_5), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_65), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_11), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_89), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_121), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_81), .B(n_0), .Y(n_128) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_78), .A2(n_38), .B(n_75), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_102), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_118), .B(n_0), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_80), .B(n_2), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_106), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_87), .B(n_3), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_102), .B(n_5), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_97), .B(n_43), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_101), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_105), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_108), .Y(n_145) );
INVxp67_ASAP7_75t_L g146 ( .A(n_85), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_110), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_120), .Y(n_154) );
INVxp67_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_86), .A2(n_46), .B(n_74), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_93), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_84), .B(n_40), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_99), .B(n_6), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_100), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_103), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_83), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_82), .Y(n_165) );
INVx3_ASAP7_75t_R g166 ( .A(n_139), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_137), .B(n_99), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_165), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_126), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_146), .A2(n_109), .B1(n_90), .B2(n_92), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_128), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_126), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_126), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_128), .B(n_91), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_126), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_126), .Y(n_178) );
INVx8_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_126), .Y(n_180) );
AND2x6_ASAP7_75t_L g181 ( .A(n_139), .B(n_117), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_133), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_164), .B(n_91), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_155), .B(n_96), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_124), .B(n_113), .Y(n_188) );
OR2x2_ASAP7_75t_SL g189 ( .A(n_160), .B(n_112), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_127), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_124), .B(n_107), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_164), .B(n_77), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_164), .B(n_96), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_141), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_164), .B(n_77), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_164), .B(n_107), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_127), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_152), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_138), .B(n_116), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_133), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_138), .B(n_79), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_130), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_130), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_158), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_152), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_125), .B(n_111), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_125), .B(n_109), .Y(n_210) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_157), .A2(n_104), .B(n_50), .Y(n_211) );
INVxp67_ASAP7_75t_SL g212 ( .A(n_131), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_140), .B(n_92), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_133), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_140), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_133), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_141), .Y(n_217) );
OR2x6_ASAP7_75t_L g218 ( .A(n_157), .B(n_104), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_152), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_156), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_148), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_156), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_208), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_212), .B(n_145), .Y(n_225) );
INVx5_ASAP7_75t_L g226 ( .A(n_179), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_213), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_208), .Y(n_228) );
AND2x4_ASAP7_75t_SL g229 ( .A(n_213), .B(n_90), .Y(n_229) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_181), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_208), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_219), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_219), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_215), .B(n_147), .Y(n_234) );
OR2x2_ASAP7_75t_L g235 ( .A(n_168), .B(n_163), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_219), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_173), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_215), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_196), .B(n_156), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_220), .Y(n_240) );
AND2x6_ASAP7_75t_SL g241 ( .A(n_213), .B(n_132), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_220), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_181), .A2(n_147), .B1(n_145), .B2(n_154), .Y(n_243) );
BUFx3_ASAP7_75t_L g244 ( .A(n_179), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_196), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_172), .A2(n_112), .B1(n_163), .B2(n_162), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_200), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_170), .Y(n_248) );
BUFx4f_ASAP7_75t_L g249 ( .A(n_181), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_169), .A2(n_154), .B1(n_162), .B2(n_158), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_223), .B(n_156), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_209), .B(n_161), .Y(n_252) );
AOI22xp33_ASAP7_75t_SL g253 ( .A1(n_176), .A2(n_141), .B1(n_136), .B2(n_153), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_183), .B(n_144), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_167), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_185), .Y(n_256) );
NOR2xp67_ASAP7_75t_L g257 ( .A(n_190), .B(n_143), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_176), .B(n_161), .Y(n_258) );
INVx5_ASAP7_75t_L g259 ( .A(n_179), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_205), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_185), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_191), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_179), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_181), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_209), .B(n_143), .Y(n_265) );
BUFx5_ASAP7_75t_L g266 ( .A(n_181), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_205), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_206), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_200), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_196), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_167), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_196), .B(n_217), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_209), .B(n_144), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_221), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_196), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_221), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_194), .B(n_142), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_190), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_191), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_190), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_194), .B(n_142), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_181), .A2(n_191), .B1(n_188), .B2(n_169), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_199), .Y(n_285) );
OR2x2_ASAP7_75t_SL g286 ( .A(n_189), .B(n_129), .Y(n_286) );
INVx4_ASAP7_75t_L g287 ( .A(n_226), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_225), .Y(n_288) );
INVx3_ASAP7_75t_L g289 ( .A(n_226), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_237), .B(n_204), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_284), .A2(n_167), .B1(n_217), .B2(n_189), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_251), .A2(n_239), .B(n_242), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_225), .Y(n_293) );
BUFx4f_ASAP7_75t_L g294 ( .A(n_227), .Y(n_294) );
AOI21xp33_ASAP7_75t_L g295 ( .A1(n_238), .A2(n_198), .B(n_197), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_229), .B(n_188), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_240), .A2(n_129), .B(n_192), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_226), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_226), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_239), .A2(n_218), .B(n_197), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_259), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_225), .B(n_188), .Y(n_302) );
NAND2x1_ASAP7_75t_SL g303 ( .A(n_256), .B(n_129), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_259), .Y(n_304) );
AND2x2_ASAP7_75t_SL g305 ( .A(n_230), .B(n_129), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_259), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_235), .B(n_191), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_254), .A2(n_207), .B(n_201), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_259), .B(n_191), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_244), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_234), .B(n_191), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_248), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_244), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_243), .A2(n_218), .B1(n_166), .B2(n_199), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_229), .B(n_199), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_248), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_263), .Y(n_317) );
INVx4_ASAP7_75t_L g318 ( .A(n_263), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_258), .Y(n_319) );
INVx4_ASAP7_75t_SL g320 ( .A(n_264), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_264), .Y(n_321) );
BUFx10_ASAP7_75t_L g322 ( .A(n_241), .Y(n_322) );
BUFx2_ASAP7_75t_SL g323 ( .A(n_266), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_230), .Y(n_324) );
INVx4_ASAP7_75t_L g325 ( .A(n_230), .Y(n_325) );
BUFx4_ASAP7_75t_SL g326 ( .A(n_281), .Y(n_326) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_249), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_240), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_255), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_261), .B(n_166), .Y(n_330) );
NAND2x1_ASAP7_75t_L g331 ( .A(n_255), .B(n_141), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_255), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_278), .A2(n_218), .B1(n_141), .B2(n_153), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_246), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_252), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_252), .B(n_149), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_302), .B(n_252), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_328), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_302), .A2(n_243), .B1(n_286), .B2(n_253), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_328), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_334), .A2(n_249), .B1(n_265), .B2(n_274), .Y(n_341) );
CKINVDCx6p67_ASAP7_75t_R g342 ( .A(n_312), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_316), .A2(n_249), .B1(n_281), .B2(n_250), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_297), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_319), .A2(n_279), .B1(n_262), .B2(n_218), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_302), .A2(n_271), .B1(n_283), .B2(n_254), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_290), .B(n_260), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_299), .B(n_266), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_288), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g350 ( .A1(n_294), .A2(n_283), .B1(n_271), .B2(n_257), .C(n_231), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_307), .A2(n_268), .B1(n_272), .B2(n_267), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_293), .B(n_271), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_329), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_294), .A2(n_232), .B1(n_224), .B2(n_228), .Y(n_354) );
BUFx2_ASAP7_75t_SL g355 ( .A(n_299), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_296), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_299), .Y(n_357) );
INVxp33_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
AOI332xp33_ASAP7_75t_L g359 ( .A1(n_336), .A2(n_135), .A3(n_134), .B1(n_149), .B2(n_282), .B3(n_280), .C1(n_285), .C2(n_9), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_299), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_332), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_331), .A2(n_273), .B(n_275), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_292), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_307), .B(n_232), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_301), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_335), .B(n_232), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_308), .B(n_266), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_291), .A2(n_228), .B1(n_224), .B2(n_233), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_339), .A2(n_333), .B1(n_314), .B2(n_311), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g370 ( .A1(n_359), .A2(n_330), .B(n_134), .C(n_135), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_339), .A2(n_322), .B1(n_330), .B2(n_309), .Y(n_371) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_359), .A2(n_295), .B(n_303), .C(n_300), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_365), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_347), .B(n_322), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_347), .A2(n_285), .B1(n_236), .B2(n_233), .C(n_310), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_356), .A2(n_327), .B1(n_287), .B2(n_310), .C(n_313), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_367), .A2(n_322), .B1(n_309), .B2(n_318), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_358), .B(n_313), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_342), .A2(n_318), .B1(n_287), .B2(n_301), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_342), .Y(n_380) );
AOI22x1_ASAP7_75t_SL g381 ( .A1(n_349), .A2(n_287), .B1(n_289), .B2(n_326), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_351), .A2(n_305), .B1(n_317), .B2(n_327), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_337), .B(n_289), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g385 ( .A1(n_346), .A2(n_317), .B1(n_236), .B2(n_306), .C(n_298), .Y(n_385) );
OR2x6_ASAP7_75t_L g386 ( .A(n_355), .B(n_301), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_367), .A2(n_309), .B1(n_141), .B2(n_306), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_351), .A2(n_141), .B1(n_298), .B2(n_301), .Y(n_388) );
OAI221xp5_ASAP7_75t_SL g389 ( .A1(n_341), .A2(n_277), .B1(n_269), .B2(n_247), .C(n_326), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
OAI332xp33_ASAP7_75t_L g391 ( .A1(n_350), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_14), .B3(n_15), .C1(n_203), .C2(n_193), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_365), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_353), .Y(n_394) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_364), .A2(n_297), .B(n_305), .C(n_247), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_345), .A2(n_323), .B1(n_304), .B2(n_325), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_386), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_371), .A2(n_343), .B1(n_354), .B2(n_361), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_389), .A2(n_340), .B1(n_338), .B2(n_366), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_393), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_382), .A2(n_361), .B1(n_363), .B2(n_366), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_386), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_386), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_382), .B(n_355), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_369), .A2(n_338), .B1(n_340), .B2(n_352), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_380), .A2(n_340), .B1(n_338), .B2(n_304), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_394), .B(n_357), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_383), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
OAI211xp5_ASAP7_75t_SL g411 ( .A1(n_370), .A2(n_368), .B(n_363), .C(n_203), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_373), .B(n_357), .Y(n_413) );
OAI33xp33_ASAP7_75t_L g414 ( .A1(n_379), .A2(n_193), .A3(n_184), .B1(n_187), .B2(n_214), .B3(n_202), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_390), .B(n_360), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_390), .B(n_360), .Y(n_416) );
AOI21xp5_ASAP7_75t_SL g417 ( .A1(n_396), .A2(n_325), .B(n_304), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_372), .A2(n_362), .B(n_344), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_392), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_369), .A2(n_211), .B1(n_304), .B2(n_159), .Y(n_420) );
NAND4xp25_ASAP7_75t_SL g421 ( .A(n_377), .B(n_10), .C(n_15), .D(n_344), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_392), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_392), .B(n_211), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_384), .B(n_211), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_159), .B1(n_325), .B2(n_344), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_375), .B(n_151), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_391), .A2(n_187), .B1(n_184), .B2(n_151), .C(n_148), .Y(n_427) );
OAI33xp33_ASAP7_75t_L g428 ( .A1(n_381), .A2(n_202), .A3(n_175), .B1(n_178), .B2(n_222), .B3(n_214), .Y(n_428) );
NAND4xp25_ASAP7_75t_L g429 ( .A(n_378), .B(n_178), .C(n_174), .D(n_222), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_376), .A2(n_148), .B1(n_151), .B2(n_269), .C(n_277), .Y(n_430) );
AOI31xp33_ASAP7_75t_L g431 ( .A1(n_399), .A2(n_388), .A3(n_387), .B(n_385), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_409), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_412), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_401), .B(n_395), .Y(n_434) );
NOR2x1_ASAP7_75t_SL g435 ( .A(n_405), .B(n_403), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
INVx5_ASAP7_75t_SL g437 ( .A(n_405), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_418), .A2(n_348), .B(n_180), .Y(n_438) );
AND2x2_ASAP7_75t_SL g439 ( .A(n_402), .B(n_324), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_409), .B(n_159), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_424), .B(n_151), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_410), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_405), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_424), .B(n_151), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_397), .Y(n_445) );
OAI31xp33_ASAP7_75t_L g446 ( .A1(n_421), .A2(n_273), .A3(n_180), .B(n_175), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_405), .B(n_404), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_408), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
OR2x6_ASAP7_75t_L g451 ( .A(n_417), .B(n_321), .Y(n_451) );
AND2x4_ASAP7_75t_SL g452 ( .A(n_397), .B(n_321), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_408), .B(n_423), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_427), .B(n_174), .C(n_151), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_423), .B(n_148), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_411), .A2(n_159), .B1(n_321), .B2(n_266), .Y(n_457) );
AO22x2_ASAP7_75t_L g458 ( .A1(n_397), .A2(n_320), .B1(n_159), .B2(n_321), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_398), .A2(n_159), .B1(n_266), .B2(n_324), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_413), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_419), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_404), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_422), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_422), .B(n_148), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
INVx6_ASAP7_75t_L g466 ( .A(n_416), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_403), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_430), .B(n_148), .C(n_186), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_416), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_415), .Y(n_470) );
OAI211xp5_ASAP7_75t_L g471 ( .A1(n_417), .A2(n_324), .B(n_186), .C(n_216), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_415), .B(n_21), .Y(n_472) );
AND2x4_ASAP7_75t_SL g473 ( .A(n_426), .B(n_324), .Y(n_473) );
INVx5_ASAP7_75t_L g474 ( .A(n_426), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_428), .A2(n_186), .B1(n_171), .B2(n_177), .C(n_216), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_400), .B(n_22), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_420), .B(n_23), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
AOI221x1_ASAP7_75t_L g479 ( .A1(n_458), .A2(n_429), .B1(n_414), .B2(n_407), .C(n_425), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_442), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_453), .B(n_27), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_433), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_453), .B(n_28), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_435), .B(n_30), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_470), .B(n_31), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_448), .B(n_33), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_469), .B(n_159), .Y(n_489) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_467), .B(n_216), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_436), .Y(n_492) );
AOI31xp33_ASAP7_75t_L g493 ( .A1(n_447), .A2(n_320), .A3(n_36), .B(n_37), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_466), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_442), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_466), .Y(n_496) );
OAI211xp5_ASAP7_75t_L g497 ( .A1(n_443), .A2(n_216), .B(n_195), .C(n_186), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_465), .B(n_216), .C(n_195), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_441), .B(n_48), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_441), .B(n_49), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_456), .B(n_53), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_444), .B(n_54), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_444), .B(n_55), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_448), .B(n_56), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_467), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_450), .B(n_447), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_455), .Y(n_507) );
BUFx2_ASAP7_75t_SL g508 ( .A(n_467), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_460), .B(n_57), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_466), .B(n_58), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_454), .A2(n_266), .B1(n_320), .B2(n_177), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_439), .A2(n_266), .B1(n_177), .B2(n_195), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_450), .B(n_461), .Y(n_513) );
XNOR2xp5_ASAP7_75t_L g514 ( .A(n_439), .B(n_61), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_461), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_463), .B(n_62), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_434), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_452), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_464), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_443), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_465), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_437), .B(n_66), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_462), .B(n_472), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_437), .B(n_67), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_464), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_478), .Y(n_527) );
OAI21x1_ASAP7_75t_L g528 ( .A1(n_490), .A2(n_445), .B(n_475), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_492), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_491), .B(n_431), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_493), .A2(n_473), .B(n_446), .C(n_476), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_506), .B(n_437), .Y(n_532) );
NOR3xp33_ASAP7_75t_SL g533 ( .A(n_514), .B(n_471), .C(n_468), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_505), .B(n_474), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_487), .Y(n_535) );
OAI31xp33_ASAP7_75t_L g536 ( .A1(n_514), .A2(n_473), .A3(n_476), .B(n_477), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_518), .B(n_474), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_494), .B(n_437), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_487), .B(n_435), .Y(n_539) );
AOI221xp5_ASAP7_75t_SL g540 ( .A1(n_496), .A2(n_477), .B1(n_459), .B2(n_457), .C(n_171), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_508), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_484), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_518), .B(n_474), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_482), .B(n_474), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_522), .B(n_451), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_497), .A2(n_451), .B(n_458), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_513), .B(n_452), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_521), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_482), .B(n_438), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_480), .Y(n_550) );
NAND2x1_ASAP7_75t_L g551 ( .A(n_505), .B(n_451), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_495), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_521), .B(n_451), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_505), .B(n_438), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_485), .B(n_440), .Y(n_555) );
BUFx8_ASAP7_75t_SL g556 ( .A(n_485), .Y(n_556) );
OAI22xp33_ASAP7_75t_L g557 ( .A1(n_488), .A2(n_458), .B1(n_438), .B2(n_76), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_513), .B(n_458), .Y(n_558) );
AOI211xp5_ASAP7_75t_L g559 ( .A1(n_481), .A2(n_186), .B(n_195), .C(n_171), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_515), .B(n_71), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_479), .A2(n_72), .B(n_171), .Y(n_561) );
AOI211x1_ASAP7_75t_SL g562 ( .A1(n_524), .A2(n_171), .B(n_177), .C(n_182), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_516), .B(n_177), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_520), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_526), .B(n_182), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_508), .Y(n_566) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_541), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_527), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_531), .A2(n_498), .B(n_485), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_541), .B(n_519), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_564), .B(n_526), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_564), .B(n_507), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_548), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_542), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_548), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_531), .A2(n_483), .B1(n_481), .B2(n_512), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_550), .Y(n_577) );
AOI32xp33_ASAP7_75t_L g578 ( .A1(n_530), .A2(n_523), .A3(n_519), .B1(n_500), .B2(n_503), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_552), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_530), .B(n_507), .Y(n_580) );
XOR2x2_ASAP7_75t_L g581 ( .A(n_556), .B(n_523), .Y(n_581) );
AO21x1_ASAP7_75t_L g582 ( .A1(n_536), .A2(n_525), .B(n_504), .Y(n_582) );
XNOR2x1_ASAP7_75t_L g583 ( .A(n_532), .B(n_525), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_566), .A2(n_479), .B(n_500), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_535), .B(n_566), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_545), .B(n_509), .Y(n_586) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_561), .A2(n_486), .B1(n_503), .B2(n_502), .C1(n_499), .C2(n_501), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_553), .B(n_517), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_553), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_547), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_537), .Y(n_591) );
AOI31xp33_ASAP7_75t_L g592 ( .A1(n_534), .A2(n_502), .A3(n_510), .B(n_517), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_538), .B(n_511), .Y(n_593) );
NOR2xp67_ASAP7_75t_L g594 ( .A(n_546), .B(n_489), .Y(n_594) );
O2A1O1Ixp5_ASAP7_75t_L g595 ( .A1(n_551), .A2(n_182), .B(n_195), .C(n_245), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_539), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_563), .Y(n_597) );
XNOR2x1_ASAP7_75t_L g598 ( .A(n_539), .B(n_534), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_559), .B(n_245), .Y(n_599) );
AO22x1_ASAP7_75t_L g600 ( .A1(n_544), .A2(n_245), .B1(n_270), .B2(n_276), .Y(n_600) );
OAI22xp5_ASAP7_75t_SL g601 ( .A1(n_554), .A2(n_245), .B1(n_270), .B2(n_276), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_558), .B(n_270), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_533), .A2(n_270), .B1(n_276), .B2(n_557), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_543), .A2(n_276), .B1(n_557), .B2(n_554), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_549), .Y(n_605) );
NAND3xp33_ASAP7_75t_SL g606 ( .A(n_533), .B(n_562), .C(n_543), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g607 ( .A1(n_555), .A2(n_560), .B1(n_540), .B2(n_565), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_555), .B(n_528), .Y(n_608) );
OAI322xp33_ASAP7_75t_L g609 ( .A1(n_530), .A2(n_527), .A3(n_478), .B1(n_491), .B2(n_506), .C1(n_552), .C2(n_550), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_530), .A2(n_527), .B1(n_478), .B2(n_491), .C(n_391), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_527), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_527), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_529), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_599), .Y(n_614) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_567), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_591), .B(n_575), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_598), .A2(n_569), .B(n_581), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
AND3x4_ASAP7_75t_L g619 ( .A(n_594), .B(n_582), .C(n_596), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_584), .B(n_606), .C(n_603), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_571), .B(n_572), .Y(n_621) );
AOI322xp5_ASAP7_75t_L g622 ( .A1(n_610), .A2(n_567), .A3(n_608), .B1(n_570), .B2(n_585), .C1(n_607), .C2(n_580), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_589), .B(n_605), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_SL g624 ( .A1(n_570), .A2(n_569), .B(n_576), .C(n_585), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_574), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_606), .A2(n_590), .B1(n_593), .B2(n_583), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_568), .B(n_612), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_624), .A2(n_617), .B(n_619), .Y(n_628) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_614), .A2(n_603), .B(n_586), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_627), .Y(n_630) );
NAND4xp75_ASAP7_75t_L g631 ( .A(n_622), .B(n_610), .C(n_604), .D(n_595), .Y(n_631) );
NOR4xp75_ASAP7_75t_SL g632 ( .A(n_622), .B(n_588), .C(n_609), .D(n_578), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_627), .Y(n_633) );
OAI211xp5_ASAP7_75t_SL g634 ( .A1(n_626), .A2(n_587), .B(n_611), .C(n_595), .Y(n_634) );
XNOR2xp5_ASAP7_75t_L g635 ( .A(n_620), .B(n_577), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_630), .Y(n_636) );
AO22x2_ASAP7_75t_L g637 ( .A1(n_631), .A2(n_615), .B1(n_618), .B2(n_616), .Y(n_637) );
NAND5xp2_ASAP7_75t_L g638 ( .A(n_628), .B(n_586), .C(n_623), .D(n_602), .E(n_597), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_633), .Y(n_639) );
NOR3xp33_ASAP7_75t_SL g640 ( .A(n_628), .B(n_601), .C(n_614), .Y(n_640) );
OR3x1_ASAP7_75t_L g641 ( .A(n_638), .B(n_632), .C(n_634), .Y(n_641) );
NAND3xp33_ASAP7_75t_SL g642 ( .A(n_640), .B(n_635), .C(n_629), .Y(n_642) );
AOI31xp33_ASAP7_75t_L g643 ( .A1(n_637), .A2(n_621), .A3(n_579), .B(n_614), .Y(n_643) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_641), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_643), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_644), .A2(n_637), .B1(n_639), .B2(n_636), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_645), .B(n_642), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_647), .A2(n_625), .B1(n_592), .B2(n_613), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_648), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_649), .A2(n_646), .B(n_600), .Y(n_650) );
endmodule