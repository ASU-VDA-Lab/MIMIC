module fake_jpeg_3585_n_398 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_398);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_398;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_20),
.Y(n_58)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_7),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_60),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_22),
.B(n_42),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_7),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_63),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_6),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_68),
.Y(n_131)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_6),
.B(n_1),
.Y(n_67)
);

OR2x2_ASAP7_75t_SL g159 ( 
.A(n_67),
.B(n_32),
.Y(n_159)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_30),
.B(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_69),
.B(n_75),
.Y(n_149)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_70),
.Y(n_179)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_39),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g167 ( 
.A(n_72),
.Y(n_167)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_73),
.Y(n_174)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_30),
.B(n_3),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g177 ( 
.A(n_78),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_79),
.B(n_80),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_82),
.B(n_83),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_5),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_106),
.Y(n_137)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_31),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_92),
.B(n_93),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_13),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_24),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_31),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_102),
.B(n_105),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_14),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_45),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_36),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_46),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_113),
.B(n_145),
.C(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_38),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_115),
.B(n_126),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_118),
.B(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_84),
.B(n_38),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_55),
.A2(n_46),
.B1(n_27),
.B2(n_29),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_142),
.A2(n_130),
.B1(n_136),
.B2(n_128),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_65),
.A2(n_40),
.B1(n_52),
.B2(n_50),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_180),
.B1(n_181),
.B2(n_100),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_29),
.C(n_53),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_56),
.A2(n_40),
.B1(n_52),
.B2(n_50),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_157),
.B1(n_160),
.B2(n_165),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_54),
.A2(n_36),
.B1(n_49),
.B2(n_48),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_152),
.A2(n_150),
.B1(n_156),
.B2(n_125),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_161),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_57),
.A2(n_33),
.B1(n_49),
.B2(n_48),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_81),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_76),
.B(n_53),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_85),
.A2(n_44),
.B1(n_15),
.B2(n_16),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_96),
.B(n_15),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_113),
.Y(n_200)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_61),
.Y(n_173)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_90),
.A2(n_0),
.B1(n_16),
.B2(n_110),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_145),
.B1(n_166),
.B2(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_91),
.B(n_0),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_133),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_74),
.A2(n_96),
.B1(n_71),
.B2(n_77),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_87),
.A2(n_111),
.B1(n_86),
.B2(n_101),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_117),
.B(n_70),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_184),
.B(n_186),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_94),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_185),
.B(n_187),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_73),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_115),
.A2(n_94),
.B(n_103),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_188),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_202),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_131),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_192),
.B(n_200),
.Y(n_254)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_195),
.A2(n_225),
.B1(n_242),
.B2(n_190),
.Y(n_271)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_137),
.B(n_122),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_198),
.B(n_207),
.Y(n_283)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_199),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_164),
.C(n_126),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_122),
.B(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_208),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_176),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_209),
.B(n_215),
.Y(n_277)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_SL g212 ( 
.A(n_149),
.B(n_144),
.C(n_175),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_213),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_142),
.A2(n_127),
.B1(n_129),
.B2(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_214),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_134),
.B(n_141),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_226),
.Y(n_243)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_114),
.A2(n_116),
.B1(n_124),
.B2(n_163),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_213),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_149),
.A2(n_119),
.B1(n_153),
.B2(n_120),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_143),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_235),
.Y(n_269)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_227),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_181),
.A2(n_168),
.B1(n_154),
.B2(n_170),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_132),
.B(n_139),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_121),
.B(n_177),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_123),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_229),
.Y(n_257)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_231),
.Y(n_261)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_232),
.Y(n_284)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_117),
.B(n_115),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_115),
.B(n_126),
.Y(n_235)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_156),
.A2(n_142),
.B(n_97),
.C(n_145),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_188),
.B(n_233),
.C(n_216),
.Y(n_275)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_158),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_238),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_122),
.B(n_117),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_131),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_240),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_155),
.B(n_117),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_122),
.B(n_117),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_241),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_175),
.A2(n_115),
.B1(n_178),
.B2(n_126),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_234),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_246),
.B(n_247),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_196),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_209),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_230),
.Y(n_296)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_253),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_255),
.A2(n_280),
.B1(n_264),
.B2(n_244),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_185),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_276),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_221),
.A2(n_242),
.B1(n_206),
.B2(n_187),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_264),
.A2(n_277),
.B1(n_246),
.B2(n_272),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_271),
.A2(n_274),
.B1(n_280),
.B2(n_253),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_191),
.A2(n_236),
.B1(n_188),
.B2(n_229),
.Y(n_274)
);

HAxp5_ASAP7_75t_SL g314 ( 
.A(n_275),
.B(n_256),
.CON(n_314),
.SN(n_314)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_216),
.B(n_205),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_199),
.B(n_231),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_279),
.B(n_281),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_211),
.B(n_194),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_188),
.B(n_201),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_286),
.A2(n_287),
.B(n_300),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_245),
.A2(n_225),
.B1(n_201),
.B2(n_223),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_252),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_292),
.Y(n_325)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_289),
.Y(n_333)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_232),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_290),
.B(n_296),
.Y(n_319)
);

OAI31xp33_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_217),
.A3(n_223),
.B(n_197),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_SL g330 ( 
.A1(n_291),
.A2(n_314),
.B(n_262),
.C(n_268),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_279),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_303),
.Y(n_326)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_294),
.Y(n_320)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_260),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_298),
.B(n_311),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_265),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_299),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_269),
.A2(n_249),
.B(n_243),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_301),
.A2(n_282),
.B1(n_267),
.B2(n_278),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_302),
.A2(n_307),
.B1(n_309),
.B2(n_266),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_247),
.B(n_269),
.C(n_243),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_308),
.C(n_262),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_254),
.B(n_271),
.C(n_259),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_249),
.A2(n_283),
.B1(n_256),
.B2(n_259),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_250),
.B(n_285),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_273),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_313),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_276),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_266),
.B(n_265),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_315),
.B(n_268),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_248),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_318),
.A2(n_287),
.B1(n_295),
.B2(n_316),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_267),
.Y(n_323)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_282),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_330),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_270),
.B(n_248),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_327),
.A2(n_331),
.B(n_334),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_306),
.Y(n_342)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_286),
.A2(n_308),
.B(n_305),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_337),
.C(n_325),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_310),
.B(n_301),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_310),
.A2(n_303),
.B(n_313),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_325),
.A2(n_291),
.B1(n_293),
.B2(n_290),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_339),
.A2(n_345),
.B1(n_330),
.B2(n_320),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_295),
.B1(n_304),
.B2(n_306),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_340),
.A2(n_348),
.B1(n_327),
.B2(n_322),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_312),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_347),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_343),
.C(n_344),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_298),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_317),
.C(n_295),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_297),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_333),
.A2(n_294),
.B1(n_311),
.B2(n_337),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_323),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_349),
.B(n_351),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_326),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_321),
.B(n_326),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_319),
.C(n_338),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_343),
.C(n_344),
.Y(n_359)
);

AO21x1_ASAP7_75t_L g370 ( 
.A1(n_356),
.A2(n_368),
.B(n_338),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_363),
.Y(n_375)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_348),
.Y(n_360)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_352),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_319),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_352),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_364),
.B(n_336),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_365),
.B(n_367),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_318),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_366),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_340),
.B(n_321),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_368),
.A2(n_353),
.B1(n_346),
.B2(n_355),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_373),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_357),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_324),
.Y(n_374)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_374),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_320),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_372),
.A2(n_365),
.B(n_358),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_378),
.B(n_379),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_358),
.B(n_359),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_382),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_373),
.B(n_361),
.Y(n_383)
);

INVx11_ASAP7_75t_L g385 ( 
.A(n_383),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_375),
.C(n_363),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_386),
.B(n_387),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_375),
.C(n_376),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_376),
.B1(n_356),
.B2(n_369),
.Y(n_389)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_387),
.Y(n_390)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_390),
.A2(n_391),
.B(n_388),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_386),
.B(n_370),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_394),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_392),
.C(n_384),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_395),
.A2(n_396),
.B(n_384),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_397),
.B(n_391),
.Y(n_398)
);


endmodule