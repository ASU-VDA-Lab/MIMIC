module fake_jpeg_13160_n_194 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_194);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_13),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_70),
.Y(n_91)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_3),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_85),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_79),
.B1(n_63),
.B2(n_61),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_94),
.B(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_62),
.B1(n_70),
.B2(n_56),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_64),
.B1(n_55),
.B2(n_73),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_99),
.B1(n_68),
.B2(n_58),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_57),
.B1(n_54),
.B2(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_58),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_100),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_52),
.Y(n_131)
);

NOR2xp67_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_76),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_96),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_114),
.Y(n_133)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_122),
.Y(n_134)
);

BUFx2_ASAP7_75t_SL g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_7),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_4),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_82),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_81),
.B(n_78),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_135)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_131),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_40),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_5),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_27),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_7),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_142),
.B1(n_134),
.B2(n_143),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_115),
.B1(n_123),
.B2(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_8),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_22),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_9),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_10),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_11),
.B(n_14),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_35),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_155),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_153),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_15),
.B(n_21),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_159),
.B(n_166),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_24),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_160),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_29),
.B(n_31),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_32),
.A3(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_38),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_167),
.B(n_168),
.Y(n_170)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_126),
.B(n_132),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_171),
.B1(n_149),
.B2(n_160),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_147),
.B1(n_146),
.B2(n_46),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_159),
.B(n_165),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_151),
.B1(n_162),
.B2(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_182),
.B(n_184),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_175),
.C(n_178),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_41),
.B1(n_43),
.B2(n_49),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_180),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_185),
.B(n_174),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_186),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_184),
.B(n_176),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_170),
.B(n_175),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_179),
.Y(n_194)
);


endmodule