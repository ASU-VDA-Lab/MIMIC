module fake_jpeg_12440_n_146 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_2),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_30),
.B(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_10),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_12),
.B(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_18),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_15),
.Y(n_70)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_12),
.B(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_48),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_20),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_11),
.Y(n_50)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_24),
.B(n_14),
.C(n_28),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_70),
.B(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_11),
.B1(n_28),
.B2(n_16),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_74),
.B(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_31),
.A2(n_11),
.B1(n_14),
.B2(n_16),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_74),
.B1(n_40),
.B2(n_32),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_25),
.B(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_65),
.B(n_71),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_15),
.B1(n_20),
.B2(n_25),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_73),
.B(n_53),
.C(n_63),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_37),
.A2(n_4),
.B1(n_0),
.B2(n_1),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_33),
.B1(n_45),
.B2(n_32),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_48),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_87),
.B1(n_90),
.B2(n_94),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_48),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_59),
.C(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_79),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_83),
.Y(n_98)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_60),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_54),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_93),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_52),
.B(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_111),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_52),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_79),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_94),
.B(n_87),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_119),
.A2(n_121),
.B(n_110),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_101),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_80),
.B1(n_87),
.B2(n_88),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_121),
.B(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_109),
.C(n_103),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_126),
.B(n_129),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_108),
.C(n_97),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_127),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_105),
.C(n_87),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_86),
.B(n_134),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_112),
.B1(n_116),
.B2(n_105),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_135),
.B1(n_125),
.B2(n_105),
.Y(n_136)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_126),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_138),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_142),
.A2(n_143),
.B(n_140),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_135),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_144),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_133),
.Y(n_146)
);


endmodule