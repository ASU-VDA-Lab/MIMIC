module fake_jpeg_11403_n_171 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_171);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_25),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_30),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_63),
.Y(n_93)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_53),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_72),
.B1(n_64),
.B2(n_58),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_95),
.B(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_72),
.B1(n_70),
.B2(n_56),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_92),
.B1(n_75),
.B2(n_82),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_67),
.B1(n_65),
.B2(n_54),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_69),
.B(n_54),
.C(n_62),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_116),
.B(n_1),
.Y(n_120)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_109),
.B1(n_113),
.B2(n_114),
.Y(n_130)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_110),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_73),
.B1(n_71),
.B2(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_51),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_115),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_62),
.B1(n_52),
.B2(n_3),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_15),
.B1(n_47),
.B2(n_46),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_2),
.C(n_3),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_50),
.B(n_44),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_11),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_120),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_41),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_126),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_127),
.Y(n_152)
);

CKINVDCx10_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_39),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_132),
.B1(n_136),
.B2(n_17),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_135),
.B1(n_126),
.B2(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_7),
.B(n_8),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_19),
.B(n_20),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_24),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_142),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_13),
.B(n_14),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_141),
.B(n_149),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_13),
.B(n_14),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_138),
.B(n_122),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_159),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.C(n_35),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_160),
.B(n_140),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_148),
.C(n_152),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_148),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_166),
.B(n_141),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_162),
.B(n_164),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_143),
.B1(n_153),
.B2(n_147),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_158),
.B(n_146),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);


endmodule