module fake_jpeg_13717_n_48 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_48);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_48;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_0),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_20),
.A2(n_21),
.B1(n_17),
.B2(n_11),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_20),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_32),
.B(n_33),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_26),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_38),
.C(n_34),
.Y(n_39)
);

A2O1A1O1Ixp25_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_24),
.B(n_18),
.C(n_17),
.D(n_10),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_28),
.B(n_16),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_33),
.C(n_6),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_4),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_42),
.C(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_32),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_46),
.A2(n_44),
.B(n_28),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_4),
.Y(n_48)
);


endmodule