module fake_ariane_2810_n_1753 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1753);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1753;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1733;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_SL g173 ( 
.A(n_162),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_21),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_60),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_42),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_171),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_18),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_129),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_80),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_88),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_81),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_46),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_99),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_4),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_25),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_54),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_83),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_100),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_61),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_57),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_105),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_21),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_96),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_51),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_67),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_141),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_45),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_90),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_98),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_137),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_35),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_94),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_86),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_166),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_27),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_26),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_170),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_6),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_32),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_14),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_118),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_4),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_24),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_66),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_106),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_26),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_138),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_12),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_164),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_156),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_44),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_69),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_38),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_42),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_48),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_120),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_124),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_115),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_116),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_133),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_65),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_50),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_72),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_0),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_91),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_25),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_145),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_23),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_114),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_49),
.Y(n_264)
);

BUFx2_ASAP7_75t_SL g265 ( 
.A(n_123),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_19),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_1),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_110),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_46),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_79),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_35),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_107),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_82),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_132),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_11),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_32),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_14),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_1),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_30),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_37),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_165),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_15),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_126),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_39),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_31),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_150),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_64),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_48),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_155),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_55),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_76),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_104),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_37),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_160),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_9),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_6),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_63),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_92),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_49),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_5),
.Y(n_305)
);

BUFx2_ASAP7_75t_SL g306 ( 
.A(n_27),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_36),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_12),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_73),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_13),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_59),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_97),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_29),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_40),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_158),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_8),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_93),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_22),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_28),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_50),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_40),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_101),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_172),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_117),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_53),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_119),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_23),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_68),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_78),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_70),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_95),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_108),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_134),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_154),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_28),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_41),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_153),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_102),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_45),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_58),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_10),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_31),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_11),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_53),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_258),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_258),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_297),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_180),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_206),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_199),
.B(n_0),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_269),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_216),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_258),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_258),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_221),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_258),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_2),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_244),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_178),
.B(n_2),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_258),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_175),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_244),
.B(n_3),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_258),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_225),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_303),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_192),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_177),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_303),
.Y(n_369)
);

INVxp33_ASAP7_75t_SL g370 ( 
.A(n_175),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_226),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_177),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_214),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_303),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_228),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_303),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_214),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_303),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_283),
.B(n_3),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_182),
.B(n_5),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_283),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_241),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_189),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_182),
.B(n_189),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_229),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_303),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_230),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_232),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

BUFx6f_ASAP7_75t_SL g391 ( 
.A(n_201),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_233),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_238),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_194),
.B(n_7),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_238),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_237),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_194),
.B(n_8),
.Y(n_400)
);

INVxp33_ASAP7_75t_SL g401 ( 
.A(n_195),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_239),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_241),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_242),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_279),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_279),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_240),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_193),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_193),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_193),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_240),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_245),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_193),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_249),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_210),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_210),
.Y(n_420)
);

INVxp33_ASAP7_75t_SL g421 ( 
.A(n_195),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_210),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_318),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_210),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_246),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_187),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_187),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_260),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_261),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_262),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_275),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_383),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_368),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_345),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_366),
.A2(n_198),
.B(n_191),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_372),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_373),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_358),
.B(n_344),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_346),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_378),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_346),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_393),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_353),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_397),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_383),
.B(n_336),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_410),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_354),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_354),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_356),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_415),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_418),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_356),
.B(n_202),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_367),
.B(n_201),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_348),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_361),
.B(n_203),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_382),
.B(n_344),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_349),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_364),
.B(n_205),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_364),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_347),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_412),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_369),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_403),
.B(n_336),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_352),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_374),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_355),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_420),
.Y(n_477)
);

OA21x2_ASAP7_75t_L g478 ( 
.A1(n_374),
.A2(n_213),
.B(n_208),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_375),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_365),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_375),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_377),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_377),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_379),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_371),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_376),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_387),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_386),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_413),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_367),
.B(n_215),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_390),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_385),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_390),
.B(n_196),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_R g496 ( 
.A(n_388),
.B(n_313),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_429),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_429),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_389),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_392),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_399),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_402),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_426),
.B(n_173),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_461),
.B(n_405),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_434),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_446),
.Y(n_511)
);

BUFx4f_ASAP7_75t_L g512 ( 
.A(n_478),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_465),
.B(n_416),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_446),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_495),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_446),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_448),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_500),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_500),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_448),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_474),
.B(n_425),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_448),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_490),
.B(n_428),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_440),
.B(n_423),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_478),
.A2(n_350),
.B1(n_360),
.B2(n_357),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_437),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_490),
.B(n_432),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_478),
.A2(n_381),
.B1(n_401),
.B2(n_370),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_435),
.B(n_398),
.C(n_395),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

BUFx6f_ASAP7_75t_SL g531 ( 
.A(n_442),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_500),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_442),
.B(n_430),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_459),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_442),
.B(n_359),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_442),
.B(n_398),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_432),
.B(n_404),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_384),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_501),
.Y(n_539)
);

BUFx4f_ASAP7_75t_L g540 ( 
.A(n_478),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_452),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_452),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_471),
.B(n_404),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_496),
.A2(n_296),
.B1(n_311),
.B2(n_309),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_436),
.A2(n_463),
.B(n_458),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_459),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_471),
.B(n_406),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_500),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_503),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_495),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_440),
.A2(n_381),
.B1(n_421),
.B2(n_391),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_455),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_471),
.B(n_391),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_464),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_469),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_464),
.A2(n_380),
.B1(n_363),
.B2(n_311),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_469),
.A2(n_296),
.B1(n_309),
.B2(n_267),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_475),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_450),
.B(n_407),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_476),
.B(n_408),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_475),
.A2(n_256),
.B1(n_176),
.B2(n_212),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_475),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_435),
.B(n_406),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_443),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_443),
.B(n_409),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_444),
.B(n_409),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_458),
.A2(n_278),
.B1(n_316),
.B2(n_325),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_450),
.B(n_426),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_484),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_480),
.B(n_186),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_484),
.A2(n_497),
.B1(n_506),
.B2(n_493),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_493),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_444),
.B(n_427),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_493),
.A2(n_506),
.B1(n_497),
.B2(n_450),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_497),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_438),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_494),
.B(n_427),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_445),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_494),
.B(n_200),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_453),
.Y(n_586)
);

INVx6_ASAP7_75t_L g587 ( 
.A(n_450),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_441),
.A2(n_321),
.B1(n_291),
.B2(n_288),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_453),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_462),
.B(n_411),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_462),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_486),
.B(n_186),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_473),
.A2(n_247),
.B1(n_305),
.B2(n_271),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_467),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_487),
.B(n_489),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_467),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_473),
.A2(n_310),
.B1(n_320),
.B2(n_327),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_499),
.A2(n_321),
.B1(n_291),
.B2(n_288),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_473),
.B(n_441),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_472),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_472),
.B(n_411),
.Y(n_602)
);

OR2x6_ASAP7_75t_L g603 ( 
.A(n_505),
.B(n_396),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_479),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_495),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_473),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_481),
.Y(n_608)
);

BUFx4f_ASAP7_75t_L g609 ( 
.A(n_481),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_460),
.B(n_217),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_459),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_482),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_491),
.B(n_222),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_482),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_483),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_483),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_485),
.B(n_223),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_485),
.B(n_414),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_488),
.B(n_414),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_492),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_502),
.B(n_188),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_499),
.B(n_313),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_504),
.A2(n_400),
.B1(n_325),
.B2(n_343),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_459),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_507),
.B(n_188),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_463),
.A2(n_276),
.B1(n_252),
.B2(n_266),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_459),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_495),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_466),
.B(n_284),
.C(n_264),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_505),
.B(n_224),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_466),
.A2(n_314),
.B1(n_341),
.B2(n_285),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_468),
.B(n_190),
.Y(n_634)
);

OAI21xp33_ASAP7_75t_SL g635 ( 
.A1(n_436),
.A2(n_174),
.B(n_173),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_508),
.A2(n_319),
.B1(n_343),
.B2(n_339),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_508),
.A2(n_279),
.B1(n_215),
.B2(n_273),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_468),
.B(n_190),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_436),
.B(n_424),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_470),
.Y(n_640)
);

AND2x2_ASAP7_75t_SL g641 ( 
.A(n_470),
.B(n_196),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_495),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_470),
.B(n_424),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_495),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_470),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_470),
.B(n_417),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_495),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_470),
.B(n_417),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_433),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_477),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_477),
.B(n_419),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_477),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_512),
.A2(n_235),
.B(n_234),
.Y(n_655)
);

OAI21xp33_ASAP7_75t_L g656 ( 
.A1(n_632),
.A2(n_299),
.B(n_308),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_567),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_559),
.B(n_304),
.C(n_307),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_527),
.B(n_315),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_557),
.B(n_322),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_635),
.A2(n_281),
.B(n_243),
.C(n_236),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_557),
.B(n_331),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_524),
.B(n_197),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_523),
.B(n_277),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_524),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_510),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_526),
.B(n_439),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_587),
.B(n_280),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_567),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_518),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_528),
.B(n_197),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_587),
.B(n_607),
.Y(n_672)
);

AND2x6_ASAP7_75t_SL g673 ( 
.A(n_603),
.B(n_419),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_610),
.A2(n_174),
.B1(n_259),
.B2(n_323),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_538),
.B(n_259),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_609),
.A2(n_536),
.B(n_566),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_625),
.B(n_323),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_594),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_609),
.B(n_326),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_570),
.B(n_447),
.Y(n_680)
);

NAND2xp33_ASAP7_75t_L g681 ( 
.A(n_533),
.B(n_326),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_594),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_580),
.B(n_449),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_581),
.B(n_329),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_613),
.A2(n_329),
.B1(n_265),
.B2(n_254),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_556),
.B(n_607),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_596),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_625),
.B(n_287),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_530),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_518),
.B(n_293),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_584),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_530),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_525),
.A2(n_248),
.B1(n_251),
.B2(n_289),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_596),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_587),
.B(n_295),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_535),
.B(n_300),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_561),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_518),
.B(n_335),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_599),
.B(n_451),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_519),
.B(n_532),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_587),
.A2(n_294),
.B1(n_301),
.B2(n_302),
.Y(n_701)
);

AO221x1_ASAP7_75t_L g702 ( 
.A1(n_598),
.A2(n_196),
.B1(n_211),
.B2(n_255),
.C(n_340),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_599),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_561),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_554),
.B(n_456),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_574),
.B(n_317),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_624),
.B(n_457),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_561),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_560),
.B(n_215),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_585),
.B(n_334),
.C(n_333),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_606),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_592),
.B(n_324),
.Y(n_712)
);

NAND2x1_ASAP7_75t_L g713 ( 
.A(n_515),
.B(n_477),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_562),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_562),
.A2(n_257),
.B1(n_181),
.B2(n_183),
.Y(n_715)
);

AND2x6_ASAP7_75t_SL g716 ( 
.A(n_603),
.B(n_422),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_609),
.A2(n_179),
.B1(n_184),
.B2(n_185),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_606),
.A2(n_270),
.B1(n_218),
.B2(n_204),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_519),
.B(n_207),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_608),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_654),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_519),
.B(n_209),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_576),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_608),
.A2(n_274),
.B1(n_231),
.B2(n_219),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_515),
.B(n_553),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_532),
.B(n_196),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_532),
.B(n_220),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_603),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_623),
.B(n_273),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_612),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_551),
.B(n_227),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_612),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_551),
.B(n_512),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_509),
.B(n_273),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_635),
.A2(n_422),
.B(n_268),
.C(n_338),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_576),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_576),
.Y(n_737)
);

OAI22xp33_ASAP7_75t_L g738 ( 
.A1(n_546),
.A2(n_268),
.B1(n_338),
.B2(n_250),
.Y(n_738)
);

AND2x6_ASAP7_75t_SL g739 ( 
.A(n_603),
.B(n_9),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_627),
.B(n_16),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_551),
.B(n_16),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_614),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_603),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_572),
.B(n_290),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_572),
.B(n_292),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_614),
.Y(n_746)
);

AND2x6_ASAP7_75t_L g747 ( 
.A(n_639),
.B(n_340),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_634),
.B(n_17),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_616),
.B(n_286),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_582),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_534),
.Y(n_751)
);

BUFx6f_ASAP7_75t_SL g752 ( 
.A(n_650),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_L g753 ( 
.A(n_616),
.B(n_298),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_621),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_638),
.B(n_17),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_621),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_540),
.B(n_211),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_622),
.B(n_282),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_617),
.A2(n_312),
.B(n_253),
.C(n_337),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_582),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_513),
.B(n_521),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_622),
.B(n_578),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_552),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_641),
.A2(n_498),
.B1(n_340),
.B2(n_211),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_540),
.A2(n_639),
.B(n_511),
.C(n_544),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_582),
.B(n_272),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_537),
.B(n_19),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_L g768 ( 
.A(n_595),
.B(n_263),
.C(n_328),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_641),
.A2(n_498),
.B1(n_340),
.B2(n_255),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_540),
.B(n_255),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_586),
.A2(n_330),
.B1(n_255),
.B2(n_211),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_552),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_586),
.B(n_498),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_589),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_589),
.B(n_498),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_539),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_642),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_545),
.B(n_20),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_568),
.A2(n_498),
.B(n_74),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_591),
.B(n_20),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_591),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_600),
.B(n_604),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_600),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_604),
.B(n_22),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_550),
.B(n_24),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_539),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_563),
.B(n_636),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_643),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_641),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_546),
.B(n_34),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_615),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_615),
.B(n_620),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_620),
.B(n_34),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_588),
.B(n_38),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_577),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_541),
.Y(n_796)
);

INVx5_ASAP7_75t_L g797 ( 
.A(n_642),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_511),
.B(n_39),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_514),
.B(n_41),
.Y(n_799)
);

BUFx8_ASAP7_75t_L g800 ( 
.A(n_531),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_514),
.B(n_43),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_516),
.B(n_43),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_636),
.B(n_44),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_516),
.B(n_47),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_628),
.B(n_51),
.C(n_52),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_631),
.B(n_52),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_517),
.B(n_54),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_590),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_631),
.A2(n_547),
.B1(n_555),
.B2(n_579),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_643),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_571),
.A2(n_55),
.B1(n_56),
.B2(n_62),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_602),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_517),
.B(n_56),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_534),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_531),
.B(n_71),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_520),
.B(n_75),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_520),
.B(n_77),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_522),
.A2(n_85),
.B(n_89),
.C(n_103),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_522),
.B(n_167),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_691),
.B(n_588),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_676),
.A2(n_569),
.B(n_558),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_699),
.B(n_593),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_SL g823 ( 
.A1(n_733),
.A2(n_555),
.B(n_543),
.C(n_579),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_669),
.B(n_686),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_691),
.B(n_571),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_664),
.A2(n_633),
.B1(n_637),
.B2(n_547),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_810),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_664),
.B(n_597),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_733),
.A2(n_558),
.B(n_544),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_669),
.B(n_553),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_787),
.B(n_543),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_666),
.Y(n_832)
);

AOI22x1_ASAP7_75t_L g833 ( 
.A1(n_678),
.A2(n_541),
.B1(n_542),
.B2(n_548),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_700),
.A2(n_792),
.B(n_782),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_SL g835 ( 
.A(n_752),
.B(n_531),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_667),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_795),
.B(n_565),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_659),
.B(n_565),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_682),
.A2(n_529),
.B1(n_575),
.B2(n_573),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_721),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_687),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_763),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_665),
.B(n_703),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_703),
.B(n_564),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_672),
.A2(n_605),
.B1(n_515),
.B2(n_601),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_679),
.A2(n_583),
.B(n_651),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_SL g847 ( 
.A1(n_679),
.A2(n_618),
.B(n_619),
.C(n_645),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_765),
.A2(n_645),
.B(n_653),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_694),
.A2(n_583),
.B1(n_649),
.B2(n_651),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_808),
.B(n_651),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_719),
.A2(n_649),
.B(n_583),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_812),
.B(n_649),
.Y(n_852)
);

CKINVDCx10_ASAP7_75t_R g853 ( 
.A(n_752),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_663),
.B(n_653),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_722),
.A2(n_640),
.B(n_626),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_772),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_684),
.B(n_644),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_714),
.B(n_644),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_773),
.A2(n_652),
.B(n_648),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_775),
.A2(n_720),
.B(n_711),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_748),
.A2(n_601),
.B1(n_629),
.B2(n_611),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_680),
.B(n_601),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_730),
.A2(n_646),
.B(n_534),
.Y(n_863)
);

NOR2xp67_ASAP7_75t_L g864 ( 
.A(n_776),
.B(n_630),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_732),
.A2(n_654),
.B(n_534),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_728),
.B(n_654),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_683),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_721),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_707),
.B(n_654),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_689),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_743),
.B(n_654),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_790),
.A2(n_709),
.B1(n_738),
.B2(n_658),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_738),
.A2(n_642),
.B1(n_647),
.B2(n_629),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_742),
.A2(n_629),
.B(n_611),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_788),
.B(n_629),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_768),
.B(n_629),
.Y(n_876)
);

AOI21x1_ASAP7_75t_L g877 ( 
.A1(n_726),
.A2(n_611),
.B(n_549),
.Y(n_877)
);

AOI21x1_ASAP7_75t_L g878 ( 
.A1(n_726),
.A2(n_611),
.B(n_549),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_727),
.A2(n_611),
.B(n_549),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_721),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_794),
.A2(n_647),
.B1(n_642),
.B2(n_630),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_706),
.B(n_549),
.Y(n_882)
);

AOI21x1_ASAP7_75t_L g883 ( 
.A1(n_816),
.A2(n_534),
.B(n_647),
.Y(n_883)
);

NOR2x1p5_ASAP7_75t_SL g884 ( 
.A(n_697),
.B(n_630),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_712),
.B(n_630),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_746),
.A2(n_754),
.B1(n_756),
.B2(n_693),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_721),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_655),
.A2(n_630),
.B(n_112),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_755),
.A2(n_109),
.B1(n_121),
.B2(n_128),
.Y(n_889)
);

OAI21xp33_ASAP7_75t_L g890 ( 
.A1(n_656),
.A2(n_131),
.B(n_139),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_786),
.B(n_660),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_677),
.B(n_140),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_704),
.A2(n_142),
.B(n_143),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_755),
.A2(n_151),
.B1(n_152),
.B2(n_159),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_675),
.B(n_761),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_662),
.B(n_668),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_708),
.A2(n_750),
.B(n_736),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_803),
.Y(n_898)
);

O2A1O1Ixp5_ASAP7_75t_L g899 ( 
.A1(n_696),
.A2(n_785),
.B(n_778),
.C(n_767),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_668),
.B(n_695),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_695),
.B(n_657),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_819),
.A2(n_762),
.B(n_774),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_751),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_781),
.A2(n_791),
.B(n_767),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_731),
.A2(n_723),
.B(n_737),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_692),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_766),
.A2(n_758),
.B(n_749),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_690),
.A2(n_698),
.B(n_753),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_670),
.A2(n_760),
.B(n_681),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_670),
.A2(n_760),
.B(n_713),
.Y(n_910)
);

AOI21x1_ASAP7_75t_L g911 ( 
.A1(n_796),
.A2(n_799),
.B(n_802),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_729),
.B(n_745),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_673),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_729),
.B(n_705),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_688),
.B(n_744),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_783),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_674),
.B(n_740),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_740),
.B(n_685),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_780),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_817),
.A2(n_725),
.B(n_814),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_778),
.A2(n_785),
.B(n_817),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_715),
.B(n_734),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_725),
.A2(n_751),
.B(n_814),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_798),
.A2(n_813),
.B(n_807),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_800),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_735),
.A2(n_661),
.B(n_801),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_789),
.A2(n_741),
.B1(n_804),
.B2(n_769),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_671),
.B(n_789),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_741),
.B(n_793),
.Y(n_929)
);

AOI21x1_ASAP7_75t_L g930 ( 
.A1(n_784),
.A2(n_779),
.B(n_771),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_751),
.Y(n_931)
);

NOR2x1_ASAP7_75t_L g932 ( 
.A(n_805),
.B(n_710),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_751),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_806),
.A2(n_759),
.B(n_804),
.C(n_793),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_814),
.A2(n_818),
.B(n_764),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_777),
.B(n_797),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_701),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_814),
.A2(n_764),
.B(n_769),
.Y(n_938)
);

OAI21x1_ASAP7_75t_SL g939 ( 
.A1(n_811),
.A2(n_717),
.B(n_718),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_724),
.A2(n_815),
.B(n_777),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_777),
.A2(n_797),
.B(n_811),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_777),
.A2(n_797),
.B(n_702),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_747),
.B(n_800),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_797),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_739),
.A2(n_716),
.B(n_747),
.C(n_803),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_747),
.A2(n_803),
.B(n_748),
.C(n_755),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_747),
.B(n_699),
.Y(n_947)
);

AOI22x1_ASAP7_75t_L g948 ( 
.A1(n_747),
.A2(n_676),
.B1(n_589),
.B2(n_591),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_810),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_669),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_748),
.A2(n_755),
.B(n_740),
.C(n_655),
.Y(n_952)
);

CKINVDCx8_ASAP7_75t_R g953 ( 
.A(n_786),
.Y(n_953)
);

CKINVDCx8_ASAP7_75t_R g954 ( 
.A(n_786),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_955)
);

BUFx2_ASAP7_75t_SL g956 ( 
.A(n_752),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_678),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_678),
.A2(n_687),
.B1(n_694),
.B2(n_682),
.Y(n_958)
);

BUFx4f_ASAP7_75t_L g959 ( 
.A(n_667),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_748),
.A2(n_755),
.B(n_740),
.C(n_655),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_664),
.B(n_557),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_664),
.B(n_557),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_963)
);

OAI321xp33_ASAP7_75t_L g964 ( 
.A1(n_789),
.A2(n_811),
.A3(n_738),
.B1(n_588),
.B2(n_693),
.C(n_598),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_664),
.B(n_557),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_664),
.B(n_557),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_SL g968 ( 
.A(n_752),
.B(n_650),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_810),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_752),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_669),
.B(n_474),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_748),
.A2(n_755),
.B(n_740),
.C(n_655),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_L g975 ( 
.A1(n_709),
.A2(n_712),
.B(n_706),
.Y(n_975)
);

BUFx6f_ASAP7_75t_SL g976 ( 
.A(n_772),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_664),
.B(n_557),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_721),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_979)
);

AOI21x1_ASAP7_75t_L g980 ( 
.A1(n_757),
.A2(n_770),
.B(n_733),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_664),
.B(n_557),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_699),
.B(n_546),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_678),
.A2(n_687),
.B1(n_694),
.B2(n_682),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_664),
.B(n_557),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_752),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_664),
.B(n_557),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_721),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_699),
.B(n_546),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_721),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_691),
.B(n_368),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_676),
.A2(n_733),
.B(n_700),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_676),
.A2(n_809),
.B(n_765),
.Y(n_994)
);

OAI21x1_ASAP7_75t_SL g995 ( 
.A1(n_921),
.A2(n_939),
.B(n_926),
.Y(n_995)
);

OAI22x1_ASAP7_75t_L g996 ( 
.A1(n_820),
.A2(n_914),
.B1(n_825),
.B2(n_922),
.Y(n_996)
);

NAND2x1p5_ASAP7_75t_L g997 ( 
.A(n_903),
.B(n_951),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_896),
.B(n_912),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_953),
.Y(n_999)
);

INVx3_ASAP7_75t_SL g1000 ( 
.A(n_970),
.Y(n_1000)
);

AND2x6_ASAP7_75t_L g1001 ( 
.A(n_944),
.B(n_947),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_964),
.B(n_975),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_841),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_899),
.A2(n_960),
.B(n_952),
.Y(n_1004)
);

AOI221x1_ASAP7_75t_L g1005 ( 
.A1(n_973),
.A2(n_927),
.B1(n_900),
.B2(n_938),
.C(n_994),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_982),
.B(n_990),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_SL g1007 ( 
.A1(n_929),
.A2(n_917),
.B(n_901),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_907),
.A2(n_924),
.B(n_950),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_856),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_918),
.A2(n_828),
.B(n_946),
.C(n_934),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_822),
.B(n_867),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_961),
.B(n_962),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_903),
.B(n_951),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_950),
.A2(n_971),
.B(n_955),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_959),
.B(n_891),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_954),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_831),
.A2(n_826),
.B(n_892),
.C(n_928),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_985),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_965),
.B(n_967),
.Y(n_1019)
);

AOI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_992),
.A2(n_872),
.B(n_836),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_977),
.B(n_981),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_959),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_842),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_955),
.A2(n_974),
.B(n_971),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_827),
.B(n_949),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_984),
.B(n_986),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_924),
.A2(n_993),
.B(n_974),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_937),
.B(n_862),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_993),
.A2(n_966),
.B(n_963),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_979),
.A2(n_989),
.B(n_987),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_883),
.A2(n_821),
.B(n_948),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_843),
.B(n_844),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_832),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_869),
.B(n_895),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_886),
.A2(n_983),
.B1(n_958),
.B2(n_957),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_868),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_821),
.A2(n_848),
.B(n_829),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_920),
.A2(n_908),
.B(n_857),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_834),
.A2(n_847),
.B(n_865),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_865),
.A2(n_874),
.B(n_905),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_848),
.A2(n_902),
.B(n_879),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_976),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_913),
.B(n_969),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_956),
.B(n_925),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_874),
.A2(n_823),
.B(n_855),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_860),
.A2(n_863),
.B(n_897),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_840),
.B(n_880),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_976),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_916),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_863),
.A2(n_897),
.B(n_904),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_898),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_851),
.A2(n_935),
.B(n_824),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_980),
.A2(n_878),
.B(n_877),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_968),
.B(n_915),
.Y(n_1054)
);

CKINVDCx6p67_ASAP7_75t_R g1055 ( 
.A(n_853),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_935),
.A2(n_919),
.B(n_910),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_972),
.B(n_943),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_837),
.B(n_838),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_868),
.Y(n_1059)
);

AOI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_932),
.A2(n_858),
.B(n_854),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_923),
.A2(n_833),
.B(n_930),
.Y(n_1061)
);

OR2x6_ASAP7_75t_L g1062 ( 
.A(n_945),
.B(n_941),
.Y(n_1062)
);

OA22x2_ASAP7_75t_L g1063 ( 
.A1(n_850),
.A2(n_852),
.B1(n_889),
.B2(n_894),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_835),
.B(n_882),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_840),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_940),
.B(n_906),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_870),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_888),
.A2(n_938),
.A3(n_839),
.B(n_859),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_940),
.B(n_880),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_875),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_864),
.B(n_991),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_888),
.A2(n_890),
.B(n_941),
.C(n_893),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_859),
.A2(n_846),
.B(n_942),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_942),
.A2(n_849),
.A3(n_893),
.B(n_909),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_936),
.A2(n_944),
.B(n_876),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_868),
.B(n_991),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_936),
.A2(n_871),
.B(n_866),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_887),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_861),
.A2(n_830),
.B(n_885),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_887),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_931),
.B(n_933),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_931),
.A2(n_933),
.B(n_988),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_933),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_884),
.A2(n_845),
.B(n_873),
.C(n_881),
.Y(n_1084)
);

BUFx10_ASAP7_75t_L g1085 ( 
.A(n_978),
.Y(n_1085)
);

CKINVDCx8_ASAP7_75t_R g1086 ( 
.A(n_978),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_978),
.B(n_988),
.Y(n_1087)
);

AO31x2_ASAP7_75t_L g1088 ( 
.A1(n_988),
.A2(n_927),
.A3(n_924),
.B(n_765),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_921),
.A2(n_960),
.B(n_973),
.C(n_952),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_912),
.B(n_964),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_921),
.A2(n_960),
.B(n_973),
.C(n_952),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_902),
.A2(n_911),
.B(n_924),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_959),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_832),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_921),
.A2(n_899),
.B(n_952),
.Y(n_1095)
);

O2A1O1Ixp5_ASAP7_75t_L g1096 ( 
.A1(n_921),
.A2(n_927),
.B(n_899),
.C(n_929),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_921),
.A2(n_960),
.B(n_973),
.C(n_952),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_921),
.A2(n_899),
.B(n_952),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_921),
.A2(n_929),
.B(n_900),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_950),
.A2(n_971),
.B(n_955),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_896),
.B(n_665),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_896),
.B(n_665),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_921),
.A2(n_899),
.B(n_952),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_950),
.A2(n_971),
.B(n_955),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_896),
.B(n_665),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_982),
.B(n_990),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_950),
.A2(n_971),
.B(n_955),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_856),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_950),
.A2(n_971),
.B(n_955),
.Y(n_1109)
);

AOI31xp33_ASAP7_75t_L g1110 ( 
.A1(n_872),
.A2(n_546),
.A3(n_560),
.B(n_588),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_896),
.B(n_665),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_953),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_982),
.B(n_990),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_902),
.A2(n_911),
.B(n_924),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_959),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_950),
.A2(n_971),
.B(n_955),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_841),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_921),
.A2(n_899),
.B(n_952),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_868),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_976),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_902),
.A2(n_911),
.B(n_924),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_952),
.A2(n_973),
.B(n_960),
.C(n_921),
.Y(n_1122)
);

O2A1O1Ixp5_ASAP7_75t_L g1123 ( 
.A1(n_921),
.A2(n_927),
.B(n_899),
.C(n_929),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_921),
.A2(n_929),
.B(n_900),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_921),
.A2(n_929),
.B(n_900),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_953),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_921),
.A2(n_899),
.B(n_952),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_832),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_896),
.B(n_665),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_896),
.B(n_665),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_950),
.A2(n_971),
.B(n_955),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_917),
.A2(n_918),
.B(n_975),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_953),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_842),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_976),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_950),
.A2(n_971),
.B(n_955),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_921),
.A2(n_929),
.B(n_927),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1086),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_1135),
.Y(n_1139)
);

INVxp67_ASAP7_75t_SL g1140 ( 
.A(n_1028),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1003),
.Y(n_1141)
);

NOR2xp67_ASAP7_75t_L g1142 ( 
.A(n_1022),
.B(n_1093),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_998),
.B(n_1015),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_SL g1144 ( 
.A1(n_996),
.A2(n_1002),
.B1(n_1090),
.B2(n_1113),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1006),
.B(n_1106),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1089),
.A2(n_1091),
.B(n_1097),
.C(n_1122),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1090),
.A2(n_1002),
.B1(n_1011),
.B2(n_1054),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1034),
.B(n_1134),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1035),
.A2(n_1122),
.B1(n_1124),
.B2(n_1125),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1124),
.A2(n_1125),
.B(n_1072),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_999),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1023),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_SL g1153 ( 
.A(n_1017),
.B(n_1042),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1132),
.B(n_1012),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1115),
.B(n_1119),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_999),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1019),
.B(n_1021),
.Y(n_1157)
);

CKINVDCx11_ASAP7_75t_R g1158 ( 
.A(n_1055),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1119),
.B(n_1087),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1026),
.B(n_1058),
.Y(n_1160)
);

AO32x1_ASAP7_75t_L g1161 ( 
.A1(n_1005),
.A2(n_1137),
.A3(n_1070),
.B1(n_1004),
.B2(n_1049),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1119),
.B(n_1087),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1120),
.B(n_1133),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_1009),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1120),
.B(n_1133),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1043),
.B(n_1009),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1095),
.A2(n_1098),
.B1(n_1118),
.B2(n_1103),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1038),
.A2(n_1127),
.B(n_1008),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1094),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1096),
.A2(n_1123),
.B(n_1030),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1036),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1112),
.A2(n_1000),
.B1(n_1044),
.B2(n_1062),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1030),
.A2(n_1029),
.B(n_995),
.Y(n_1173)
);

O2A1O1Ixp5_ASAP7_75t_SL g1174 ( 
.A1(n_1020),
.A2(n_1046),
.B(n_1060),
.C(n_1050),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_1052),
.A2(n_1010),
.B(n_1056),
.C(n_1027),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1101),
.B(n_1102),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1032),
.B(n_1001),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1135),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1117),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1001),
.B(n_1062),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1108),
.B(n_1051),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1056),
.A2(n_1039),
.B(n_1063),
.Y(n_1182)
);

INVx3_ASAP7_75t_SL g1183 ( 
.A(n_1112),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1108),
.B(n_1105),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1044),
.B(n_1001),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1110),
.A2(n_1063),
.B1(n_1062),
.B2(n_1129),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_1092),
.A2(n_1121),
.B(n_1114),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1016),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1111),
.B(n_1130),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1126),
.Y(n_1190)
);

AOI221x1_ASAP7_75t_L g1191 ( 
.A1(n_1052),
.A2(n_1039),
.B1(n_1069),
.B2(n_1040),
.C(n_1066),
.Y(n_1191)
);

O2A1O1Ixp5_ASAP7_75t_SL g1192 ( 
.A1(n_1064),
.A2(n_1083),
.B(n_1059),
.C(n_1067),
.Y(n_1192)
);

BUFx12f_ASAP7_75t_L g1193 ( 
.A(n_1018),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1040),
.A2(n_1045),
.B(n_1131),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1001),
.B(n_1128),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1025),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1045),
.A2(n_1136),
.B(n_1116),
.Y(n_1197)
);

AOI21x1_ASAP7_75t_SL g1198 ( 
.A1(n_1007),
.A2(n_1071),
.B(n_1081),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1044),
.B(n_1001),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1048),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1025),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1048),
.B(n_1065),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1037),
.A2(n_1109),
.B(n_1107),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1078),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1000),
.B(n_1057),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1076),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1036),
.B(n_1080),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1036),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1085),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1085),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1059),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1083),
.Y(n_1212)
);

OAI21xp33_ASAP7_75t_L g1213 ( 
.A1(n_997),
.A2(n_1013),
.B(n_1047),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1084),
.A2(n_1047),
.B1(n_1082),
.B2(n_1088),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1077),
.A2(n_1082),
.B1(n_1079),
.B2(n_1075),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1014),
.A2(n_1104),
.B(n_1024),
.Y(n_1216)
);

BUFx12f_ASAP7_75t_L g1217 ( 
.A(n_1074),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1068),
.B(n_1073),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1100),
.A2(n_1031),
.B(n_1061),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1041),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1068),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1009),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1089),
.A2(n_1097),
.B1(n_1091),
.B2(n_921),
.Y(n_1223)
);

OAI21xp33_ASAP7_75t_L g1224 ( 
.A1(n_1089),
.A2(n_960),
.B(n_952),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1099),
.A2(n_921),
.B(n_929),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1006),
.B(n_1106),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1023),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1003),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1099),
.A2(n_921),
.B(n_929),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1055),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1086),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1086),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1009),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1003),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1009),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1003),
.Y(n_1237)
);

CKINVDCx8_ASAP7_75t_R g1238 ( 
.A(n_1134),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1055),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1002),
.A2(n_546),
.B1(n_709),
.B2(n_820),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1086),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1006),
.B(n_1106),
.Y(n_1243)
);

BUFx12f_ASAP7_75t_L g1244 ( 
.A(n_1135),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1089),
.A2(n_1097),
.B1(n_1091),
.B2(n_921),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1099),
.A2(n_921),
.B(n_929),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1002),
.A2(n_546),
.B1(n_709),
.B2(n_820),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1090),
.B(n_815),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1061),
.A2(n_1031),
.B(n_1053),
.Y(n_1249)
);

INVx5_ASAP7_75t_L g1250 ( 
.A(n_1001),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1006),
.B(n_1106),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1006),
.B(n_1106),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1033),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1089),
.A2(n_1097),
.B1(n_1091),
.B2(n_921),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1135),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1135),
.Y(n_1257)
);

CKINVDCx6p67_ASAP7_75t_R g1258 ( 
.A(n_1055),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1009),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1006),
.B(n_1106),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1055),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1099),
.A2(n_921),
.B(n_929),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1090),
.B(n_1028),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1009),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1006),
.B(n_1106),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1135),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1185),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1218),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1183),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1140),
.B(n_1226),
.Y(n_1275)
);

AO21x1_ASAP7_75t_L g1276 ( 
.A1(n_1186),
.A2(n_1248),
.B(n_1167),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1248),
.A2(n_1144),
.B1(n_1186),
.B2(n_1153),
.Y(n_1277)
);

CKINVDCx6p67_ASAP7_75t_R g1278 ( 
.A(n_1158),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1240),
.A2(n_1247),
.B1(n_1254),
.B2(n_1241),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1218),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1226),
.A2(n_1260),
.B1(n_1263),
.B2(n_1264),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1222),
.Y(n_1282)
);

NAND2x1_ASAP7_75t_L g1283 ( 
.A(n_1215),
.B(n_1149),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1219),
.A2(n_1249),
.B(n_1197),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_R g1285 ( 
.A1(n_1148),
.A2(n_1176),
.B1(n_1262),
.B2(n_1251),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1153),
.A2(n_1263),
.B1(n_1261),
.B2(n_1265),
.Y(n_1286)
);

BUFx2_ASAP7_75t_R g1287 ( 
.A(n_1231),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1241),
.A2(n_1264),
.B1(n_1261),
.B2(n_1260),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1238),
.B(n_1151),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1254),
.A2(n_1268),
.B1(n_1265),
.B2(n_1243),
.Y(n_1290)
);

BUFx12f_ASAP7_75t_L g1291 ( 
.A(n_1239),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1268),
.A2(n_1143),
.B1(n_1147),
.B2(n_1145),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1179),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1250),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1227),
.A2(n_1270),
.B1(n_1252),
.B2(n_1154),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1185),
.B(n_1199),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1199),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1223),
.A2(n_1255),
.B1(n_1245),
.B2(n_1154),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1170),
.A2(n_1194),
.B(n_1168),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1223),
.A2(n_1245),
.B1(n_1255),
.B2(n_1224),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1229),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1266),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1167),
.A2(n_1267),
.B(n_1225),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1235),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1196),
.A2(n_1201),
.B1(n_1253),
.B2(n_1169),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1173),
.A2(n_1175),
.B(n_1216),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1187),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1237),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1146),
.A2(n_1164),
.B1(n_1149),
.B2(n_1234),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1191),
.A2(n_1150),
.B(n_1216),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1177),
.A2(n_1217),
.B1(n_1166),
.B2(n_1189),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1171),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1184),
.B(n_1180),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1180),
.B(n_1206),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1177),
.A2(n_1160),
.B1(n_1157),
.B2(n_1221),
.Y(n_1315)
);

BUFx10_ASAP7_75t_L g1316 ( 
.A(n_1163),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1204),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1236),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1259),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1160),
.A2(n_1195),
.B1(n_1172),
.B2(n_1214),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1138),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1214),
.A2(n_1138),
.B1(n_1205),
.B2(n_1232),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1159),
.B(n_1162),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1195),
.A2(n_1181),
.B1(n_1156),
.B2(n_1269),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1161),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1138),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1161),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1208),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1171),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1258),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1203),
.A2(n_1182),
.B(n_1267),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1202),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1202),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1161),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1188),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1232),
.A2(n_1233),
.B1(n_1242),
.B2(n_1190),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1225),
.A2(n_1246),
.B(n_1230),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1220),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1233),
.A2(n_1242),
.B1(n_1200),
.B2(n_1152),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1228),
.B(n_1211),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1174),
.A2(n_1192),
.B(n_1213),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1207),
.A2(n_1198),
.B(n_1142),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1212),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1155),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1155),
.A2(n_1139),
.B(n_1178),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1209),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1209),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1209),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1210),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1210),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1163),
.A2(n_1165),
.B1(n_1244),
.B2(n_1256),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1271),
.A2(n_1210),
.B(n_1257),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1193),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_1165),
.Y(n_1354)
);

INVxp33_ASAP7_75t_L g1355 ( 
.A(n_1271),
.Y(n_1355)
);

BUFx8_ASAP7_75t_SL g1356 ( 
.A(n_1231),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1141),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1240),
.A2(n_1002),
.B1(n_1247),
.B2(n_709),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1141),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1141),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1218),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1158),
.Y(n_1362)
);

CKINVDCx11_ASAP7_75t_R g1363 ( 
.A(n_1158),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1158),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1138),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1141),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1145),
.B(n_1227),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1222),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_1158),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1240),
.A2(n_1002),
.B1(n_1247),
.B2(n_709),
.Y(n_1370)
);

CKINVDCx11_ASAP7_75t_R g1371 ( 
.A(n_1158),
.Y(n_1371)
);

CKINVDCx11_ASAP7_75t_R g1372 ( 
.A(n_1158),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1140),
.B(n_1226),
.Y(n_1373)
);

AO21x1_ASAP7_75t_L g1374 ( 
.A1(n_1186),
.A2(n_921),
.B(n_1248),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1141),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_1164),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1248),
.A2(n_372),
.B1(n_373),
.B2(n_368),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1141),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1141),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1273),
.B(n_1280),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1376),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1314),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1313),
.B(n_1273),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1280),
.B(n_1361),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1282),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1338),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1281),
.B(n_1288),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1345),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1293),
.B(n_1301),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1304),
.B(n_1308),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1275),
.B(n_1373),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1284),
.A2(n_1306),
.B(n_1337),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1283),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1283),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1356),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1368),
.B(n_1318),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1290),
.B(n_1298),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1360),
.B(n_1366),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1319),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1309),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1306),
.A2(n_1303),
.B(n_1341),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1379),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1345),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1378),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1375),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1328),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1299),
.A2(n_1307),
.B(n_1374),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1310),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1300),
.B(n_1292),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1316),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1325),
.A2(n_1334),
.B(n_1327),
.Y(n_1412)
);

OA21x2_ASAP7_75t_L g1413 ( 
.A1(n_1325),
.A2(n_1334),
.B(n_1327),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1331),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1367),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1316),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1335),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1354),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1374),
.A2(n_1276),
.B(n_1317),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1367),
.B(n_1295),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1344),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1276),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1342),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1320),
.A2(n_1315),
.B(n_1279),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1311),
.B(n_1333),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1342),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1342),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1332),
.B(n_1324),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1286),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1294),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1294),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1344),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1343),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1329),
.Y(n_1434)
);

INVxp67_ASAP7_75t_L g1435 ( 
.A(n_1340),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1364),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1358),
.A2(n_1370),
.B(n_1305),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1418),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1414),
.B(n_1277),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1401),
.B(n_1339),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1412),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1409),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1412),
.B(n_1322),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1393),
.B(n_1336),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1412),
.B(n_1274),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1391),
.B(n_1348),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1409),
.B(n_1312),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1398),
.B(n_1346),
.Y(n_1448)
);

AOI33xp33_ASAP7_75t_L g1449 ( 
.A1(n_1422),
.A2(n_1377),
.A3(n_1285),
.B1(n_1351),
.B2(n_1350),
.B3(n_1347),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1391),
.B(n_1348),
.Y(n_1450)
);

AOI31xp33_ASAP7_75t_L g1451 ( 
.A1(n_1410),
.A2(n_1296),
.A3(n_1272),
.B(n_1355),
.Y(n_1451)
);

INVxp67_ASAP7_75t_SL g1452 ( 
.A(n_1381),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1383),
.B(n_1297),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1386),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1407),
.Y(n_1455)
);

OAI31xp33_ASAP7_75t_L g1456 ( 
.A1(n_1410),
.A2(n_1285),
.A3(n_1326),
.B(n_1321),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1386),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1422),
.B(n_1352),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1387),
.A2(n_1278),
.B1(n_1335),
.B2(n_1364),
.Y(n_1459)
);

NAND2xp33_ASAP7_75t_R g1460 ( 
.A(n_1380),
.B(n_1353),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1413),
.B(n_1382),
.Y(n_1461)
);

BUFx12f_ASAP7_75t_L g1462 ( 
.A(n_1395),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1424),
.A2(n_1369),
.B1(n_1362),
.B2(n_1323),
.Y(n_1463)
);

AND2x2_ASAP7_75t_SL g1464 ( 
.A(n_1380),
.B(n_1323),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1393),
.B(n_1289),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_1440),
.B(n_1433),
.C(n_1400),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1439),
.A2(n_1437),
.B1(n_1429),
.B2(n_1424),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1464),
.B(n_1393),
.Y(n_1468)
);

OAI211xp5_ASAP7_75t_L g1469 ( 
.A1(n_1440),
.A2(n_1456),
.B(n_1455),
.C(n_1444),
.Y(n_1469)
);

NAND3xp33_ASAP7_75t_L g1470 ( 
.A(n_1445),
.B(n_1426),
.C(n_1427),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1459),
.A2(n_1429),
.B1(n_1424),
.B2(n_1394),
.Y(n_1471)
);

NAND4xp25_ASAP7_75t_L g1472 ( 
.A(n_1459),
.B(n_1396),
.C(n_1435),
.D(n_1417),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1452),
.B(n_1385),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1439),
.A2(n_1419),
.B1(n_1420),
.B2(n_1405),
.C(n_1403),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1452),
.B(n_1396),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1461),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1449),
.A2(n_1415),
.B1(n_1420),
.B2(n_1384),
.C(n_1394),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1455),
.B(n_1389),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1446),
.B(n_1450),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1446),
.B(n_1389),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1453),
.B(n_1394),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1439),
.A2(n_1437),
.B1(n_1424),
.B2(n_1425),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1456),
.A2(n_1384),
.B(n_1355),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1463),
.A2(n_1437),
.B1(n_1432),
.B2(n_1421),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_SL g1485 ( 
.A(n_1460),
.B(n_1353),
.C(n_1302),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1464),
.A2(n_1437),
.B1(n_1421),
.B2(n_1436),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1464),
.B(n_1451),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1454),
.B(n_1390),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1442),
.A2(n_1392),
.B(n_1423),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1444),
.A2(n_1428),
.B(n_1430),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1445),
.B(n_1458),
.C(n_1448),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1443),
.A2(n_1411),
.B1(n_1416),
.B2(n_1278),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1454),
.B(n_1397),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1457),
.B(n_1397),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1457),
.B(n_1399),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1462),
.B(n_1362),
.Y(n_1496)
);

XNOR2x1_ASAP7_75t_SL g1497 ( 
.A(n_1460),
.B(n_1428),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1445),
.B(n_1426),
.C(n_1427),
.Y(n_1498)
);

NOR3xp33_ASAP7_75t_L g1499 ( 
.A(n_1458),
.B(n_1408),
.C(n_1434),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1453),
.B(n_1388),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1443),
.A2(n_1431),
.B1(n_1430),
.B2(n_1349),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1449),
.B(n_1402),
.C(n_1406),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1443),
.A2(n_1419),
.B1(n_1404),
.B2(n_1425),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1476),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1489),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1472),
.B(n_1465),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1489),
.Y(n_1507)
);

INVx4_ASAP7_75t_L g1508 ( 
.A(n_1489),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1479),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1500),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1481),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1475),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1478),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1488),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1493),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1491),
.B(n_1441),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1494),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1470),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1498),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_1461),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1480),
.B(n_1441),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1466),
.B(n_1465),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1495),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1468),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1468),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1502),
.B(n_1461),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1499),
.B(n_1447),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1501),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1447),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1528),
.B(n_1497),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1504),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1504),
.Y(n_1532)
);

AND2x4_ASAP7_75t_SL g1533 ( 
.A(n_1529),
.B(n_1465),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1509),
.B(n_1490),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1520),
.B(n_1438),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1504),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1526),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1514),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1505),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1505),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1505),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1505),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1514),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1514),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1512),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1509),
.B(n_1469),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1515),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1515),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1515),
.Y(n_1549)
);

OAI21xp33_ASAP7_75t_L g1550 ( 
.A1(n_1526),
.A2(n_1477),
.B(n_1471),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1517),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1507),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1512),
.Y(n_1553)
);

AO21x1_ASAP7_75t_L g1554 ( 
.A1(n_1508),
.A2(n_1486),
.B(n_1487),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1517),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1517),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1520),
.B(n_1438),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1523),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1509),
.B(n_1474),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1512),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1526),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1520),
.B(n_1438),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1507),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1523),
.Y(n_1564)
);

NAND2x1p5_ASAP7_75t_L g1565 ( 
.A(n_1525),
.B(n_1487),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1518),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1523),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1513),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1513),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1566),
.B(n_1518),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1531),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1530),
.B(n_1528),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1566),
.B(n_1506),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1566),
.B(n_1546),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1531),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1537),
.B(n_1518),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1561),
.B(n_1516),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1550),
.B(n_1518),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1530),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1532),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1516),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1539),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1532),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1536),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1533),
.B(n_1528),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1533),
.B(n_1511),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1506),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1565),
.Y(n_1589)
);

NOR2xp67_ASAP7_75t_SL g1590 ( 
.A(n_1559),
.B(n_1369),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1536),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1565),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1553),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1560),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1539),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1568),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1533),
.B(n_1529),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1568),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1535),
.B(n_1519),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1569),
.B(n_1519),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1569),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1538),
.B(n_1519),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1538),
.B(n_1529),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1543),
.B(n_1519),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1565),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1554),
.B(n_1511),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1554),
.B(n_1511),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1543),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1544),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1544),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1547),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1547),
.B(n_1363),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1572),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1606),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1579),
.A2(n_1503),
.B1(n_1508),
.B2(n_1507),
.C(n_1482),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1606),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1576),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1588),
.A2(n_1574),
.B1(n_1607),
.B2(n_1575),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1607),
.B(n_1527),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1597),
.B(n_1508),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1597),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1603),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1573),
.B(n_1548),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1612),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1573),
.B(n_1548),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1603),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1586),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1586),
.B(n_1527),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1588),
.B(n_1549),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1508),
.Y(n_1630)
);

AND2x4_ASAP7_75t_SL g1631 ( 
.A(n_1587),
.B(n_1485),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1580),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1581),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1584),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1578),
.B(n_1577),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1610),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1585),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1570),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1591),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1610),
.B(n_1549),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1596),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1587),
.B(n_1527),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1574),
.A2(n_1522),
.B1(n_1525),
.B2(n_1529),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1598),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1590),
.B(n_1363),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1601),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1578),
.B(n_1551),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1612),
.A2(n_1467),
.B1(n_1484),
.B2(n_1508),
.Y(n_1648)
);

NOR2xp67_ASAP7_75t_L g1649 ( 
.A(n_1621),
.B(n_1599),
.Y(n_1649)
);

AOI31xp33_ASAP7_75t_L g1650 ( 
.A1(n_1618),
.A2(n_1496),
.A3(n_1599),
.B(n_1302),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1615),
.A2(n_1600),
.B(n_1604),
.C(n_1602),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1613),
.Y(n_1652)
);

NAND2x1_ASAP7_75t_L g1653 ( 
.A(n_1621),
.B(n_1603),
.Y(n_1653)
);

O2A1O1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1614),
.A2(n_1605),
.B(n_1592),
.C(n_1589),
.Y(n_1654)
);

A2O1A1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1648),
.A2(n_1571),
.B(n_1507),
.C(n_1582),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1632),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1614),
.A2(n_1508),
.B1(n_1542),
.B2(n_1541),
.C(n_1563),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1613),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

NOR4xp25_ASAP7_75t_L g1660 ( 
.A(n_1616),
.B(n_1593),
.C(n_1594),
.D(n_1582),
.Y(n_1660)
);

NAND2x1p5_ASAP7_75t_L g1661 ( 
.A(n_1645),
.B(n_1321),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1627),
.B(n_1326),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1617),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1636),
.B(n_1527),
.Y(n_1664)
);

AOI21xp33_ASAP7_75t_L g1665 ( 
.A1(n_1638),
.A2(n_1616),
.B(n_1629),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_SL g1666 ( 
.A1(n_1635),
.A2(n_1583),
.B1(n_1595),
.B2(n_1552),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1633),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1638),
.B(n_1551),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1633),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1634),
.Y(n_1670)
);

OAI21xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1619),
.A2(n_1609),
.B(n_1608),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1631),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1622),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1640),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1672),
.B(n_1622),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1662),
.B(n_1624),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1656),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1652),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1672),
.B(n_1371),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1660),
.B(n_1619),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1658),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1649),
.B(n_1626),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1660),
.B(n_1626),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1664),
.B(n_1674),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1659),
.B(n_1663),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1673),
.B(n_1623),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1653),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1661),
.B(n_1631),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1650),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1661),
.B(n_1628),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1665),
.B(n_1628),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1667),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1671),
.B(n_1642),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1669),
.B(n_1642),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1680),
.A2(n_1655),
.B1(n_1650),
.B2(n_1651),
.Y(n_1695)
);

AOI222xp33_ASAP7_75t_L g1696 ( 
.A1(n_1683),
.A2(n_1657),
.B1(n_1670),
.B2(n_1668),
.C1(n_1643),
.C2(n_1666),
.Y(n_1696)
);

NOR3x1_ASAP7_75t_L g1697 ( 
.A(n_1684),
.B(n_1635),
.C(n_1625),
.Y(n_1697)
);

AOI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1683),
.A2(n_1654),
.B(n_1630),
.C(n_1620),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1679),
.B(n_1620),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1691),
.A2(n_1634),
.B1(n_1637),
.B2(n_1646),
.C(n_1644),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1676),
.A2(n_1693),
.B(n_1689),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1693),
.A2(n_1662),
.B(n_1639),
.Y(n_1702)
);

OAI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1691),
.A2(n_1647),
.B(n_1639),
.Y(n_1703)
);

AOI21xp33_ASAP7_75t_SL g1704 ( 
.A1(n_1687),
.A2(n_1647),
.B(n_1630),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1682),
.A2(n_1595),
.B1(n_1583),
.B2(n_1620),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1681),
.A2(n_1552),
.B(n_1542),
.C(n_1541),
.Y(n_1706)
);

AOI211x1_ASAP7_75t_L g1707 ( 
.A1(n_1701),
.A2(n_1677),
.B(n_1675),
.C(n_1682),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1703),
.B(n_1675),
.Y(n_1708)
);

AND3x1_ASAP7_75t_L g1709 ( 
.A(n_1698),
.B(n_1688),
.C(n_1677),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1699),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1697),
.B(n_1690),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1695),
.B(n_1686),
.C(n_1685),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1704),
.B(n_1688),
.Y(n_1713)
);

NOR3xp33_ASAP7_75t_L g1714 ( 
.A(n_1702),
.B(n_1700),
.C(n_1685),
.Y(n_1714)
);

NAND2x1p5_ASAP7_75t_L g1715 ( 
.A(n_1705),
.B(n_1371),
.Y(n_1715)
);

NAND5xp2_ASAP7_75t_L g1716 ( 
.A(n_1696),
.B(n_1690),
.C(n_1694),
.D(n_1692),
.E(n_1678),
.Y(n_1716)
);

NAND3xp33_ASAP7_75t_SL g1717 ( 
.A(n_1706),
.B(n_1681),
.C(n_1694),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1711),
.B(n_1681),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1716),
.B(n_1678),
.Y(n_1719)
);

AOI311xp33_ASAP7_75t_L g1720 ( 
.A1(n_1714),
.A2(n_1692),
.A3(n_1646),
.B(n_1644),
.C(n_1641),
.Y(n_1720)
);

NOR3xp33_ASAP7_75t_L g1721 ( 
.A(n_1712),
.B(n_1372),
.C(n_1330),
.Y(n_1721)
);

NOR4xp25_ASAP7_75t_L g1722 ( 
.A(n_1717),
.B(n_1641),
.C(n_1637),
.D(n_1611),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_L g1723 ( 
.A(n_1713),
.B(n_1372),
.C(n_1330),
.Y(n_1723)
);

OAI211xp5_ASAP7_75t_SL g1724 ( 
.A1(n_1710),
.A2(n_1287),
.B(n_1562),
.C(n_1557),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1723),
.B(n_1709),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1719),
.A2(n_1708),
.B1(n_1715),
.B2(n_1630),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1718),
.A2(n_1721),
.B1(n_1724),
.B2(n_1722),
.Y(n_1727)
);

AO22x1_ASAP7_75t_L g1728 ( 
.A1(n_1720),
.A2(n_1707),
.B1(n_1356),
.B2(n_1291),
.Y(n_1728)
);

OAI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1719),
.A2(n_1563),
.B1(n_1540),
.B2(n_1291),
.Y(n_1729)
);

INVxp67_ASAP7_75t_SL g1730 ( 
.A(n_1719),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1718),
.Y(n_1731)
);

NAND2x1p5_ASAP7_75t_SL g1732 ( 
.A(n_1719),
.B(n_1525),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1731),
.B(n_1620),
.Y(n_1733)
);

NOR3xp33_ASAP7_75t_L g1734 ( 
.A(n_1730),
.B(n_1630),
.C(n_1540),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1725),
.B(n_1462),
.Y(n_1735)
);

NOR4xp25_ASAP7_75t_L g1736 ( 
.A(n_1729),
.B(n_1567),
.C(n_1564),
.D(n_1555),
.Y(n_1736)
);

NAND3x1_ASAP7_75t_L g1737 ( 
.A(n_1726),
.B(n_1462),
.C(n_1555),
.Y(n_1737)
);

NOR2x1_ASAP7_75t_L g1738 ( 
.A(n_1732),
.B(n_1535),
.Y(n_1738)
);

XNOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1735),
.B(n_1727),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1738),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1733),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1740),
.A2(n_1734),
.B1(n_1737),
.B2(n_1728),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1742),
.B(n_1741),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1743),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1743),
.B(n_1739),
.Y(n_1745)
);

AOI31xp33_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1736),
.A3(n_1525),
.B(n_1524),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1744),
.B(n_1556),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1567),
.B1(n_1564),
.B2(n_1556),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1746),
.A2(n_1558),
.B(n_1521),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1558),
.B(n_1521),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1748),
.B1(n_1365),
.B2(n_1492),
.Y(n_1751)
);

OAI221xp5_ASAP7_75t_R g1752 ( 
.A1(n_1751),
.A2(n_1562),
.B1(n_1557),
.B2(n_1510),
.C(n_1497),
.Y(n_1752)
);

AOI211xp5_ASAP7_75t_L g1753 ( 
.A1(n_1752),
.A2(n_1522),
.B(n_1483),
.C(n_1524),
.Y(n_1753)
);


endmodule