module real_aes_633_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_316;
wire n_284;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g530 ( .A(n_0), .B(n_141), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_1), .B(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_2), .B(n_123), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_3), .B(n_139), .Y(n_158) );
INVx1_ASAP7_75t_L g130 ( .A(n_4), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_5), .B(n_123), .Y(n_461) );
NAND2xp33_ASAP7_75t_SL g515 ( .A(n_6), .B(n_129), .Y(n_515) );
INVx1_ASAP7_75t_L g508 ( .A(n_7), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g761 ( .A(n_8), .Y(n_761) );
AND2x2_ASAP7_75t_L g459 ( .A(n_9), .B(n_144), .Y(n_459) );
AND2x2_ASAP7_75t_L g160 ( .A(n_10), .B(n_148), .Y(n_160) );
AND2x2_ASAP7_75t_L g169 ( .A(n_11), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g145 ( .A(n_12), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_13), .B(n_139), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_14), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g759 ( .A(n_14), .B(n_760), .C(n_762), .Y(n_759) );
AOI221x1_ASAP7_75t_L g511 ( .A1(n_15), .A2(n_132), .B1(n_170), .B2(n_512), .C(n_514), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_16), .B(n_123), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_17), .B(n_123), .Y(n_203) );
INVx1_ASAP7_75t_L g447 ( .A(n_18), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_19), .A2(n_92), .B1(n_123), .B2(n_233), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_20), .A2(n_73), .B1(n_746), .B2(n_747), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_20), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_21), .A2(n_132), .B(n_463), .Y(n_462) );
AOI221xp5_ASAP7_75t_SL g520 ( .A1(n_22), .A2(n_37), .B1(n_123), .B2(n_132), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_23), .B(n_141), .Y(n_464) );
OR2x2_ASAP7_75t_L g146 ( .A(n_24), .B(n_91), .Y(n_146) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_24), .A2(n_91), .B(n_145), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_25), .B(n_139), .Y(n_502) );
INVxp67_ASAP7_75t_L g510 ( .A(n_26), .Y(n_510) );
AND2x2_ASAP7_75t_L g483 ( .A(n_27), .B(n_143), .Y(n_483) );
AOI22xp5_ASAP7_75t_SL g727 ( .A1(n_28), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_28), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_29), .A2(n_132), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_30), .B(n_751), .Y(n_750) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_31), .A2(n_170), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_32), .B(n_139), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_33), .A2(n_132), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_34), .B(n_139), .Y(n_187) );
AND2x2_ASAP7_75t_L g129 ( .A(n_35), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g133 ( .A(n_35), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g241 ( .A(n_35), .Y(n_241) );
OR2x6_ASAP7_75t_L g445 ( .A(n_36), .B(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_L g762 ( .A(n_36), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_38), .B(n_123), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_39), .A2(n_84), .B1(n_132), .B2(n_239), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_40), .B(n_139), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_41), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_42), .B(n_141), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_43), .A2(n_132), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_44), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g533 ( .A(n_45), .B(n_143), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_46), .B(n_143), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_47), .B(n_123), .Y(n_175) );
INVx1_ASAP7_75t_L g126 ( .A(n_48), .Y(n_126) );
INVx1_ASAP7_75t_L g136 ( .A(n_48), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_49), .B(n_139), .Y(n_167) );
AND2x2_ASAP7_75t_L g194 ( .A(n_50), .B(n_143), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_51), .B(n_123), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_52), .B(n_141), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_53), .B(n_141), .Y(n_186) );
AND2x2_ASAP7_75t_L g474 ( .A(n_54), .B(n_143), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_55), .B(n_123), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_56), .B(n_139), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_57), .B(n_123), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_58), .A2(n_132), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_59), .B(n_141), .Y(n_472) );
AND2x2_ASAP7_75t_SL g503 ( .A(n_60), .B(n_144), .Y(n_503) );
AND2x2_ASAP7_75t_L g209 ( .A(n_61), .B(n_144), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_62), .A2(n_132), .B(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_63), .B(n_139), .Y(n_465) );
INVxp33_ASAP7_75t_L g765 ( .A(n_64), .Y(n_765) );
AND2x2_ASAP7_75t_SL g493 ( .A(n_65), .B(n_148), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_66), .B(n_141), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_67), .B(n_141), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_68), .A2(n_95), .B1(n_132), .B2(n_239), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_69), .A2(n_744), .B1(n_748), .B2(n_749), .Y(n_743) );
INVx1_ASAP7_75t_L g749 ( .A(n_69), .Y(n_749) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_70), .A2(n_80), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx14_ASAP7_75t_R g732 ( .A(n_70), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_71), .B(n_139), .Y(n_206) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
INVx1_ASAP7_75t_L g134 ( .A(n_72), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_73), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_74), .A2(n_727), .B1(n_734), .B2(n_736), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_75), .B(n_141), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_76), .A2(n_132), .B(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_77), .A2(n_132), .B(n_137), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_78), .A2(n_132), .B(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g189 ( .A(n_79), .B(n_144), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_80), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_81), .B(n_143), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_82), .B(n_123), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_83), .A2(n_86), .B1(n_123), .B2(n_233), .Y(n_491) );
INVx1_ASAP7_75t_L g448 ( .A(n_85), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_87), .B(n_141), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_88), .B(n_141), .Y(n_523) );
AND2x2_ASAP7_75t_L g147 ( .A(n_89), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_90), .A2(n_132), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_93), .B(n_139), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_94), .A2(n_132), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_96), .B(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g208 ( .A(n_97), .Y(n_208) );
INVxp67_ASAP7_75t_L g513 ( .A(n_98), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_99), .B(n_139), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_100), .A2(n_132), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_101), .B(n_123), .Y(n_532) );
BUFx2_ASAP7_75t_L g109 ( .A(n_102), .Y(n_109) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_755), .B(n_764), .Y(n_103) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_110), .B(n_738), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2x1_ASAP7_75t_R g740 ( .A(n_109), .B(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g110 ( .A1(n_111), .A2(n_727), .B(n_733), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI21x1_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_440), .B(n_449), .Y(n_112) );
AO22x2_ASAP7_75t_L g734 ( .A1(n_113), .A2(n_441), .B1(n_450), .B2(n_735), .Y(n_734) );
INVx4_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_348), .Y(n_114) );
NOR3xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_271), .C(n_306), .Y(n_115) );
OAI211xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_171), .B(n_223), .C(n_261), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_150), .Y(n_118) );
AND2x2_ASAP7_75t_L g254 ( .A(n_119), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_119), .B(n_260), .Y(n_294) );
AND2x2_ASAP7_75t_L g319 ( .A(n_119), .B(n_274), .Y(n_319) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g226 ( .A(n_120), .Y(n_226) );
OR2x2_ASAP7_75t_L g257 ( .A(n_120), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g265 ( .A(n_120), .B(n_161), .Y(n_265) );
AND2x2_ASAP7_75t_L g273 ( .A(n_120), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g300 ( .A(n_120), .B(n_301), .Y(n_300) );
NOR2x1_ASAP7_75t_L g311 ( .A(n_120), .B(n_303), .Y(n_311) );
AND2x4_ASAP7_75t_L g328 ( .A(n_120), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g366 ( .A(n_120), .Y(n_366) );
AND2x4_ASAP7_75t_SL g371 ( .A(n_120), .B(n_151), .Y(n_371) );
OR2x6_ASAP7_75t_L g120 ( .A(n_121), .B(n_147), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_131), .B(n_143), .Y(n_121) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
INVx1_ASAP7_75t_L g516 ( .A(n_124), .Y(n_516) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
AND2x6_ASAP7_75t_L g141 ( .A(n_125), .B(n_134), .Y(n_141) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g139 ( .A(n_127), .B(n_136), .Y(n_139) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx5_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
AND2x2_ASAP7_75t_L g135 ( .A(n_130), .B(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_130), .Y(n_236) );
AND2x6_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
BUFx3_ASAP7_75t_L g237 ( .A(n_133), .Y(n_237) );
INVx2_ASAP7_75t_L g243 ( .A(n_134), .Y(n_243) );
AND2x4_ASAP7_75t_L g239 ( .A(n_135), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g235 ( .A(n_136), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_142), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_141), .B(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_142), .A2(n_157), .B(n_158), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_142), .A2(n_166), .B(n_167), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_142), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_142), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_142), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_142), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_142), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_142), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_142), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_142), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_142), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_142), .A2(n_530), .B(n_531), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_143), .Y(n_153) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_143), .A2(n_232), .B(n_238), .Y(n_231) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_143), .A2(n_520), .B(n_524), .Y(n_519) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g180 ( .A(n_145), .B(n_146), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_148), .A2(n_203), .B(n_204), .Y(n_202) );
INVx2_ASAP7_75t_SL g489 ( .A(n_148), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_148), .A2(n_498), .B(n_499), .Y(n_497) );
BUFx4f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_150), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_150), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_161), .Y(n_150) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_151), .Y(n_266) );
INVx2_ASAP7_75t_L g302 ( .A(n_151), .Y(n_302) );
INVx1_ASAP7_75t_L g329 ( .A(n_151), .Y(n_329) );
AND2x2_ASAP7_75t_L g428 ( .A(n_151), .B(n_338), .Y(n_428) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_152), .Y(n_260) );
AND2x2_ASAP7_75t_L g274 ( .A(n_152), .B(n_161), .Y(n_274) );
AOI21x1_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_160), .Y(n_152) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_153), .A2(n_468), .B(n_474), .Y(n_467) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_153), .A2(n_477), .B(n_483), .Y(n_476) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_153), .A2(n_477), .B(n_483), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_159), .Y(n_154) );
INVx2_ASAP7_75t_L g303 ( .A(n_161), .Y(n_303) );
INVx2_ASAP7_75t_L g338 ( .A(n_161), .Y(n_338) );
OR2x2_ASAP7_75t_L g423 ( .A(n_161), .B(n_255), .Y(n_423) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_169), .Y(n_161) );
INVx4_ASAP7_75t_L g170 ( .A(n_162), .Y(n_170) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_162), .A2(n_527), .B(n_533), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_168), .Y(n_163) );
INVx3_ASAP7_75t_L g182 ( .A(n_170), .Y(n_182) );
AOI211xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_190), .B(n_210), .C(n_217), .Y(n_171) );
INVx2_ASAP7_75t_SL g312 ( .A(n_172), .Y(n_312) );
AND2x2_ASAP7_75t_L g318 ( .A(n_172), .B(n_191), .Y(n_318) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_181), .Y(n_172) );
INVx1_ASAP7_75t_L g214 ( .A(n_173), .Y(n_214) );
INVx1_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
INVx2_ASAP7_75t_L g245 ( .A(n_173), .Y(n_245) );
AND2x2_ASAP7_75t_L g269 ( .A(n_173), .B(n_193), .Y(n_269) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_173), .Y(n_298) );
OR2x2_ASAP7_75t_L g378 ( .A(n_173), .B(n_201), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_180), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_180), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_180), .A2(n_461), .B(n_462), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_180), .B(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_180), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_180), .B(n_513), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_180), .B(n_515), .C(n_516), .Y(n_514) );
AND2x2_ASAP7_75t_L g244 ( .A(n_181), .B(n_245), .Y(n_244) );
NOR2x1_ASAP7_75t_SL g276 ( .A(n_181), .B(n_201), .Y(n_276) );
AO21x1_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_181) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_182), .A2(n_183), .B(n_189), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_188), .Y(n_183) );
INVxp67_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g290 ( .A(n_191), .B(n_213), .Y(n_290) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_201), .Y(n_191) );
OR2x2_ASAP7_75t_L g222 ( .A(n_192), .B(n_201), .Y(n_222) );
BUFx2_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_192), .B(n_298), .Y(n_297) );
INVx4_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_193), .Y(n_249) );
AND2x2_ASAP7_75t_L g275 ( .A(n_193), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g285 ( .A(n_193), .Y(n_285) );
NAND2x1_ASAP7_75t_L g323 ( .A(n_193), .B(n_201), .Y(n_323) );
OR2x2_ASAP7_75t_L g398 ( .A(n_193), .B(n_215), .Y(n_398) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx2_ASAP7_75t_SL g211 ( .A(n_201), .Y(n_211) );
AND2x2_ASAP7_75t_L g270 ( .A(n_201), .B(n_215), .Y(n_270) );
AND2x2_ASAP7_75t_L g341 ( .A(n_201), .B(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g362 ( .A(n_201), .Y(n_362) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_209), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
INVx1_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g284 ( .A(n_213), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
BUFx2_ASAP7_75t_L g279 ( .A(n_214), .Y(n_279) );
AND2x2_ASAP7_75t_L g251 ( .A(n_215), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g342 ( .A(n_215), .Y(n_342) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_221), .Y(n_218) );
OR2x2_ASAP7_75t_L g288 ( .A(n_219), .B(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_SL g330 ( .A(n_219), .B(n_331), .Y(n_330) );
AOI322xp5_ASAP7_75t_L g367 ( .A1(n_219), .A2(n_246), .A3(n_368), .B1(n_370), .B2(n_373), .C1(n_375), .C2(n_377), .Y(n_367) );
AND2x2_ASAP7_75t_L g432 ( .A(n_219), .B(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_220), .B(n_246), .Y(n_256) );
AOI322xp5_ASAP7_75t_L g307 ( .A1(n_221), .A2(n_308), .A3(n_312), .B1(n_313), .B2(n_316), .C1(n_318), .C2(n_319), .Y(n_307) );
INVx2_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g359 ( .A(n_222), .B(n_312), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_222), .A2(n_419), .B1(n_421), .B2(n_424), .Y(n_418) );
OR2x2_ASAP7_75t_L g436 ( .A(n_222), .B(n_385), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_246), .B(n_247), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
AOI221xp5_ASAP7_75t_SL g286 ( .A1(n_225), .A2(n_262), .B1(n_287), .B2(n_290), .C(n_291), .Y(n_286) );
AND2x2_ASAP7_75t_L g313 ( .A(n_225), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_226), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g355 ( .A(n_226), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g384 ( .A(n_227), .Y(n_384) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_244), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_228), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g326 ( .A(n_228), .Y(n_326) );
OR2x2_ASAP7_75t_L g333 ( .A(n_228), .B(n_334), .Y(n_333) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g376 ( .A(n_229), .B(n_338), .Y(n_376) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AND2x4_ASAP7_75t_L g255 ( .A(n_230), .B(n_231), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_233), .A2(n_239), .B1(n_507), .B2(n_509), .Y(n_506) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_237), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NOR2x1p5_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_244), .B(n_305), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_244), .B(n_285), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_244), .Y(n_385) );
INVx1_ASAP7_75t_L g252 ( .A(n_245), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_253), .B1(n_256), .B2(n_257), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_SL g363 ( .A(n_251), .Y(n_363) );
AND2x2_ASAP7_75t_L g420 ( .A(n_252), .B(n_276), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_254), .B(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_SL g292 ( .A(n_254), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_254), .B(n_413), .Y(n_412) );
BUFx3_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
INVx2_ASAP7_75t_L g310 ( .A(n_255), .Y(n_310) );
AND2x2_ASAP7_75t_L g353 ( .A(n_255), .B(n_337), .Y(n_353) );
INVx1_ASAP7_75t_L g267 ( .A(n_257), .Y(n_267) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI21xp5_ASAP7_75t_SL g261 ( .A1(n_262), .A2(n_267), .B(n_268), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g346 ( .A(n_265), .Y(n_346) );
INVx2_ASAP7_75t_L g334 ( .A(n_266), .Y(n_334) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x2_ASAP7_75t_L g331 ( .A(n_270), .B(n_285), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_270), .A2(n_368), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_272), .B(n_286), .Y(n_271) );
AOI32xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_275), .A3(n_277), .B1(n_281), .B2(n_284), .Y(n_272) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_273), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_273), .A2(n_362), .B1(n_380), .B2(n_382), .C(n_388), .Y(n_379) );
AND2x2_ASAP7_75t_L g399 ( .A(n_273), .B(n_280), .Y(n_399) );
BUFx2_ASAP7_75t_L g283 ( .A(n_274), .Y(n_283) );
INVx1_ASAP7_75t_L g408 ( .A(n_274), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_274), .Y(n_413) );
INVx1_ASAP7_75t_SL g406 ( .A(n_275), .Y(n_406) );
INVx2_ASAP7_75t_L g289 ( .A(n_276), .Y(n_289) );
AND2x2_ASAP7_75t_L g401 ( .A(n_277), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g373 ( .A(n_279), .B(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g345 ( .A(n_280), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_280), .B(n_371), .Y(n_393) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g305 ( .A(n_285), .Y(n_305) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g295 ( .A(n_289), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g304 ( .A(n_289), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g409 ( .A(n_290), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B1(n_299), .B2(n_304), .Y(n_291) );
INVx2_ASAP7_75t_SL g383 ( .A(n_293), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_293), .B(n_422), .Y(n_424) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_295), .A2(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g340 ( .A(n_297), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g368 ( .A(n_300), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g315 ( .A(n_301), .Y(n_315) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g357 ( .A(n_303), .Y(n_357) );
INVx1_ASAP7_75t_L g402 ( .A(n_304), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_320), .C(n_343), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx2_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
AND2x2_ASAP7_75t_L g387 ( .A(n_309), .B(n_328), .Y(n_387) );
OR2x2_ASAP7_75t_L g426 ( .A(n_309), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_310), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g322 ( .A(n_312), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g389 ( .A(n_315), .B(n_326), .Y(n_389) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_318), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g430 ( .A(n_318), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_324), .B1(n_328), .B2(n_330), .C(n_332), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_321), .A2(n_344), .B(n_347), .Y(n_343) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx3_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_323), .B(n_417), .Y(n_416) );
INVxp33_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g335 ( .A(n_331), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_336), .B2(n_339), .Y(n_332) );
INVx2_ASAP7_75t_L g438 ( .A(n_334), .Y(n_438) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVxp67_ASAP7_75t_L g417 ( .A(n_342), .Y(n_417) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NOR2x1_ASAP7_75t_L g348 ( .A(n_349), .B(n_394), .Y(n_348) );
NAND4xp25_ASAP7_75t_L g349 ( .A(n_350), .B(n_367), .C(n_379), .D(n_391), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B(n_358), .C(n_360), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_355), .A2(n_361), .B(n_364), .Y(n_360) );
INVx2_ASAP7_75t_L g439 ( .A(n_356), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_357), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g372 ( .A(n_357), .Y(n_372) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
OR2x2_ASAP7_75t_L g434 ( .A(n_362), .B(n_398), .Y(n_434) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_369), .Y(n_405) );
AND2x2_ASAP7_75t_SL g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x2_ASAP7_75t_L g375 ( .A(n_371), .B(n_376), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_371), .A2(n_401), .B(n_403), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_371), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g429 ( .A(n_371), .Y(n_429) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI22xp33_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_384), .B1(n_385), .B2(n_386), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_395), .B(n_400), .C(n_410), .D(n_431), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_407), .B2(n_409), .Y(n_403) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI211xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_414), .B(n_418), .C(n_425), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_429), .B(n_430), .Y(n_425) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
OAI21xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_435), .B(n_437), .Y(n_431) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
CKINVDCx11_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
OR2x6_ASAP7_75t_SL g442 ( .A(n_443), .B(n_444), .Y(n_442) );
AND2x6_ASAP7_75t_SL g450 ( .A(n_443), .B(n_445), .Y(n_450) );
OR2x2_ASAP7_75t_L g737 ( .A(n_443), .B(n_445), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_443), .B(n_444), .Y(n_742) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_447), .B(n_448), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx2_ASAP7_75t_L g735 ( .A(n_451), .Y(n_735) );
XNOR2xp5_ASAP7_75t_L g744 ( .A(n_451), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_649), .Y(n_451) );
NOR3xp33_ASAP7_75t_SL g452 ( .A(n_453), .B(n_573), .C(n_623), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_553), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_494), .B(n_534), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_484), .Y(n_456) );
INVx1_ASAP7_75t_SL g659 ( .A(n_457), .Y(n_659) );
AOI32xp33_ASAP7_75t_L g690 ( .A1(n_457), .A2(n_672), .A3(n_691), .B1(n_692), .B2(n_693), .Y(n_690) );
AND2x2_ASAP7_75t_L g692 ( .A(n_457), .B(n_549), .Y(n_692) );
AND2x4_ASAP7_75t_SL g457 ( .A(n_458), .B(n_466), .Y(n_457) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_458), .Y(n_485) );
INVx5_ASAP7_75t_L g552 ( .A(n_458), .Y(n_552) );
OR2x2_ASAP7_75t_L g559 ( .A(n_458), .B(n_551), .Y(n_559) );
INVx2_ASAP7_75t_L g564 ( .A(n_458), .Y(n_564) );
AND2x2_ASAP7_75t_L g576 ( .A(n_458), .B(n_467), .Y(n_576) );
AND2x2_ASAP7_75t_L g581 ( .A(n_458), .B(n_475), .Y(n_581) );
OR2x2_ASAP7_75t_L g588 ( .A(n_458), .B(n_487), .Y(n_588) );
AND2x4_ASAP7_75t_L g597 ( .A(n_458), .B(n_476), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_SL g639 ( .A1(n_458), .A2(n_555), .B(n_590), .C(n_628), .Y(n_639) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx3_ASAP7_75t_SL g589 ( .A(n_466), .Y(n_589) );
AND2x2_ASAP7_75t_L g635 ( .A(n_466), .B(n_552), .Y(n_635) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
AND2x2_ASAP7_75t_L g486 ( .A(n_467), .B(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g566 ( .A(n_467), .B(n_476), .Y(n_566) );
AND2x2_ASAP7_75t_L g570 ( .A(n_467), .B(n_549), .Y(n_570) );
INVx1_ASAP7_75t_L g596 ( .A(n_467), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_467), .B(n_476), .Y(n_618) );
INVx2_ASAP7_75t_L g622 ( .A(n_467), .Y(n_622) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_467), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_467), .B(n_552), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g633 ( .A(n_476), .B(n_487), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g643 ( .A(n_485), .Y(n_643) );
NAND2xp33_ASAP7_75t_SL g668 ( .A(n_485), .B(n_560), .Y(n_668) );
AND2x2_ASAP7_75t_L g710 ( .A(n_486), .B(n_552), .Y(n_710) );
AND2x2_ASAP7_75t_L g621 ( .A(n_487), .B(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g684 ( .A(n_487), .Y(n_684) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_488), .Y(n_549) );
AOI21x1_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_493), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_494), .A2(n_575), .B1(n_677), .B2(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_517), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_495), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_495), .B(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_504), .Y(n_495) );
INVx2_ASAP7_75t_L g540 ( .A(n_496), .Y(n_540) );
OR2x2_ASAP7_75t_L g544 ( .A(n_496), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_496), .B(n_557), .Y(n_562) );
AND2x4_ASAP7_75t_SL g572 ( .A(n_496), .B(n_505), .Y(n_572) );
OR2x2_ASAP7_75t_L g579 ( .A(n_496), .B(n_519), .Y(n_579) );
OR2x2_ASAP7_75t_L g591 ( .A(n_496), .B(n_505), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_496), .B(n_519), .Y(n_605) );
INVx1_ASAP7_75t_L g610 ( .A(n_496), .Y(n_610) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_496), .Y(n_628) );
AND2x2_ASAP7_75t_L g691 ( .A(n_496), .B(n_611), .Y(n_691) );
INVx2_ASAP7_75t_L g695 ( .A(n_496), .Y(n_695) );
OR2x2_ASAP7_75t_L g702 ( .A(n_496), .B(n_592), .Y(n_702) );
OR2x2_ASAP7_75t_L g724 ( .A(n_496), .B(n_725), .Y(n_724) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
AND2x2_ASAP7_75t_L g541 ( .A(n_504), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_504), .B(n_525), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_504), .B(n_601), .Y(n_663) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g560 ( .A(n_505), .Y(n_560) );
AND2x4_ASAP7_75t_L g611 ( .A(n_505), .B(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_505), .B(n_556), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_505), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_505), .B(n_545), .Y(n_704) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
AND2x2_ASAP7_75t_L g571 ( .A(n_517), .B(n_572), .Y(n_571) );
AO221x1_ASAP7_75t_L g645 ( .A1(n_517), .A2(n_560), .B1(n_591), .B2(n_646), .C(n_647), .Y(n_645) );
OAI322xp33_ASAP7_75t_L g697 ( .A1(n_517), .A2(n_617), .A3(n_698), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_703), .Y(n_697) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_525), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g539 ( .A(n_519), .Y(n_539) );
INVx2_ASAP7_75t_L g545 ( .A(n_519), .Y(n_545) );
AND2x2_ASAP7_75t_L g557 ( .A(n_519), .B(n_525), .Y(n_557) );
INVx1_ASAP7_75t_L g602 ( .A(n_519), .Y(n_602) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_519), .Y(n_658) );
INVx1_ASAP7_75t_L g542 ( .A(n_525), .Y(n_542) );
OR2x2_ASAP7_75t_L g592 ( .A(n_525), .B(n_545), .Y(n_592) );
INVx2_ASAP7_75t_L g612 ( .A(n_525), .Y(n_612) );
INVx1_ASAP7_75t_L g665 ( .A(n_525), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_525), .B(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .Y(n_527) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI21xp33_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_543), .B(n_546), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_536), .A2(n_575), .B1(n_577), .B2(n_581), .C(n_582), .Y(n_574) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .Y(n_537) );
NOR2x1p5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g661 ( .A(n_540), .Y(n_661) );
INVx1_ASAP7_75t_SL g580 ( .A(n_541), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_541), .A2(n_686), .B(n_688), .Y(n_685) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_542), .Y(n_585) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_545), .Y(n_648) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
OAI211xp5_ASAP7_75t_L g623 ( .A1(n_548), .A2(n_624), .B(n_629), .C(n_640), .Y(n_623) );
OR2x2_ASAP7_75t_L g713 ( .A(n_548), .B(n_618), .Y(n_713) );
AND2x2_ASAP7_75t_L g715 ( .A(n_548), .B(n_581), .Y(n_715) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g555 ( .A(n_549), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g617 ( .A(n_549), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g655 ( .A(n_549), .B(n_622), .Y(n_655) );
OA33x2_ASAP7_75t_L g662 ( .A1(n_549), .A2(n_579), .A3(n_663), .B1(n_664), .B2(n_666), .B3(n_668), .Y(n_662) );
OR2x2_ASAP7_75t_L g673 ( .A(n_549), .B(n_658), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_549), .B(n_597), .Y(n_687) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g575 ( .A(n_551), .B(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_551), .A2(n_581), .B1(n_625), .B2(n_626), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_552), .B(n_632), .C(n_665), .Y(n_664) );
AOI322xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_558), .A3(n_560), .B1(n_561), .B2(n_563), .C1(n_567), .C2(n_571), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g660 ( .A(n_556), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g615 ( .A1(n_557), .A2(n_572), .B(n_616), .C(n_619), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_558), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
NAND4xp25_ASAP7_75t_SL g679 ( .A(n_559), .B(n_588), .C(n_680), .D(n_682), .Y(n_679) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g569 ( .A(n_564), .Y(n_569) );
OR2x2_ASAP7_75t_L g614 ( .A(n_564), .B(n_566), .Y(n_614) );
AND2x2_ASAP7_75t_L g683 ( .A(n_565), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g688 ( .A(n_569), .B(n_683), .Y(n_688) );
BUFx2_ASAP7_75t_L g681 ( .A(n_570), .Y(n_681) );
INVx1_ASAP7_75t_SL g711 ( .A(n_571), .Y(n_711) );
AND2x4_ASAP7_75t_L g647 ( .A(n_572), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g700 ( .A(n_572), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_593), .C(n_615), .Y(n_573) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_SL g637 ( .A(n_579), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_579), .A2(n_706), .B(n_707), .C(n_716), .Y(n_705) );
OR2x2_ASAP7_75t_L g627 ( .A(n_580), .B(n_628), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_586), .B1(n_589), .B2(n_590), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_584), .B(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_587), .B(n_644), .Y(n_726) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g701 ( .A(n_588), .B(n_589), .Y(n_701) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g646 ( .A(n_592), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_598), .B1(n_603), .B2(n_607), .C1(n_608), .C2(n_613), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_596), .Y(n_607) );
AND2x2_ASAP7_75t_L g654 ( .A(n_597), .B(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_597), .A2(n_670), .B1(n_675), .B2(n_679), .Y(n_669) );
INVx2_ASAP7_75t_SL g722 ( .A(n_597), .Y(n_722) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g678 ( .A(n_602), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_602), .B(n_665), .Y(n_725) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g638 ( .A(n_606), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_608), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g676 ( .A(n_610), .Y(n_676) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_611), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g719 ( .A(n_611), .B(n_648), .Y(n_719) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g644 ( .A(n_618), .Y(n_644) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g723 ( .A(n_621), .Y(n_723) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_622), .Y(n_667) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_634), .B(n_636), .C(n_639), .Y(n_629) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g674 ( .A(n_636), .Y(n_674) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_645), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_689), .C(n_705), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_669), .C(n_685), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B1(n_659), .B2(n_660), .C(n_662), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_674), .Y(n_670) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g698 ( .A(n_684), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g706 ( .A(n_688), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_696), .Y(n_689) );
INVx2_ASAP7_75t_L g712 ( .A(n_691), .Y(n_712) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g703 ( .A(n_694), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B1(n_712), .B2(n_713), .C(n_714), .Y(n_708) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_720), .B1(n_724), .B2(n_726), .Y(n_717) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI21xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_743), .B(n_750), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
BUFx3_ASAP7_75t_L g754 ( .A(n_742), .Y(n_754) );
INVx2_ASAP7_75t_L g748 ( .A(n_744), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
CKINVDCx11_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_756), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx3_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_759), .B(n_763), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
endmodule