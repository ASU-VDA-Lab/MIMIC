module fake_jpeg_744_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_38),
.Y(n_59)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_35),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_30),
.B1(n_35),
.B2(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_49),
.B1(n_48),
.B2(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_30),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_60),
.C(n_61),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_37),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_65),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_58),
.B1(n_57),
.B2(n_60),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_47),
.B(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_47),
.B1(n_15),
.B2(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_65),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_78),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_13),
.C(n_28),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_76),
.C(n_23),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_47),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_1),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_26),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_25),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_24),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_92),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_88),
.C(n_93),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_91),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_81),
.C(n_82),
.Y(n_93)
);

OAI322xp33_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_21),
.A3(n_20),
.B1(n_18),
.B2(n_11),
.C1(n_7),
.C2(n_3),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_86),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_98),
.C(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_99),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_87),
.C(n_97),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_90),
.C(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

OAI221xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_4),
.C(n_8),
.Y(n_108)
);


endmodule