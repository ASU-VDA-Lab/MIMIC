module fake_jpeg_12264_n_420 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_420);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_420;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_45),
.Y(n_100)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_47),
.B(n_59),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_0),
.B(n_1),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_53),
.C(n_24),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_60),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_31),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_0),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_18),
.B(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_65),
.Y(n_102)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_21),
.B(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_76),
.Y(n_122)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx2_ASAP7_75t_SL g115 ( 
.A(n_77),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_30),
.B(n_15),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_79),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_35),
.Y(n_83)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_83),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_42),
.B1(n_25),
.B2(n_38),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_88),
.A2(n_94),
.B1(n_117),
.B2(n_118),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_42),
.B1(n_25),
.B2(n_29),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_107),
.B1(n_120),
.B2(n_20),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_42),
.B1(n_25),
.B2(n_29),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_95),
.B(n_113),
.Y(n_163)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_26),
.B1(n_34),
.B2(n_29),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_105),
.B1(n_119),
.B2(n_73),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_30),
.B1(n_21),
.B2(n_19),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_82),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_26),
.B1(n_19),
.B2(n_68),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_25),
.B1(n_42),
.B2(n_41),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_49),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_48),
.A2(n_43),
.B1(n_40),
.B2(n_28),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_62),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_51),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_53),
.B(n_52),
.C(n_72),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_131),
.A2(n_153),
.B1(n_161),
.B2(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_50),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_110),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_73),
.B(n_57),
.C(n_44),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_83),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_141),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_80),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_143),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_84),
.B1(n_116),
.B2(n_112),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_144),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_93),
.A2(n_79),
.B(n_61),
.C(n_76),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_70),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_46),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_85),
.B(n_73),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_146),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_150),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_86),
.B(n_69),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

OR2x2_ASAP7_75t_SL g151 ( 
.A(n_104),
.B(n_55),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_152),
.C(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_63),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_101),
.A2(n_81),
.B1(n_75),
.B2(n_66),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_14),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_156),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_35),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_14),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_160),
.Y(n_191)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_91),
.B(n_2),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_10),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_96),
.A2(n_111),
.B1(n_108),
.B2(n_106),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_90),
.A2(n_77),
.B1(n_35),
.B2(n_5),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_103),
.B(n_77),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_177),
.Y(n_205)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_100),
.A3(n_77),
.B1(n_90),
.B2(n_97),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_192),
.B(n_195),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_193),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_134),
.B1(n_133),
.B2(n_156),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_146),
.A2(n_100),
.B1(n_123),
.B2(n_121),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_148),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_139),
.A2(n_123),
.B1(n_121),
.B2(n_109),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_156),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_137),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_201),
.C(n_207),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_138),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_199),
.B(n_203),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_194),
.A2(n_152),
.B(n_163),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_219),
.B(n_225),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_163),
.C(n_144),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_143),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_193),
.B1(n_179),
.B2(n_183),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_186),
.C(n_163),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_134),
.B1(n_130),
.B2(n_135),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_208),
.A2(n_221),
.B1(n_188),
.B2(n_192),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_140),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_220),
.C(n_174),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_216),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_141),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_141),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_223),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_151),
.B(n_129),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_129),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_159),
.B1(n_154),
.B2(n_136),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_155),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_183),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_188),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_154),
.B(n_160),
.Y(n_225)
);

INVxp33_ASAP7_75t_SL g228 ( 
.A(n_214),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_181),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_241),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_221),
.A2(n_185),
.B1(n_187),
.B2(n_195),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_245),
.B1(n_224),
.B2(n_204),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_235),
.A2(n_242),
.B1(n_136),
.B2(n_157),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_243),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_180),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_239),
.C(n_248),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_181),
.C(n_169),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_191),
.A3(n_173),
.B1(n_176),
.B2(n_182),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_191),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_185),
.B1(n_171),
.B2(n_196),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_205),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_247),
.A2(n_208),
.B(n_223),
.Y(n_269)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_174),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_252),
.C(n_219),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_200),
.B(n_176),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_210),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_253),
.B(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_203),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_256),
.B(n_267),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_257),
.A2(n_273),
.B1(n_279),
.B2(n_282),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_237),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_244),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_275),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_206),
.C(n_225),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_265),
.C(n_251),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_206),
.C(n_209),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_199),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_269),
.B(n_283),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_211),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_211),
.Y(n_272)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

AOI22x1_ASAP7_75t_L g273 ( 
.A1(n_233),
.A2(n_149),
.B1(n_222),
.B2(n_198),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_232),
.Y(n_274)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_239),
.B1(n_252),
.B2(n_241),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_277),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_231),
.A2(n_190),
.B1(n_198),
.B2(n_149),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_229),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_284),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_234),
.A2(n_149),
.B1(n_190),
.B2(n_168),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_242),
.A2(n_178),
.B(n_170),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_232),
.A2(n_248),
.B1(n_238),
.B2(n_254),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_262),
.B1(n_260),
.B2(n_257),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_258),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_291),
.B(n_296),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_230),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_311),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_300),
.C(n_306),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_258),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_249),
.Y(n_297)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_190),
.B1(n_158),
.B2(n_116),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_303),
.A2(n_279),
.B1(n_281),
.B2(n_280),
.Y(n_313)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_165),
.C(n_161),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_268),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_307),
.B(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_278),
.B1(n_270),
.B2(n_273),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_161),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_286),
.A2(n_275),
.B(n_272),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_312),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_304),
.B1(n_301),
.B2(n_289),
.Y(n_346)
);

XNOR2x1_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_264),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_316),
.C(n_321),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_265),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_261),
.C(n_271),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_317),
.B(n_168),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_276),
.B1(n_259),
.B2(n_283),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_318),
.A2(n_323),
.B1(n_324),
.B2(n_327),
.Y(n_352)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_292),
.A2(n_273),
.B1(n_278),
.B2(n_158),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_292),
.A2(n_285),
.B1(n_293),
.B2(n_299),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_326),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_299),
.A2(n_168),
.B1(n_109),
.B2(n_87),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_108),
.C(n_103),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_332),
.C(n_308),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_87),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_336),
.B(n_342),
.Y(n_369)
);

BUFx12_ASAP7_75t_L g340 ( 
.A(n_313),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_340),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_306),
.C(n_286),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_341),
.B(n_344),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_312),
.A2(n_333),
.B(n_310),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_318),
.A2(n_297),
.B(n_298),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_343),
.B(n_345),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_302),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_302),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_311),
.B1(n_298),
.B2(n_302),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_348),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_315),
.A2(n_302),
.B1(n_288),
.B2(n_303),
.Y(n_348)
);

NOR2x1_ASAP7_75t_L g358 ( 
.A(n_351),
.B(n_331),
.Y(n_358)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_330),
.Y(n_353)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_353),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_161),
.Y(n_354)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_349),
.A2(n_323),
.B(n_327),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_357),
.Y(n_379)
);

NAND2x1_ASAP7_75t_SL g357 ( 
.A(n_350),
.B(n_315),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_340),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_352),
.A2(n_329),
.B1(n_332),
.B2(n_314),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_365),
.B1(n_366),
.B2(n_339),
.Y(n_372)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_353),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_363),
.A2(n_349),
.B1(n_350),
.B2(n_338),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_337),
.A2(n_112),
.B1(n_125),
.B2(n_124),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_337),
.A2(n_125),
.B1(n_124),
.B2(n_92),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_161),
.C(n_111),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_335),
.C(n_340),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_106),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_370),
.Y(n_382)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_372),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_376),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_338),
.B1(n_342),
.B2(n_336),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_360),
.B1(n_368),
.B2(n_357),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_348),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_378),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_356),
.A2(n_346),
.B1(n_347),
.B2(n_340),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_362),
.A2(n_335),
.B(n_343),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_381),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_380),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_84),
.C(n_115),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_371),
.A2(n_10),
.B(n_14),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_383),
.B(n_384),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_358),
.A2(n_13),
.B(n_12),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_84),
.C(n_35),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_370),
.C(n_355),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_379),
.A2(n_361),
.B(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_395),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_390),
.A2(n_382),
.B1(n_13),
.B2(n_12),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_380),
.B(n_359),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_394),
.B(n_385),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_365),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_396),
.B(n_366),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_378),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_400),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_403),
.C(n_401),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_389),
.C(n_388),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_402),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_392),
.Y(n_402)
);

AOI21x1_ASAP7_75t_L g403 ( 
.A1(n_395),
.A2(n_381),
.B(n_382),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_404),
.A2(n_405),
.B1(n_393),
.B2(n_13),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_393),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_407),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_398),
.Y(n_409)
);

A2O1A1O1Ixp25_ASAP7_75t_L g415 ( 
.A1(n_409),
.A2(n_410),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_404),
.A2(n_11),
.B(n_4),
.Y(n_411)
);

OAI21xp33_ASAP7_75t_L g414 ( 
.A1(n_411),
.A2(n_4),
.B(n_5),
.Y(n_414)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g412 ( 
.A1(n_406),
.A2(n_3),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_412),
.A2(n_414),
.B1(n_408),
.B2(n_7),
.Y(n_416)
);

AOI21x1_ASAP7_75t_L g417 ( 
.A1(n_415),
.A2(n_6),
.B(n_8),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_416),
.B(n_417),
.C(n_413),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_9),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_419),
.B(n_9),
.Y(n_420)
);


endmodule