module real_jpeg_24721_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_1),
.A2(n_56),
.B1(n_67),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_1),
.A2(n_26),
.B1(n_29),
.B2(n_71),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_71),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_5),
.A2(n_26),
.B1(n_29),
.B2(n_46),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_5),
.A2(n_46),
.B1(n_63),
.B2(n_64),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_6),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_26),
.B1(n_29),
.B2(n_76),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_6),
.A2(n_57),
.B1(n_68),
.B2(n_76),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_76),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_7),
.B(n_69),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_7),
.B(n_26),
.C(n_40),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_106),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_7),
.B(n_85),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_7),
.A2(n_25),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_10),
.A2(n_67),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_10),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_115),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_115),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_10),
.A2(n_26),
.B1(n_29),
.B2(n_115),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_11),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_58),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_11),
.A2(n_26),
.B1(n_29),
.B2(n_58),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_26),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_13),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_13),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_14),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_14),
.A2(n_30),
.B1(n_43),
.B2(n_44),
.Y(n_96)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_15),
.Y(n_103)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_15),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_144),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_143),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_20),
.B(n_120),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_86),
.C(n_97),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_23),
.B(n_54),
.C(n_72),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_24),
.B(n_37),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_31),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_25),
.B(n_35),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_25),
.A2(n_28),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_25),
.A2(n_33),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_25),
.A2(n_90),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_25),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_25),
.A2(n_206),
.B1(n_213),
.B2(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_27),
.Y(n_178)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_27),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_29),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_32),
.A2(n_92),
.B(n_204),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B(n_47),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_38),
.A2(n_42),
.B1(n_50),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_38),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_38),
.A2(n_50),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_38),
.A2(n_50),
.B1(n_191),
.B2(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_38),
.B(n_106),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_51)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_44),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_43),
.B(n_64),
.C(n_81),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_44),
.B(n_187),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_44),
.A2(n_80),
.B(n_231),
.C(n_232),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_48),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_49),
.A2(n_128),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_50),
.A2(n_96),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_50),
.A2(n_127),
.B(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_50),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_72),
.B2(n_73),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_69),
.B2(n_70),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_55),
.Y(n_119)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_62),
.C(n_63),
.Y(n_107)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_59),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_59),
.A2(n_69),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_60),
.A2(n_113),
.B1(n_114),
.B2(n_119),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_64),
.B(n_105),
.C(n_107),
.Y(n_104)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_64),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g231 ( 
.A(n_64),
.B(n_106),
.CON(n_231),
.SN(n_231)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_68),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_69),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_70),
.Y(n_134)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B(n_83),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_85),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_109),
.B(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_79),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_84),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_78),
.A2(n_85),
.B1(n_110),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_78),
.A2(n_85),
.B1(n_172),
.B2(n_231),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_79),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_86),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_94),
.B2(n_95),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_92),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_93),
.A2(n_102),
.B(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_97),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.C(n_112),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_98),
.A2(n_99),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_104),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_106),
.B(n_116),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_106),
.B(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_108),
.B(n_112),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_142),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_130),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_129),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_128),
.B(n_155),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_179),
.B(n_264),
.C(n_269),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_164),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_146),
.B(n_164),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_161),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_148),
.B(n_151),
.C(n_161),
.Y(n_265)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.C(n_158),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_165),
.B(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_168),
.B(n_169),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.C(n_176),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_170),
.B(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_248)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_263),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_258),
.B(n_262),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_243),
.B(n_257),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_227),
.B(n_242),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_201),
.B(n_226),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_192),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_188),
.B1(n_189),
.B2(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_200),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_210),
.B(n_225),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_208),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_221),
.B(n_224),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_241),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_241),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_237),
.C(n_240),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_239),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_244),
.B(n_245),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_252),
.C(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_252),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);


endmodule