module fake_jpeg_761_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

AND2x6_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_4),
.Y(n_12)
);

OAI21xp33_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_3),
.B(n_10),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_17),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_15),
.B1(n_7),
.B2(n_6),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_16),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_11),
.B1(n_10),
.B2(n_8),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_14),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_14),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_18),
.C(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_14),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_19),
.B1(n_18),
.B2(n_8),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_29),
.B(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_23),
.Y(n_33)
);

MAJx2_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_16),
.C(n_3),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_33),
.B(n_34),
.Y(n_36)
);


endmodule