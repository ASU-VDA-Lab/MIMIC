module fake_jpeg_18217_n_68 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_40),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_12),
.B1(n_27),
.B2(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_1),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_36),
.B(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_48),
.B1(n_50),
.B2(n_3),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_33),
.C(n_30),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_39),
.C(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_46),
.B1(n_51),
.B2(n_49),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.C(n_16),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_11),
.B(n_5),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_18),
.C(n_6),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_20),
.C(n_8),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_9),
.C(n_10),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_21),
.B(n_24),
.C(n_28),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_4),
.Y(n_68)
);


endmodule