module fake_netlist_6_3950_n_835 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_835);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_835;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_796;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_24),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_72),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_45),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_78),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g192 ( 
.A(n_110),
.B(n_115),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_130),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_108),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_92),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_12),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_65),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_152),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_47),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_95),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_41),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_96),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_121),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_3),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_139),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_74),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_17),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_11),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_0),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_102),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_54),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_46),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_86),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_89),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_148),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_179),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_33),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_109),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_124),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_71),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_84),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_85),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_63),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_68),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_L g236 ( 
.A(n_73),
.B(n_136),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_44),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_69),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_70),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_88),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_167),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_16),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_5),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_34),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_61),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_18),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_161),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_38),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g253 ( 
.A1(n_200),
.A2(n_0),
.B(n_1),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_213),
.A2(n_1),
.B(n_2),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_20),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_209),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_184),
.Y(n_266)
);

BUFx8_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_189),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_2),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_191),
.Y(n_274)
);

CKINVDCx6p67_ASAP7_75t_R g275 ( 
.A(n_211),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_197),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_198),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_216),
.B(n_4),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_21),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_222),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_229),
.Y(n_286)
);

BUFx8_ASAP7_75t_L g287 ( 
.A(n_193),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_233),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_239),
.B(n_4),
.Y(n_291)
);

AND2x6_ASAP7_75t_L g292 ( 
.A(n_235),
.B(n_22),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_239),
.B(n_5),
.Y(n_293)
);

OAI22x1_ASAP7_75t_SL g294 ( 
.A1(n_249),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_246),
.B(n_6),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_248),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_192),
.B(n_23),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_184),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_212),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_252),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_194),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_255),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_265),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_293),
.A2(n_225),
.B1(n_245),
.B2(n_218),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_263),
.A2(n_236),
.B(n_218),
.C(n_245),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

AO21x2_ASAP7_75t_L g320 ( 
.A1(n_279),
.A2(n_251),
.B(n_195),
.Y(n_320)
);

AO21x2_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_196),
.B(n_187),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_275),
.A2(n_225),
.B1(n_241),
.B2(n_231),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_256),
.Y(n_325)
);

CKINVDCx6p67_ASAP7_75t_R g326 ( 
.A(n_275),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_256),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_L g329 ( 
.A(n_273),
.B(n_242),
.C(n_230),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_266),
.B(n_227),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_263),
.B(n_202),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_263),
.B(n_203),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_300),
.B(n_282),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_300),
.B(n_204),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_268),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_282),
.B(n_205),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_268),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

NOR2x1p5_ASAP7_75t_L g343 ( 
.A(n_302),
.B(n_206),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_266),
.B(n_224),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_287),
.A2(n_276),
.B1(n_289),
.B2(n_260),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_207),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_287),
.B(n_208),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_276),
.B(n_210),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_219),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_298),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_270),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_296),
.Y(n_355)
);

NOR2x1p5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_302),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_309),
.B(n_296),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_299),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_264),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_325),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_297),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_299),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_273),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_287),
.Y(n_367)
);

BUFx8_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g369 ( 
.A1(n_317),
.A2(n_253),
.B1(n_258),
.B2(n_259),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_297),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_341),
.A2(n_253),
.B1(n_258),
.B2(n_292),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_299),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_334),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_343),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_347),
.A2(n_258),
.B1(n_253),
.B2(n_288),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_345),
.B(n_267),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_323),
.B(n_267),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_299),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_303),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_327),
.B(n_299),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_261),
.Y(n_382)
);

O2A1O1Ixp5_ASAP7_75t_L g383 ( 
.A1(n_331),
.A2(n_285),
.B(n_290),
.C(n_274),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_338),
.B(n_269),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_283),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_332),
.A2(n_292),
.B1(n_285),
.B2(n_284),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_354),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_332),
.B(n_292),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_344),
.B(n_270),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_320),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_305),
.B(n_285),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_321),
.A2(n_292),
.B1(n_272),
.B2(n_286),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_311),
.B(n_270),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_307),
.B(n_267),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_335),
.B(n_270),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_307),
.B(n_223),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_271),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_318),
.B(n_271),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_304),
.A2(n_294),
.B1(n_286),
.B2(n_278),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_307),
.B(n_346),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_318),
.B(n_271),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_304),
.B(n_271),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_272),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_321),
.B(n_272),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_314),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_315),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_321),
.B(n_272),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_313),
.B(n_277),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_315),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_339),
.B(n_277),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_303),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_316),
.B(n_277),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_326),
.B(n_277),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_349),
.B(n_278),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_303),
.B(n_278),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_306),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_L g419 ( 
.A(n_347),
.B(n_286),
.C(n_278),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_313),
.B(n_286),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_353),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_322),
.B(n_324),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_322),
.B(n_25),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_313),
.B(n_9),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_306),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_358),
.A2(n_313),
.B(n_324),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_363),
.B(n_313),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_342),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_366),
.A2(n_352),
.B1(n_350),
.B2(n_342),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_357),
.B(n_10),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_365),
.A2(n_340),
.B(n_336),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_366),
.B(n_10),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_371),
.B(n_336),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_373),
.A2(n_340),
.B(n_310),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_390),
.A2(n_312),
.B1(n_310),
.B2(n_308),
.Y(n_437)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_400),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_418),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_385),
.B(n_11),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_382),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_425),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_379),
.A2(n_381),
.B(n_388),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_385),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

O2A1O1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_369),
.A2(n_308),
.B(n_13),
.C(n_14),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_355),
.A2(n_101),
.B(n_182),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_395),
.A2(n_100),
.B(n_181),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_372),
.A2(n_99),
.B(n_180),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_389),
.B(n_26),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_368),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_384),
.B(n_415),
.Y(n_453)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_405),
.A2(n_103),
.B(n_178),
.Y(n_454)
);

AO22x1_ASAP7_75t_L g455 ( 
.A1(n_375),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_406),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_397),
.A2(n_104),
.B(n_177),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_389),
.A2(n_98),
.B(n_176),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_367),
.B(n_15),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_360),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_27),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_356),
.Y(n_462)
);

AOI21x1_ASAP7_75t_L g463 ( 
.A1(n_408),
.A2(n_106),
.B(n_174),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_403),
.B(n_28),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_396),
.B(n_15),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_359),
.B(n_16),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_419),
.B(n_17),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_364),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_377),
.B(n_18),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_398),
.B(n_19),
.Y(n_471)
);

OAI321xp33_ASAP7_75t_L g472 ( 
.A1(n_369),
.A2(n_19),
.A3(n_29),
.B1(n_30),
.B2(n_31),
.C(n_32),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_404),
.A2(n_35),
.B(n_36),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_372),
.B(n_37),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_394),
.B(n_39),
.Y(n_475)
);

NAND2x1p5_ASAP7_75t_L g476 ( 
.A(n_391),
.B(n_40),
.Y(n_476)
);

AND2x2_ASAP7_75t_SL g477 ( 
.A(n_386),
.B(n_42),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_409),
.A2(n_43),
.B(n_48),
.Y(n_478)
);

AO21x1_ASAP7_75t_L g479 ( 
.A1(n_376),
.A2(n_49),
.B(n_50),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_376),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_392),
.A2(n_55),
.B(n_56),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_L g482 ( 
.A1(n_383),
.A2(n_401),
.B(n_386),
.C(n_392),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_399),
.B(n_57),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_420),
.A2(n_58),
.B(n_59),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_421),
.A2(n_378),
.B1(n_362),
.B2(n_374),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_361),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_417),
.A2(n_60),
.B(n_62),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_422),
.A2(n_64),
.B(n_66),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_411),
.B(n_67),
.Y(n_489)
);

O2A1O1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_383),
.A2(n_423),
.B(n_413),
.C(n_416),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_393),
.B(n_75),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_407),
.A2(n_77),
.B(n_79),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_416),
.B(n_80),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_414),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_410),
.A2(n_412),
.B(n_380),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_412),
.A2(n_81),
.B(n_82),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_380),
.B(n_83),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_380),
.B(n_87),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_380),
.B(n_90),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_445),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_450),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_444),
.B(n_91),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_441),
.B(n_93),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_482),
.A2(n_107),
.B(n_111),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_434),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_440),
.A2(n_431),
.B(n_481),
.C(n_459),
.Y(n_506)
);

AO31x2_ASAP7_75t_L g507 ( 
.A1(n_479),
.A2(n_116),
.A3(n_117),
.B(n_119),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_456),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_443),
.A2(n_120),
.B(n_122),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_123),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_428),
.B(n_477),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_481),
.A2(n_125),
.B(n_127),
.C(n_128),
.Y(n_513)
);

OAI22x1_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_453),
.B(n_135),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_426),
.A2(n_137),
.B(n_138),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_429),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_474),
.A2(n_140),
.B(n_141),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_471),
.B(n_142),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_474),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_462),
.B(n_146),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_486),
.B(n_466),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_430),
.B(n_147),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_427),
.A2(n_149),
.B(n_153),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_430),
.B(n_155),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_491),
.A2(n_158),
.B(n_159),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_467),
.Y(n_527)
);

OA21x2_ASAP7_75t_L g528 ( 
.A1(n_449),
.A2(n_160),
.B(n_162),
.Y(n_528)
);

NOR2x1_ASAP7_75t_SL g529 ( 
.A(n_461),
.B(n_164),
.Y(n_529)
);

AOI22x1_ASAP7_75t_SL g530 ( 
.A1(n_452),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_439),
.B(n_170),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_489),
.A2(n_173),
.B(n_183),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_489),
.A2(n_490),
.B(n_451),
.Y(n_533)
);

AO31x2_ASAP7_75t_L g534 ( 
.A1(n_464),
.A2(n_485),
.A3(n_499),
.B(n_473),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_442),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_497),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_475),
.B(n_437),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_436),
.A2(n_432),
.B(n_495),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_469),
.B(n_447),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_446),
.A2(n_480),
.B(n_493),
.Y(n_540)
);

AOI211x1_ASAP7_75t_L g541 ( 
.A1(n_455),
.A2(n_492),
.B(n_483),
.C(n_485),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_498),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_465),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_438),
.B(n_433),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_492),
.A2(n_472),
.B(n_438),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_476),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_460),
.B(n_468),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_472),
.A2(n_499),
.B(n_458),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_454),
.A2(n_463),
.B(n_460),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_448),
.A2(n_457),
.B(n_488),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_487),
.A2(n_478),
.B(n_484),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_496),
.B(n_476),
.Y(n_553)
);

BUFx12f_ASAP7_75t_L g554 ( 
.A(n_465),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_444),
.B(n_363),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_444),
.B(n_337),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_444),
.B(n_337),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_444),
.B(n_370),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_486),
.Y(n_560)
);

AOI221xp5_ASAP7_75t_L g561 ( 
.A1(n_506),
.A2(n_556),
.B1(n_555),
.B2(n_559),
.C(n_541),
.Y(n_561)
);

INVx6_ASAP7_75t_L g562 ( 
.A(n_554),
.Y(n_562)
);

AO21x2_ASAP7_75t_L g563 ( 
.A1(n_545),
.A2(n_549),
.B(n_550),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_533),
.A2(n_540),
.B(n_510),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_522),
.A2(n_523),
.B1(n_560),
.B2(n_527),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_511),
.A2(n_515),
.B(n_519),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_558),
.B(n_517),
.Y(n_567)
);

AO21x2_ASAP7_75t_L g568 ( 
.A1(n_504),
.A2(n_551),
.B(n_552),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_542),
.B(n_502),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_501),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_513),
.A2(n_525),
.B(n_537),
.Y(n_571)
);

A2O1A1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_503),
.A2(n_544),
.B(n_526),
.C(n_508),
.Y(n_572)
);

AOI221xp5_ASAP7_75t_L g573 ( 
.A1(n_514),
.A2(n_557),
.B1(n_512),
.B2(n_520),
.C(n_560),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_538),
.A2(n_509),
.B(n_516),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_560),
.B(n_536),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_535),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_536),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_542),
.B(n_547),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_536),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_546),
.Y(n_580)
);

OAI21x1_ASAP7_75t_SL g581 ( 
.A1(n_529),
.A2(n_518),
.B(n_532),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_542),
.B(n_521),
.Y(n_582)
);

OAI221xp5_ASAP7_75t_L g583 ( 
.A1(n_505),
.A2(n_548),
.B1(n_531),
.B2(n_539),
.C(n_524),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_553),
.A2(n_528),
.B(n_534),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_534),
.Y(n_586)
);

OA21x2_ASAP7_75t_L g587 ( 
.A1(n_534),
.A2(n_507),
.B(n_530),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_507),
.A2(n_538),
.B(n_550),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_543),
.A2(n_440),
.B1(n_434),
.B2(n_523),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_507),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_555),
.B(n_444),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_545),
.A2(n_440),
.B1(n_434),
.B2(n_459),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_555),
.B(n_363),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_555),
.B(n_444),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_560),
.B(n_517),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_506),
.A2(n_545),
.B(n_540),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_543),
.Y(n_597)
);

CKINVDCx8_ASAP7_75t_R g598 ( 
.A(n_560),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_538),
.A2(n_550),
.B(n_443),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_555),
.B(n_363),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_500),
.Y(n_601)
);

OAI221xp5_ASAP7_75t_L g602 ( 
.A1(n_506),
.A2(n_317),
.B1(n_444),
.B2(n_366),
.C(n_440),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_506),
.A2(n_511),
.B1(n_440),
.B2(n_540),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_500),
.Y(n_604)
);

AOI21xp33_ASAP7_75t_L g605 ( 
.A1(n_506),
.A2(n_434),
.B(n_556),
.Y(n_605)
);

OA21x2_ASAP7_75t_L g606 ( 
.A1(n_533),
.A2(n_549),
.B(n_545),
.Y(n_606)
);

O2A1O1Ixp33_ASAP7_75t_L g607 ( 
.A1(n_506),
.A2(n_434),
.B(n_440),
.C(n_459),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_603),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_561),
.B(n_593),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_591),
.B(n_594),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_570),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_575),
.B(n_577),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_604),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_601),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_563),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_563),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_580),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_607),
.A2(n_605),
.B(n_603),
.Y(n_618)
);

INVx11_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_567),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_574),
.A2(n_599),
.B(n_588),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_576),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_575),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_584),
.A2(n_585),
.B(n_581),
.Y(n_624)
);

AOI21x1_ASAP7_75t_L g625 ( 
.A1(n_564),
.A2(n_566),
.B(n_606),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_597),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_577),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_606),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_602),
.B(n_589),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_598),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_568),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_600),
.B(n_571),
.Y(n_633)
);

BUFx2_ASAP7_75t_SL g634 ( 
.A(n_582),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_565),
.A2(n_571),
.B1(n_596),
.B2(n_569),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_568),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_595),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_584),
.A2(n_596),
.B(n_573),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_590),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_579),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_582),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_587),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_583),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_572),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_592),
.B(n_578),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_578),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_592),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_562),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_562),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_613),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_630),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_620),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_612),
.B(n_641),
.Y(n_653)
);

AND2x4_ASAP7_75t_SL g654 ( 
.A(n_612),
.B(n_649),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_609),
.B(n_633),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_646),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_626),
.B(n_610),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_608),
.Y(n_658)
);

AND2x4_ASAP7_75t_SL g659 ( 
.A(n_612),
.B(n_649),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_647),
.B(n_629),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_647),
.B(n_629),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_609),
.B(n_633),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_619),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_630),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_608),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_637),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_611),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_635),
.B(n_645),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_639),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_618),
.B(n_614),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_628),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_645),
.B(n_615),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_614),
.B(n_641),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_646),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_617),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_615),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_617),
.B(n_643),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_616),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_637),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_643),
.B(n_612),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_622),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_638),
.B(n_632),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_619),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_638),
.B(n_632),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_616),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_641),
.B(n_623),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_639),
.B(n_631),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_622),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_642),
.A2(n_631),
.A3(n_636),
.B(n_644),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_636),
.B(n_642),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_640),
.Y(n_691)
);

INVxp67_ASAP7_75t_SL g692 ( 
.A(n_623),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_655),
.B(n_624),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_655),
.B(n_662),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_676),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_676),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_657),
.B(n_634),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_653),
.B(n_627),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_672),
.B(n_668),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_652),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_672),
.B(n_624),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_681),
.B(n_648),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_662),
.B(n_625),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_670),
.B(n_634),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_682),
.B(n_625),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_682),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_678),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_684),
.B(n_621),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_684),
.B(n_621),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_658),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_668),
.B(n_640),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_685),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_667),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_685),
.Y(n_714)
);

AND2x4_ASAP7_75t_SL g715 ( 
.A(n_691),
.B(n_663),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_658),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_663),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_651),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_687),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_687),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_670),
.B(n_640),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_671),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_660),
.B(n_640),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_693),
.B(n_661),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_706),
.B(n_661),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_706),
.B(n_660),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_695),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_693),
.B(n_665),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_700),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_696),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_721),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_710),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_721),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_703),
.B(n_694),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_694),
.B(n_674),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_703),
.B(n_665),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_707),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_708),
.B(n_669),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_718),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_716),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_712),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_709),
.B(n_705),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_723),
.B(n_656),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_699),
.B(n_690),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_718),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_723),
.B(n_669),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_714),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_716),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_709),
.B(n_689),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_729),
.B(n_699),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_730),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_742),
.B(n_705),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_742),
.B(n_701),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_730),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_739),
.B(n_697),
.C(n_704),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_731),
.B(n_701),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_733),
.B(n_724),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_734),
.B(n_719),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_734),
.B(n_711),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_735),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_737),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_724),
.B(n_720),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_743),
.B(n_711),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_738),
.B(n_722),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_737),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_727),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_741),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_744),
.B(n_702),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_746),
.B(n_713),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_741),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_727),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_738),
.B(n_722),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_751),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_754),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_761),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_766),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_765),
.Y(n_777)
);

OAI21xp33_ASAP7_75t_L g778 ( 
.A1(n_768),
.A2(n_755),
.B(n_750),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_760),
.B(n_749),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_767),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_763),
.B(n_745),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_766),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_757),
.A2(n_725),
.B1(n_726),
.B2(n_740),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_768),
.A2(n_651),
.B(n_664),
.C(n_732),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_773),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_779),
.B(n_752),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_776),
.Y(n_787)
);

NAND4xp25_ASAP7_75t_L g788 ( 
.A(n_778),
.B(n_664),
.C(n_688),
.D(n_769),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_784),
.A2(n_726),
.B1(n_725),
.B2(n_758),
.Y(n_789)
);

AOI222xp33_ASAP7_75t_L g790 ( 
.A1(n_781),
.A2(n_736),
.B1(n_753),
.B2(n_759),
.C1(n_680),
.C2(n_728),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_SL g791 ( 
.A(n_783),
.B(n_717),
.Y(n_791)
);

OAI211xp5_ASAP7_75t_SL g792 ( 
.A1(n_789),
.A2(n_779),
.B(n_780),
.C(n_777),
.Y(n_792)
);

OAI211xp5_ASAP7_75t_L g793 ( 
.A1(n_788),
.A2(n_774),
.B(n_775),
.C(n_783),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_791),
.A2(n_756),
.B1(n_762),
.B2(n_744),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_788),
.A2(n_732),
.B(n_748),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_785),
.A2(n_748),
.B(n_770),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_SL g797 ( 
.A1(n_787),
.A2(n_782),
.B(n_648),
.C(n_747),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_797),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_793),
.B(n_796),
.Y(n_799)
);

OAI21xp33_ASAP7_75t_L g800 ( 
.A1(n_792),
.A2(n_790),
.B(n_786),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_795),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_799),
.B(n_794),
.Y(n_802)
);

NAND4xp75_ASAP7_75t_L g803 ( 
.A(n_798),
.B(n_677),
.C(n_686),
.D(n_736),
.Y(n_803)
);

NAND4xp75_ASAP7_75t_L g804 ( 
.A(n_802),
.B(n_801),
.C(n_800),
.D(n_677),
.Y(n_804)
);

INVxp33_ASAP7_75t_SL g805 ( 
.A(n_803),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_803),
.B(n_752),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_804),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_806),
.B(n_759),
.Y(n_808)
);

NOR2x1_ASAP7_75t_L g809 ( 
.A(n_805),
.B(n_683),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_805),
.B(n_771),
.Y(n_810)
);

NAND4xp75_ASAP7_75t_L g811 ( 
.A(n_806),
.B(n_675),
.C(n_680),
.D(n_764),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_809),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_808),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_810),
.Y(n_814)
);

INVxp33_ASAP7_75t_SL g815 ( 
.A(n_807),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_811),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_815),
.A2(n_740),
.B1(n_683),
.B2(n_663),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_813),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_814),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_816),
.B(n_753),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_820),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_818),
.Y(n_822)
);

AOI31xp33_ASAP7_75t_L g823 ( 
.A1(n_819),
.A2(n_812),
.A3(n_692),
.B(n_673),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_817),
.A2(n_683),
.B(n_659),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_818),
.A2(n_659),
.B(n_654),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_821),
.B(n_822),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_823),
.A2(n_654),
.B(n_666),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_825),
.B(n_772),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_824),
.A2(n_666),
.B(n_679),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_826),
.A2(n_679),
.B1(n_717),
.B2(n_698),
.Y(n_830)
);

BUFx2_ASAP7_75t_SL g831 ( 
.A(n_829),
.Y(n_831)
);

OA21x2_ASAP7_75t_L g832 ( 
.A1(n_827),
.A2(n_771),
.B(n_747),
.Y(n_832)
);

OAI31xp33_ASAP7_75t_L g833 ( 
.A1(n_831),
.A2(n_828),
.A3(n_715),
.B(n_650),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_833),
.B(n_830),
.C(n_832),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_834),
.A2(n_715),
.B(n_717),
.Y(n_835)
);


endmodule