module fake_netlist_5_1469_n_2416 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_2416);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2416;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_556;
wire n_2076;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_901;
wire n_553;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_571;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_586;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2009;
wire n_1888;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_2084;
wire n_1781;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2093;
wire n_514;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_507;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_2153;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_1458;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_783;
wire n_555;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_1115;
wire n_703;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_2104;
wire n_518;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_517;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_542;
wire n_1546;
wire n_595;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_257),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_240),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_381),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_392),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_179),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_489),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_249),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_215),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_290),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_135),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_474),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_375),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_224),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_207),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_442),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_462),
.Y(n_521)
);

BUFx5_ASAP7_75t_L g522 ( 
.A(n_469),
.Y(n_522)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_426),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_254),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_16),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_224),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_263),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_302),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_27),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_139),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_58),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_332),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_58),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_488),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_377),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_220),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_308),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_473),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_128),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_22),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_286),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_358),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_223),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_359),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_448),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_186),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_39),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_420),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_346),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_455),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_14),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_263),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_295),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_91),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_464),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_466),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_471),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_485),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_372),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_297),
.Y(n_561)
);

CKINVDCx14_ASAP7_75t_R g562 ( 
.A(n_127),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_219),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_104),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_71),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_212),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_163),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_329),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_271),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_273),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_486),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_87),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_427),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_505),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_199),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_181),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_410),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_176),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_82),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_101),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_294),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_171),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_99),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_167),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_235),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_15),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_85),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_361),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_221),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_498),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_463),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_441),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_44),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_457),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_185),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_432),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_218),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_492),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_499),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_444),
.Y(n_600)
);

BUFx5_ASAP7_75t_L g601 ( 
.A(n_470),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_347),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_38),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_460),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_106),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_317),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_422),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_458),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_231),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_110),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_495),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_480),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_221),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_345),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_119),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_479),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_497),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_468),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_144),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_7),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_214),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_116),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_262),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_219),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_477),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_115),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_114),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_289),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_481),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_11),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_254),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_443),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_253),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_233),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_404),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_360),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_456),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_161),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_214),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_81),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_292),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_218),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_234),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_351),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_171),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_117),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_50),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_96),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_491),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_112),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_13),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_222),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_411),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_155),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_271),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_298),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_437),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_323),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_490),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_209),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_50),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_467),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_235),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_284),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_496),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_298),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_126),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_213),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_54),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_403),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_459),
.Y(n_671)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_494),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_423),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_34),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_144),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_68),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_54),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_179),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_335),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_405),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_461),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_476),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_478),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_48),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_112),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_321),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_160),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_472),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_247),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_452),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_385),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_207),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_264),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_484),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_43),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_333),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_4),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_483),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_216),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_303),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_446),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_465),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_493),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_118),
.Y(n_704)
);

BUFx5_ASAP7_75t_L g705 ( 
.A(n_487),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_59),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_311),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_124),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_200),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_66),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_42),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_74),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_314),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_173),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_136),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_228),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_105),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_337),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_367),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_77),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_228),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_262),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_475),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_386),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_119),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_439),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_387),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_482),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_236),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_374),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_167),
.Y(n_731)
);

CKINVDCx16_ASAP7_75t_R g732 ( 
.A(n_512),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_540),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_639),
.Y(n_734)
);

INVxp33_ASAP7_75t_SL g735 ( 
.A(n_524),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_639),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_652),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_559),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_582),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_652),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_525),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_525),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_525),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_525),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_584),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_529),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_529),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_522),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_731),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_529),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_522),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_529),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_522),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_645),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_645),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_645),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_540),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_579),
.B(n_0),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_645),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_544),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_714),
.Y(n_761)
);

CKINVDCx16_ASAP7_75t_R g762 ( 
.A(n_557),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_714),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_714),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_714),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_716),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_716),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_716),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_709),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_562),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_716),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_562),
.Y(n_772)
);

INVxp33_ASAP7_75t_SL g773 ( 
.A(n_637),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_510),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_521),
.Y(n_775)
);

INVxp33_ASAP7_75t_L g776 ( 
.A(n_578),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_515),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_522),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_527),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_591),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_528),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_506),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_536),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_513),
.Y(n_784)
);

INVxp33_ASAP7_75t_L g785 ( 
.A(n_578),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_539),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_543),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_526),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_526),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_544),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_564),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_518),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_566),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_519),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_570),
.Y(n_795)
);

INVxp33_ASAP7_75t_SL g796 ( 
.A(n_530),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_593),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_533),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_597),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_605),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_522),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_609),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_517),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_623),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_613),
.Y(n_805)
);

INVxp33_ASAP7_75t_SL g806 ( 
.A(n_541),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_631),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_600),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_640),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_641),
.Y(n_810)
);

CKINVDCx16_ASAP7_75t_R g811 ( 
.A(n_607),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_646),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_651),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_661),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_664),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_677),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_678),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_522),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_687),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_692),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_693),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_708),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_725),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_729),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_600),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_613),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_621),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_635),
.Y(n_828)
);

INVxp33_ASAP7_75t_L g829 ( 
.A(n_581),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_635),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_618),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_581),
.B(n_0),
.Y(n_832)
);

INVx5_ASAP7_75t_L g833 ( 
.A(n_803),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_741),
.B(n_679),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_790),
.B(n_573),
.Y(n_835)
);

XNOR2x2_ASAP7_75t_L g836 ( 
.A(n_832),
.B(n_565),
.Y(n_836)
);

OA21x2_ASAP7_75t_L g837 ( 
.A1(n_748),
.A2(n_658),
.B(n_560),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_803),
.Y(n_838)
);

AND2x6_ASAP7_75t_L g839 ( 
.A(n_803),
.B(n_517),
.Y(n_839)
);

OA21x2_ASAP7_75t_L g840 ( 
.A1(n_748),
.A2(n_658),
.B(n_560),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_742),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_743),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_803),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_744),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_746),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_747),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_808),
.B(n_523),
.Y(n_847)
);

BUFx8_ASAP7_75t_SL g848 ( 
.A(n_788),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_760),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_751),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_760),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_750),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_751),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_752),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_773),
.B(n_672),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_738),
.B(n_625),
.Y(n_856)
);

BUFx8_ASAP7_75t_SL g857 ( 
.A(n_788),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_733),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_753),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_754),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_755),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_756),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_759),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_773),
.A2(n_523),
.B1(n_547),
.B2(n_546),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_753),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_778),
.A2(n_698),
.B(n_511),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_778),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_761),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_801),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_763),
.B(n_679),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_775),
.B(n_718),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_764),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_765),
.Y(n_873)
);

CKINVDCx11_ASAP7_75t_R g874 ( 
.A(n_789),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_801),
.A2(n_818),
.B(n_698),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_766),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_767),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_784),
.Y(n_878)
);

OA21x2_ASAP7_75t_L g879 ( 
.A1(n_818),
.A2(n_771),
.B(n_768),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_784),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_774),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_777),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_779),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_832),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_781),
.Y(n_885)
);

OA21x2_ASAP7_75t_L g886 ( 
.A1(n_783),
.A2(n_534),
.B(n_509),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_786),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_796),
.B(n_649),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_735),
.A2(n_624),
.B1(n_630),
.B2(n_621),
.Y(n_889)
);

CKINVDCx11_ASAP7_75t_R g890 ( 
.A(n_789),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_787),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_825),
.B(n_634),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_791),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_793),
.Y(n_894)
);

OA22x2_ASAP7_75t_SL g895 ( 
.A1(n_780),
.A2(n_710),
.B1(n_634),
.B2(n_630),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_795),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_SL g897 ( 
.A(n_762),
.B(n_558),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_879),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_879),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_879),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_888),
.B(n_811),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_879),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_850),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_855),
.B(n_831),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_834),
.B(n_659),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_850),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_850),
.B(n_828),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_838),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_875),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_859),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_849),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_859),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_859),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_875),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_853),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_834),
.B(n_690),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_838),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_849),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_865),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_849),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_853),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_865),
.Y(n_922)
);

AND2x2_ASAP7_75t_SL g923 ( 
.A(n_837),
.B(n_517),
.Y(n_923)
);

OAI21x1_ASAP7_75t_L g924 ( 
.A1(n_866),
.A2(n_550),
.B(n_545),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_865),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_867),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_867),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_836),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_867),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_853),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_853),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_874),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_848),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_869),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_869),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_884),
.B(n_830),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_884),
.B(n_892),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_834),
.B(n_571),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_851),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_869),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_869),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_851),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_837),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_884),
.B(n_785),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_894),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_884),
.B(n_733),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_834),
.B(n_592),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_836),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_884),
.B(n_601),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_837),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_837),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_840),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_838),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_894),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_840),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_840),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_838),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_840),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_866),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_894),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_SL g961 ( 
.A(n_897),
.B(n_558),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_838),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_894),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_894),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_896),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_843),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_896),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_843),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_847),
.B(n_757),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_843),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_896),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_896),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_843),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_847),
.B(n_757),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_843),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_896),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_861),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_860),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_861),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_860),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_861),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_868),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_878),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_860),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_860),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_833),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_886),
.B(n_601),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_944),
.B(n_880),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_930),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_944),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_898),
.B(n_886),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_920),
.Y(n_992)
);

CKINVDCx11_ASAP7_75t_R g993 ( 
.A(n_932),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_983),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_974),
.B(n_732),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_920),
.Y(n_996)
);

AND2x2_ASAP7_75t_SL g997 ( 
.A(n_961),
.B(n_889),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_920),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_937),
.Y(n_999)
);

BUFx4_ASAP7_75t_L g1000 ( 
.A(n_932),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_937),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_942),
.B(n_936),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_936),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_977),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_911),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_905),
.A2(n_864),
.B1(n_835),
.B2(n_871),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_977),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_928),
.B(n_782),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_979),
.Y(n_1009)
);

BUFx4f_ASAP7_75t_L g1010 ( 
.A(n_938),
.Y(n_1010)
);

OR2x6_ASAP7_75t_L g1011 ( 
.A(n_928),
.B(n_858),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_901),
.B(n_796),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_915),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_898),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_979),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_898),
.B(n_886),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_981),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_981),
.Y(n_1018)
);

BUFx8_ASAP7_75t_SL g1019 ( 
.A(n_933),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_905),
.A2(n_856),
.B1(n_806),
.B2(n_772),
.Y(n_1020)
);

OR2x6_ASAP7_75t_L g1021 ( 
.A(n_948),
.B(n_858),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_915),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_982),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_930),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_939),
.B(n_792),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_982),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_918),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_948),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_961),
.B(n_770),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_946),
.B(n_770),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_969),
.B(n_806),
.Y(n_1031)
);

AND2x2_ASAP7_75t_SL g1032 ( 
.A(n_905),
.B(n_889),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_930),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_949),
.A2(n_886),
.B1(n_735),
.B2(n_870),
.Y(n_1034)
);

INVxp33_ASAP7_75t_L g1035 ( 
.A(n_904),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_949),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_899),
.B(n_792),
.Y(n_1037)
);

AND2x6_ASAP7_75t_L g1038 ( 
.A(n_900),
.B(n_517),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_938),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_903),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_938),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_915),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_899),
.B(n_794),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_900),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_905),
.B(n_794),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_900),
.B(n_870),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_903),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_907),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_938),
.A2(n_870),
.B1(n_599),
.B2(n_602),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_907),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_916),
.B(n_772),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_916),
.B(n_798),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_L g1053 ( 
.A(n_943),
.B(n_839),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_903),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_916),
.A2(n_739),
.B1(n_769),
.B2(n_624),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_916),
.B(n_798),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_987),
.A2(n_710),
.B1(n_585),
.B2(n_655),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_947),
.B(n_670),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_906),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_947),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_947),
.A2(n_870),
.B1(n_616),
.B2(n_508),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_899),
.B(n_745),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_906),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_947),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_923),
.B(n_516),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_915),
.B(n_749),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_987),
.B(n_749),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_923),
.B(n_520),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_909),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_909),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_945),
.B(n_882),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_899),
.B(n_805),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_921),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_943),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_902),
.B(n_805),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_923),
.B(n_532),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_914),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_959),
.B(n_734),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_943),
.B(n_892),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_950),
.B(n_604),
.C(n_594),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_945),
.B(n_535),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_914),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_921),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_921),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_959),
.B(n_736),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_921),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_954),
.B(n_537),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_906),
.Y(n_1088)
);

NOR2x1p5_ASAP7_75t_L g1089 ( 
.A(n_959),
.B(n_737),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_934),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_934),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_950),
.B(n_868),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_962),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_924),
.B(n_740),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_934),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_910),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_950),
.A2(n_617),
.B1(n_682),
.B2(n_608),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_934),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_962),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_951),
.B(n_580),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_954),
.B(n_538),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_960),
.B(n_542),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_931),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_SL g1104 ( 
.A1(n_951),
.A2(n_827),
.B1(n_826),
.B2(n_514),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_931),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_935),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_902),
.B(n_826),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_962),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_960),
.B(n_548),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_951),
.B(n_868),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_952),
.B(n_610),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_935),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_952),
.A2(n_955),
.B1(n_958),
.B2(n_956),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_952),
.B(n_885),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_955),
.B(n_885),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_963),
.A2(n_551),
.B1(n_556),
.B2(n_549),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_940),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_968),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_940),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_955),
.B(n_958),
.C(n_956),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_941),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_908),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_L g1123 ( 
.A(n_956),
.B(n_839),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_958),
.B(n_776),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_910),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_902),
.B(n_885),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1103),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_994),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1105),
.Y(n_1129)
);

NOR2xp67_ASAP7_75t_SL g1130 ( 
.A(n_1014),
.B(n_1044),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1095),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_1025),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_990),
.B(n_902),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1120),
.A2(n_924),
.B(n_919),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_990),
.B(n_827),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1074),
.B(n_1113),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1106),
.Y(n_1137)
);

AND2x6_ASAP7_75t_SL g1138 ( 
.A(n_1011),
.B(n_857),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1066),
.B(n_776),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1074),
.B(n_941),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1014),
.B(n_919),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1112),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1117),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1003),
.B(n_1039),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1044),
.B(n_926),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1003),
.B(n_963),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1072),
.B(n_890),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1095),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1124),
.B(n_926),
.Y(n_1149)
);

AND2x6_ASAP7_75t_SL g1150 ( 
.A(n_1011),
.B(n_797),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1048),
.B(n_964),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1050),
.B(n_964),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1075),
.B(n_531),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1036),
.B(n_965),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1107),
.B(n_695),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_999),
.B(n_965),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1001),
.B(n_967),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1031),
.B(n_967),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1041),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_L g1160 ( 
.A(n_1100),
.B(n_971),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1119),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1062),
.B(n_971),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1037),
.B(n_1043),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1013),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1006),
.B(n_1012),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1108),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1010),
.B(n_972),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1111),
.B(n_1079),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1035),
.B(n_995),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1008),
.B(n_882),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_992),
.B(n_887),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1079),
.B(n_972),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_L g1173 ( 
.A(n_1005),
.B(n_1020),
.Y(n_1173)
);

O2A1O1Ixp5_ASAP7_75t_L g1174 ( 
.A1(n_1065),
.A2(n_976),
.B(n_980),
.C(n_978),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1010),
.B(n_976),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_SL g1176 ( 
.A(n_997),
.B(n_629),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1122),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1004),
.B(n_927),
.Y(n_1178)
);

NOR3xp33_ASAP7_75t_L g1179 ( 
.A(n_988),
.B(n_891),
.C(n_887),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1071),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1002),
.B(n_785),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1032),
.B(n_568),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1071),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1019),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1121),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_1027),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1083),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1007),
.B(n_927),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1084),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1090),
.Y(n_1190)
);

NAND2xp33_ASAP7_75t_L g1191 ( 
.A(n_1038),
.B(n_601),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1009),
.B(n_929),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1046),
.A2(n_980),
.B(n_978),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1091),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1015),
.B(n_929),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1017),
.B(n_957),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1098),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1018),
.B(n_957),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1023),
.B(n_957),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1122),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1029),
.B(n_1045),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1056),
.B(n_829),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1028),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1026),
.B(n_1034),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1060),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1114),
.B(n_957),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1099),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1067),
.B(n_829),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1114),
.B(n_966),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1067),
.B(n_552),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1064),
.A2(n_980),
.B1(n_984),
.B2(n_978),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1067),
.A2(n_985),
.B1(n_984),
.B2(n_696),
.Y(n_1212)
);

OAI221xp5_ASAP7_75t_L g1213 ( 
.A1(n_1104),
.A2(n_895),
.B1(n_758),
.B2(n_891),
.C(n_704),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1052),
.B(n_553),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1055),
.B(n_881),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1115),
.B(n_966),
.Y(n_1216)
);

NAND2xp33_ASAP7_75t_L g1217 ( 
.A(n_1038),
.B(n_1122),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1115),
.B(n_966),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1126),
.B(n_966),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1089),
.A2(n_686),
.B1(n_703),
.B2(n_702),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1126),
.B(n_910),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1120),
.B(n_912),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1099),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1030),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1046),
.B(n_912),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1078),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1092),
.B(n_912),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1092),
.B(n_913),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1085),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1068),
.A2(n_985),
.B1(n_984),
.B2(n_713),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1061),
.B(n_574),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1110),
.B(n_913),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1076),
.A2(n_1058),
.B1(n_1102),
.B2(n_1101),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_996),
.B(n_577),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_996),
.B(n_590),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1000),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1118),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_998),
.B(n_596),
.Y(n_1238)
);

O2A1O1Ixp5_ASAP7_75t_L g1239 ( 
.A1(n_1080),
.A2(n_985),
.B(n_970),
.C(n_973),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1057),
.A2(n_507),
.B1(n_555),
.B2(n_554),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_998),
.B(n_598),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1055),
.B(n_561),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1057),
.B(n_606),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1110),
.B(n_991),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1118),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1069),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_991),
.B(n_913),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1070),
.A2(n_724),
.B(n_727),
.C(n_707),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1051),
.B(n_563),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1040),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1016),
.B(n_1077),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1104),
.B(n_881),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1047),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1016),
.B(n_922),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1054),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1059),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1011),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1082),
.Y(n_1258)
);

NOR2xp67_ASAP7_75t_L g1259 ( 
.A(n_1080),
.B(n_883),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1013),
.B(n_922),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1116),
.B(n_611),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1022),
.B(n_567),
.Y(n_1262)
);

AO22x2_ASAP7_75t_L g1263 ( 
.A1(n_1093),
.A2(n_800),
.B1(n_802),
.B2(n_799),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1022),
.B(n_569),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_989),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1021),
.B(n_883),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1024),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1033),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1063),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_993),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1021),
.B(n_1094),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1097),
.B(n_922),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1088),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1096),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1021),
.B(n_804),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1042),
.B(n_1073),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1049),
.A2(n_601),
.B1(n_705),
.B2(n_694),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1042),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1125),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1073),
.B(n_612),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1086),
.B(n_572),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1086),
.B(n_614),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1123),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1038),
.B(n_925),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1038),
.B(n_925),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1053),
.B(n_925),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1094),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1094),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1109),
.B(n_893),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1081),
.B(n_632),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1087),
.A2(n_893),
.B(n_842),
.C(n_844),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1124),
.B(n_968),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_990),
.B(n_636),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1124),
.B(n_968),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1103),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1124),
.B(n_970),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_990),
.B(n_575),
.Y(n_1297)
);

NAND2xp33_ASAP7_75t_L g1298 ( 
.A(n_1124),
.B(n_601),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1103),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1008),
.B(n_807),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1124),
.B(n_970),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_990),
.A2(n_973),
.B1(n_653),
.B2(n_657),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1103),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1027),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1103),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_990),
.B(n_644),
.Y(n_1306)
);

INVxp67_ASAP7_75t_SL g1307 ( 
.A(n_1074),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1124),
.B(n_973),
.Y(n_1308)
);

NOR2xp67_ASAP7_75t_L g1309 ( 
.A(n_1031),
.B(n_809),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1019),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1124),
.B(n_908),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1027),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_SL g1313 ( 
.A(n_1011),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1074),
.B(n_908),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_990),
.B(n_576),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_990),
.A2(n_665),
.B1(n_671),
.B2(n_662),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_990),
.B(n_583),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1074),
.B(n_908),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1095),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_L g1320 ( 
.A(n_1124),
.B(n_601),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1103),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1041),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_990),
.B(n_673),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_SL g1324 ( 
.A(n_997),
.B(n_629),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1019),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1103),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_990),
.B(n_586),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1095),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1246),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1170),
.B(n_893),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1258),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1159),
.B(n_810),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1159),
.B(n_812),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1307),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1250),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1184),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1203),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1139),
.B(n_841),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1127),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1186),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1159),
.B(n_813),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1253),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1322),
.B(n_814),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1132),
.B(n_680),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1242),
.A2(n_642),
.B1(n_663),
.B2(n_619),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1165),
.B(n_681),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1168),
.B(n_854),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1163),
.A2(n_688),
.B1(n_691),
.B2(n_683),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1322),
.B(n_815),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1129),
.Y(n_1350)
);

OR2x2_ASAP7_75t_SL g1351 ( 
.A(n_1275),
.B(n_816),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1153),
.A2(n_701),
.B1(n_719),
.B2(n_700),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1202),
.B(n_731),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1137),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1155),
.A2(n_723),
.B1(n_728),
.B2(n_726),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1164),
.A2(n_917),
.B(n_908),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1176),
.A2(n_705),
.B1(n_588),
.B2(n_694),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1322),
.B(n_817),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1171),
.B(n_819),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1135),
.B(n_587),
.Y(n_1360)
);

OR2x4_ASAP7_75t_L g1361 ( 
.A(n_1147),
.B(n_820),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1310),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1304),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1142),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1325),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1300),
.B(n_821),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1180),
.B(n_730),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1312),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1226),
.B(n_873),
.Y(n_1369)
);

OR2x6_ASAP7_75t_L g1370 ( 
.A(n_1236),
.B(n_822),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1171),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_L g1372 ( 
.A(n_1270),
.Y(n_1372)
);

INVx5_ASAP7_75t_L g1373 ( 
.A(n_1177),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1128),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1271),
.B(n_823),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1229),
.B(n_873),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1143),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1166),
.B(n_824),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1161),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1176),
.A2(n_705),
.B1(n_694),
.B2(n_588),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1136),
.B(n_841),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1255),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1136),
.B(n_842),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1201),
.A2(n_844),
.B1(n_846),
.B2(n_845),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1185),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1295),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1256),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1299),
.Y(n_1388)
);

NAND2xp33_ASAP7_75t_L g1389 ( 
.A(n_1287),
.B(n_705),
.Y(n_1389)
);

AND2x2_ASAP7_75t_SL g1390 ( 
.A(n_1324),
.B(n_588),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1297),
.B(n_845),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1169),
.B(n_589),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1303),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1183),
.B(n_908),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1305),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1321),
.Y(n_1396)
);

AND2x6_ASAP7_75t_SL g1397 ( 
.A(n_1271),
.B(n_846),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1324),
.A2(n_852),
.B1(n_854),
.B2(n_917),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_R g1399 ( 
.A(n_1288),
.B(n_595),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1326),
.Y(n_1400)
);

INVx5_ASAP7_75t_L g1401 ( 
.A(n_1177),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1205),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1266),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1177),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1315),
.B(n_852),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1144),
.B(n_1271),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1200),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1200),
.Y(n_1408)
);

CKINVDCx8_ASAP7_75t_R g1409 ( 
.A(n_1138),
.Y(n_1409)
);

AND2x4_ASAP7_75t_SL g1410 ( 
.A(n_1200),
.B(n_917),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1213),
.A2(n_654),
.B1(n_675),
.B2(n_627),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1317),
.B(n_603),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1182),
.A2(n_917),
.B1(n_975),
.B2(n_953),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1314),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1327),
.B(n_615),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1269),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1181),
.B(n_620),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1309),
.B(n_917),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1164),
.B(n_917),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1173),
.B(n_304),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1257),
.B(n_305),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1224),
.B(n_1214),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1252),
.A2(n_705),
.B1(n_694),
.B2(n_588),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1208),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1274),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_R g1426 ( 
.A(n_1313),
.B(n_622),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1244),
.B(n_626),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1279),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1244),
.A2(n_1133),
.B(n_1311),
.Y(n_1429)
);

NOR2x1_ASAP7_75t_L g1430 ( 
.A(n_1234),
.B(n_1235),
.Y(n_1430)
);

AO22x1_ASAP7_75t_L g1431 ( 
.A1(n_1249),
.A2(n_633),
.B1(n_643),
.B2(n_638),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1314),
.B(n_628),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1262),
.B(n_953),
.Y(n_1433)
);

BUFx5_ASAP7_75t_L g1434 ( 
.A(n_1283),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1264),
.B(n_953),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1318),
.B(n_647),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1178),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1233),
.A2(n_650),
.B(n_656),
.C(n_648),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1215),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1281),
.B(n_953),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1204),
.A2(n_975),
.B1(n_953),
.B2(n_666),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1318),
.B(n_660),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1210),
.B(n_667),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1293),
.B(n_668),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_SL g1445 ( 
.A(n_1179),
.B(n_674),
.C(n_669),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1188),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1306),
.A2(n_953),
.B1(n_975),
.B2(n_705),
.Y(n_1447)
);

OR2x2_ASAP7_75t_SL g1448 ( 
.A(n_1150),
.B(n_676),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1289),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1313),
.Y(n_1450)
);

BUFx8_ASAP7_75t_L g1451 ( 
.A(n_1187),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1263),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1323),
.B(n_684),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1207),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1243),
.A2(n_862),
.B1(n_863),
.B2(n_860),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1131),
.B(n_306),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1192),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1316),
.B(n_1302),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1151),
.B(n_685),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1263),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1263),
.Y(n_1461)
);

NOR2xp67_ASAP7_75t_SL g1462 ( 
.A(n_1276),
.B(n_689),
.Y(n_1462)
);

AO22x1_ASAP7_75t_L g1463 ( 
.A1(n_1240),
.A2(n_699),
.B1(n_706),
.B2(n_697),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1152),
.B(n_711),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1158),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1278),
.B(n_712),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1231),
.A2(n_975),
.B1(n_863),
.B2(n_872),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1160),
.A2(n_975),
.B1(n_863),
.B2(n_872),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_R g1469 ( 
.A(n_1273),
.B(n_715),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1189),
.Y(n_1470)
);

NAND2x1p5_ASAP7_75t_L g1471 ( 
.A(n_1130),
.B(n_975),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1240),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1212),
.B(n_717),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1190),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1220),
.B(n_721),
.C(n_720),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1148),
.B(n_1319),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1328),
.B(n_722),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_R g1478 ( 
.A(n_1265),
.B(n_307),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1223),
.Y(n_1479)
);

INVx5_ASAP7_75t_L g1480 ( 
.A(n_1237),
.Y(n_1480)
);

NOR3xp33_ASAP7_75t_SL g1481 ( 
.A(n_1261),
.B(n_1),
.C(n_2),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1195),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1149),
.B(n_1156),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1251),
.A2(n_862),
.B1(n_872),
.B2(n_863),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1267),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1140),
.B(n_862),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1251),
.A2(n_862),
.B1(n_872),
.B2(n_863),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1268),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1140),
.B(n_862),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1157),
.A2(n_1194),
.B1(n_1197),
.B2(n_1259),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_SL g1491 ( 
.A(n_1248),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1149),
.B(n_872),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1245),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1196),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1141),
.Y(n_1495)
);

INVx5_ASAP7_75t_L g1496 ( 
.A(n_1217),
.Y(n_1496)
);

INVx5_ASAP7_75t_L g1497 ( 
.A(n_1191),
.Y(n_1497)
);

NAND2xp33_ASAP7_75t_L g1498 ( 
.A(n_1154),
.B(n_839),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1141),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1145),
.Y(n_1500)
);

NAND2x1p5_ASAP7_75t_L g1501 ( 
.A(n_1146),
.B(n_876),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1172),
.B(n_876),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1230),
.B(n_1238),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1198),
.Y(n_1504)
);

NAND2x2_ASAP7_75t_L g1505 ( 
.A(n_1199),
.B(n_1),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1241),
.B(n_876),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1145),
.Y(n_1507)
);

BUFx5_ASAP7_75t_L g1508 ( 
.A(n_1239),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1225),
.B(n_876),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1222),
.A2(n_839),
.B1(n_4),
.B2(n_2),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1222),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1292),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1290),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1294),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1296),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1167),
.B(n_3),
.C(n_5),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1301),
.B(n_3),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1308),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1291),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_SL g1520 ( 
.A1(n_1298),
.A2(n_839),
.B(n_877),
.C(n_876),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1175),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1286),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1286),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1211),
.B(n_309),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1260),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1260),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1277),
.A2(n_877),
.B1(n_839),
.B2(n_986),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1225),
.B(n_877),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1162),
.B(n_1227),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1280),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1247),
.Y(n_1531)
);

AND2x6_ASAP7_75t_L g1532 ( 
.A(n_1219),
.B(n_986),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1247),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1134),
.B(n_5),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1254),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1227),
.B(n_877),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1282),
.A2(n_877),
.B1(n_839),
.B2(n_986),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1422),
.B(n_1254),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1449),
.B(n_1272),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1390),
.B(n_1174),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1437),
.B(n_1228),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1446),
.B(n_1228),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_SL g1543 ( 
.A(n_1362),
.B(n_1134),
.Y(n_1543)
);

NAND2xp33_ASAP7_75t_SL g1544 ( 
.A(n_1521),
.B(n_1206),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1449),
.B(n_1221),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1353),
.B(n_1209),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1472),
.B(n_1216),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1371),
.B(n_1218),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1457),
.B(n_1232),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1371),
.B(n_1232),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1403),
.B(n_1284),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_SL g1552 ( 
.A(n_1530),
.B(n_1285),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1366),
.B(n_1193),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1403),
.B(n_1340),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1340),
.B(n_1320),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1424),
.B(n_1439),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_SL g1557 ( 
.A(n_1530),
.B(n_986),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1412),
.B(n_833),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1415),
.B(n_6),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1337),
.B(n_833),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1392),
.B(n_833),
.Y(n_1561)
);

NAND2xp33_ASAP7_75t_SL g1562 ( 
.A(n_1513),
.B(n_986),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1482),
.B(n_6),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1359),
.B(n_7),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1374),
.B(n_833),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1443),
.B(n_833),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1406),
.B(n_310),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1359),
.B(n_8),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1414),
.B(n_1531),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1420),
.B(n_986),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1420),
.B(n_8),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1391),
.B(n_9),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1512),
.B(n_9),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1405),
.B(n_10),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1330),
.B(n_10),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1360),
.B(n_11),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1406),
.B(n_504),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1513),
.B(n_12),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1332),
.B(n_12),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1332),
.B(n_13),
.Y(n_1580)
);

NAND2xp33_ASAP7_75t_SL g1581 ( 
.A(n_1516),
.B(n_1481),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1333),
.B(n_14),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1333),
.B(n_15),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1341),
.B(n_16),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1341),
.B(n_17),
.Y(n_1585)
);

NAND2xp33_ASAP7_75t_SL g1586 ( 
.A(n_1478),
.B(n_1491),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1343),
.B(n_1349),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1343),
.B(n_17),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1349),
.B(n_18),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1358),
.B(n_18),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1358),
.B(n_19),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1417),
.B(n_19),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1363),
.B(n_20),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1465),
.B(n_20),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1515),
.B(n_21),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1411),
.B(n_21),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1368),
.B(n_22),
.Y(n_1597)
);

NAND2xp33_ASAP7_75t_SL g1598 ( 
.A(n_1408),
.B(n_23),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1524),
.B(n_23),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1524),
.B(n_24),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1427),
.B(n_24),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_SL g1602 ( 
.A(n_1408),
.B(n_25),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1466),
.B(n_25),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1514),
.B(n_26),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1469),
.B(n_1453),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1470),
.B(n_26),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1375),
.B(n_503),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1378),
.B(n_27),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1518),
.B(n_28),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1474),
.B(n_28),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1375),
.B(n_312),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1373),
.B(n_29),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1373),
.B(n_29),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1373),
.B(n_30),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1401),
.B(n_30),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1401),
.B(n_31),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1401),
.B(n_31),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1450),
.B(n_32),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1459),
.B(n_1464),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1329),
.B(n_32),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1460),
.B(n_33),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1338),
.B(n_33),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1331),
.B(n_34),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1339),
.B(n_35),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1421),
.B(n_1350),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1452),
.B(n_35),
.Y(n_1626)
);

NAND2xp33_ASAP7_75t_SL g1627 ( 
.A(n_1461),
.B(n_36),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1354),
.B(n_36),
.Y(n_1628)
);

NAND2xp33_ASAP7_75t_SL g1629 ( 
.A(n_1364),
.B(n_37),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1377),
.B(n_37),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1533),
.B(n_38),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1535),
.B(n_39),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1379),
.B(n_40),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1444),
.B(n_40),
.Y(n_1635)
);

NAND2xp33_ASAP7_75t_SL g1636 ( 
.A(n_1388),
.B(n_41),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1393),
.B(n_41),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1395),
.B(n_42),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1396),
.B(n_43),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1400),
.B(n_44),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1399),
.B(n_1347),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1402),
.B(n_45),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1458),
.B(n_45),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1456),
.B(n_46),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1456),
.B(n_46),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1495),
.B(n_47),
.Y(n_1646)
);

NAND2xp33_ASAP7_75t_SL g1647 ( 
.A(n_1404),
.B(n_47),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1499),
.B(n_48),
.Y(n_1648)
);

NAND2xp33_ASAP7_75t_SL g1649 ( 
.A(n_1462),
.B(n_49),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1500),
.B(n_49),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1451),
.B(n_51),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1480),
.B(n_51),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1480),
.B(n_52),
.Y(n_1653)
);

NAND2xp33_ASAP7_75t_SL g1654 ( 
.A(n_1365),
.B(n_52),
.Y(n_1654)
);

NAND2xp33_ASAP7_75t_SL g1655 ( 
.A(n_1421),
.B(n_1426),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_SL g1656 ( 
.A(n_1507),
.B(n_1529),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1480),
.B(n_53),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1352),
.B(n_53),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1355),
.B(n_55),
.Y(n_1659)
);

NAND2xp33_ASAP7_75t_SL g1660 ( 
.A(n_1485),
.B(n_55),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1432),
.B(n_1436),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1442),
.B(n_56),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1369),
.B(n_56),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1376),
.B(n_57),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1334),
.B(n_57),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1488),
.B(n_59),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1517),
.B(n_60),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1511),
.B(n_60),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1463),
.B(n_61),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1430),
.B(n_61),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1525),
.B(n_62),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1526),
.B(n_1483),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1534),
.B(n_1346),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1438),
.B(n_62),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1434),
.B(n_63),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1434),
.B(n_63),
.Y(n_1676)
);

XNOR2xp5_ASAP7_75t_L g1677 ( 
.A(n_1448),
.B(n_313),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1434),
.B(n_64),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1434),
.B(n_64),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1335),
.B(n_1342),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1382),
.B(n_65),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1387),
.B(n_65),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1416),
.B(n_66),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1425),
.B(n_67),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1428),
.B(n_67),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1407),
.B(n_315),
.Y(n_1686)
);

NAND2xp33_ASAP7_75t_SL g1687 ( 
.A(n_1344),
.B(n_1367),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1345),
.B(n_68),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1496),
.B(n_69),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1496),
.B(n_69),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1496),
.B(n_70),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1454),
.B(n_502),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1431),
.B(n_70),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1490),
.B(n_71),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1479),
.B(n_72),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1504),
.B(n_72),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_SL g1697 ( 
.A(n_1477),
.B(n_73),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1494),
.B(n_73),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1348),
.B(n_74),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1493),
.B(n_75),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1370),
.B(n_75),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1351),
.B(n_76),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1522),
.B(n_76),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1398),
.B(n_77),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_SL g1705 ( 
.A(n_1372),
.B(n_316),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1475),
.B(n_78),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1336),
.B(n_500),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1476),
.B(n_1523),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1384),
.B(n_78),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1503),
.B(n_79),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1370),
.B(n_79),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1410),
.B(n_318),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1429),
.B(n_80),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1473),
.B(n_80),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1381),
.B(n_81),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1497),
.B(n_1519),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1497),
.B(n_82),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1497),
.B(n_83),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1357),
.B(n_83),
.Y(n_1719)
);

NAND2xp33_ASAP7_75t_SL g1720 ( 
.A(n_1380),
.B(n_84),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1383),
.B(n_84),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1510),
.B(n_85),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1423),
.B(n_86),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1433),
.B(n_86),
.Y(n_1724)
);

NAND2xp33_ASAP7_75t_SL g1725 ( 
.A(n_1506),
.B(n_87),
.Y(n_1725)
);

NAND2xp33_ASAP7_75t_SL g1726 ( 
.A(n_1418),
.B(n_88),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1435),
.B(n_88),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1440),
.B(n_89),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1492),
.B(n_89),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1413),
.B(n_90),
.Y(n_1730)
);

NAND2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1394),
.B(n_90),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1508),
.B(n_319),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1486),
.B(n_91),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1658),
.A2(n_1445),
.B1(n_1505),
.B2(n_1389),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1554),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1641),
.B(n_1501),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1634),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1586),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1538),
.B(n_1549),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1599),
.A2(n_1361),
.B1(n_1471),
.B2(n_1489),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1672),
.Y(n_1741)
);

OR2x6_ASAP7_75t_L g1742 ( 
.A(n_1716),
.B(n_1419),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1659),
.A2(n_1508),
.B1(n_1441),
.B2(n_1498),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1625),
.Y(n_1744)
);

AND2x4_ASAP7_75t_L g1745 ( 
.A(n_1625),
.B(n_1447),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1668),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1541),
.B(n_1509),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1569),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1655),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1605),
.B(n_1397),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1680),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1622),
.B(n_1409),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1587),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1556),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1541),
.B(n_1528),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1608),
.B(n_1455),
.Y(n_1756)
);

INVxp33_ASAP7_75t_L g1757 ( 
.A(n_1547),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1707),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1546),
.B(n_92),
.Y(n_1759)
);

AND3x1_ASAP7_75t_SL g1760 ( 
.A(n_1688),
.B(n_92),
.C(n_93),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1619),
.B(n_1502),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1553),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1544),
.B(n_1508),
.Y(n_1763)
);

BUFx12f_ASAP7_75t_L g1764 ( 
.A(n_1707),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1559),
.B(n_1536),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1545),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1708),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1600),
.A2(n_1468),
.B1(n_1356),
.B2(n_1527),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1542),
.B(n_1508),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1539),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1703),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1635),
.B(n_1621),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1631),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1582),
.B(n_93),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1646),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1567),
.B(n_1467),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1542),
.B(n_1532),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1571),
.B(n_320),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1567),
.B(n_1537),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1563),
.Y(n_1780)
);

AND3x1_ASAP7_75t_SL g1781 ( 
.A(n_1618),
.B(n_94),
.C(n_95),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_R g1782 ( 
.A(n_1577),
.B(n_1607),
.Y(n_1782)
);

AND3x1_ASAP7_75t_SL g1783 ( 
.A(n_1581),
.B(n_94),
.C(n_95),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1550),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1661),
.B(n_1715),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1559),
.A2(n_1532),
.B1(n_1487),
.B2(n_1484),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1686),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1577),
.B(n_1686),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1548),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1607),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1721),
.B(n_1532),
.Y(n_1791)
);

BUFx12f_ASAP7_75t_L g1792 ( 
.A(n_1611),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1564),
.B(n_96),
.Y(n_1793)
);

BUFx2_ASAP7_75t_L g1794 ( 
.A(n_1611),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1712),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1568),
.B(n_97),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1573),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1682),
.Y(n_1798)
);

A2O1A1Ixp33_ASAP7_75t_L g1799 ( 
.A1(n_1673),
.A2(n_1520),
.B(n_99),
.C(n_97),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1699),
.A2(n_101),
.B1(n_98),
.B2(n_100),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1669),
.B(n_98),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1656),
.B(n_100),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1595),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1693),
.B(n_1702),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1596),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_1712),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1665),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1702),
.B(n_1667),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1692),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1604),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1632),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1609),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1692),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1733),
.Y(n_1814)
);

O2A1O1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1576),
.A2(n_105),
.B(n_102),
.C(n_103),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1572),
.B(n_106),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1729),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1551),
.Y(n_1818)
);

BUFx2_ASAP7_75t_R g1819 ( 
.A(n_1722),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1701),
.B(n_107),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1671),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1644),
.B(n_322),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1648),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1574),
.B(n_107),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1650),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1645),
.B(n_108),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1695),
.Y(n_1827)
);

INVx4_ASAP7_75t_L g1828 ( 
.A(n_1711),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1713),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1662),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1543),
.B(n_108),
.Y(n_1831)
);

AND2x2_ASAP7_75t_SL g1832 ( 
.A(n_1705),
.B(n_109),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1710),
.B(n_109),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1687),
.B(n_110),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1555),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1709),
.A2(n_114),
.B1(n_111),
.B2(n_113),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1565),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1643),
.B(n_111),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_R g1839 ( 
.A(n_1552),
.B(n_324),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1696),
.B(n_113),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1681),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1675),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1697),
.B(n_115),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1677),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1676),
.Y(n_1845)
);

BUFx8_ASAP7_75t_L g1846 ( 
.A(n_1651),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1654),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1678),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1570),
.B(n_116),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1540),
.B(n_117),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1540),
.B(n_1694),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1670),
.B(n_1598),
.Y(n_1852)
);

CKINVDCx16_ASAP7_75t_R g1853 ( 
.A(n_1602),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1730),
.B(n_118),
.Y(n_1854)
);

AOI22x1_ASAP7_75t_L g1855 ( 
.A1(n_1649),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1663),
.B(n_1664),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1592),
.B(n_325),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1679),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1601),
.B(n_120),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1683),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1575),
.B(n_121),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1562),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1724),
.B(n_122),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1652),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1727),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1603),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1714),
.A2(n_126),
.B1(n_123),
.B2(n_125),
.Y(n_1867)
);

BUFx4f_ASAP7_75t_SL g1868 ( 
.A(n_1578),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1593),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1732),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1728),
.B(n_127),
.Y(n_1871)
);

BUFx4f_ASAP7_75t_L g1872 ( 
.A(n_1557),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1704),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1732),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1561),
.B(n_129),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1620),
.B(n_130),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1698),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1597),
.Y(n_1878)
);

INVx4_ASAP7_75t_L g1879 ( 
.A(n_1626),
.Y(n_1879)
);

BUFx6f_ASAP7_75t_L g1880 ( 
.A(n_1653),
.Y(n_1880)
);

CKINVDCx16_ASAP7_75t_R g1881 ( 
.A(n_1647),
.Y(n_1881)
);

BUFx3_ASAP7_75t_L g1882 ( 
.A(n_1579),
.Y(n_1882)
);

INVxp67_ASAP7_75t_SL g1883 ( 
.A(n_1560),
.Y(n_1883)
);

BUFx12f_ASAP7_75t_L g1884 ( 
.A(n_1580),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1674),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1623),
.B(n_131),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1657),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1566),
.B(n_132),
.Y(n_1888)
);

INVx4_ASAP7_75t_SL g1889 ( 
.A(n_1629),
.Y(n_1889)
);

BUFx3_ASAP7_75t_L g1890 ( 
.A(n_1583),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1584),
.B(n_326),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1684),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1624),
.B(n_133),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1685),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1585),
.B(n_327),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1723),
.B(n_134),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1558),
.B(n_134),
.Y(n_1897)
);

INVx8_ASAP7_75t_L g1898 ( 
.A(n_1764),
.Y(n_1898)
);

AOI22x1_ASAP7_75t_L g1899 ( 
.A1(n_1879),
.A2(n_1630),
.B1(n_1636),
.B2(n_1660),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1811),
.Y(n_1900)
);

BUFx12f_ASAP7_75t_L g1901 ( 
.A(n_1738),
.Y(n_1901)
);

CKINVDCx16_ASAP7_75t_R g1902 ( 
.A(n_1782),
.Y(n_1902)
);

OAI21x1_ASAP7_75t_L g1903 ( 
.A1(n_1747),
.A2(n_1706),
.B(n_1700),
.Y(n_1903)
);

BUFx8_ASAP7_75t_L g1904 ( 
.A(n_1792),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1748),
.Y(n_1905)
);

INVx5_ASAP7_75t_L g1906 ( 
.A(n_1742),
.Y(n_1906)
);

AOI22x1_ASAP7_75t_L g1907 ( 
.A1(n_1879),
.A2(n_1627),
.B1(n_1725),
.B2(n_1726),
.Y(n_1907)
);

NAND2x1p5_ASAP7_75t_L g1908 ( 
.A(n_1872),
.B(n_1717),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1762),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1741),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1846),
.Y(n_1911)
);

OAI21x1_ASAP7_75t_L g1912 ( 
.A1(n_1747),
.A2(n_1718),
.B(n_1690),
.Y(n_1912)
);

AO21x2_ASAP7_75t_L g1913 ( 
.A1(n_1763),
.A2(n_1666),
.B(n_1633),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1788),
.B(n_1689),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1758),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1769),
.Y(n_1916)
);

AO21x2_ASAP7_75t_L g1917 ( 
.A1(n_1799),
.A2(n_1637),
.B(n_1628),
.Y(n_1917)
);

BUFx4f_ASAP7_75t_L g1918 ( 
.A(n_1790),
.Y(n_1918)
);

BUFx10_ASAP7_75t_L g1919 ( 
.A(n_1750),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1788),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1757),
.B(n_1811),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1809),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1790),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1846),
.Y(n_1924)
);

NOR2x1_ASAP7_75t_R g1925 ( 
.A(n_1844),
.B(n_1588),
.Y(n_1925)
);

OAI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1765),
.A2(n_1719),
.B(n_1720),
.Y(n_1926)
);

BUFx3_ASAP7_75t_L g1927 ( 
.A(n_1790),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1806),
.Y(n_1928)
);

OAI21x1_ASAP7_75t_L g1929 ( 
.A1(n_1755),
.A2(n_1691),
.B(n_1639),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1806),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1751),
.Y(n_1931)
);

BUFx2_ASAP7_75t_R g1932 ( 
.A(n_1847),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1737),
.Y(n_1933)
);

BUFx4f_ASAP7_75t_L g1934 ( 
.A(n_1806),
.Y(n_1934)
);

OR2x6_ASAP7_75t_L g1935 ( 
.A(n_1870),
.B(n_1612),
.Y(n_1935)
);

OAI21x1_ASAP7_75t_SL g1936 ( 
.A1(n_1802),
.A2(n_1731),
.B(n_1640),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1807),
.B(n_1594),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1769),
.Y(n_1938)
);

BUFx3_ASAP7_75t_L g1939 ( 
.A(n_1794),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1767),
.Y(n_1940)
);

INVx6_ASAP7_75t_L g1941 ( 
.A(n_1809),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1766),
.Y(n_1942)
);

OAI21x1_ASAP7_75t_SL g1943 ( 
.A1(n_1802),
.A2(n_1642),
.B(n_1638),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1798),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1739),
.B(n_1606),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1808),
.B(n_1613),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1770),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1755),
.A2(n_1615),
.B(n_1614),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1874),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1784),
.Y(n_1950)
);

AO21x2_ASAP7_75t_L g1951 ( 
.A1(n_1850),
.A2(n_1617),
.B(n_1616),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1739),
.Y(n_1952)
);

BUFx2_ASAP7_75t_SL g1953 ( 
.A(n_1749),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1818),
.Y(n_1954)
);

OAI21x1_ASAP7_75t_L g1955 ( 
.A1(n_1777),
.A2(n_1610),
.B(n_1590),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1850),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1851),
.A2(n_1591),
.B(n_1589),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1832),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_1958)
);

BUFx2_ASAP7_75t_SL g1959 ( 
.A(n_1828),
.Y(n_1959)
);

BUFx2_ASAP7_75t_L g1960 ( 
.A(n_1744),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1777),
.A2(n_330),
.B(n_328),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1743),
.A2(n_334),
.B(n_331),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_1828),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1746),
.B(n_137),
.Y(n_1964)
);

AOI22x1_ASAP7_75t_L g1965 ( 
.A1(n_1881),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_1965)
);

CKINVDCx6p67_ASAP7_75t_R g1966 ( 
.A(n_1884),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_1837),
.Y(n_1967)
);

CKINVDCx20_ASAP7_75t_R g1968 ( 
.A(n_1853),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1789),
.Y(n_1969)
);

INVxp67_ASAP7_75t_SL g1970 ( 
.A(n_1851),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1791),
.A2(n_338),
.B(n_336),
.Y(n_1971)
);

BUFx12f_ASAP7_75t_L g1972 ( 
.A(n_1878),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1835),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1780),
.B(n_1797),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1771),
.B(n_138),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1768),
.A2(n_340),
.B(n_339),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1787),
.Y(n_1977)
);

NAND2x1p5_ASAP7_75t_L g1978 ( 
.A(n_1872),
.B(n_341),
.Y(n_1978)
);

OAI21x1_ASAP7_75t_L g1979 ( 
.A1(n_1791),
.A2(n_343),
.B(n_342),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_L g1980 ( 
.A1(n_1761),
.A2(n_1768),
.B(n_1786),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1809),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1814),
.B(n_140),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1803),
.B(n_141),
.Y(n_1983)
);

NAND2x1_ASAP7_75t_L g1984 ( 
.A(n_1742),
.B(n_344),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1773),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1810),
.B(n_141),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1775),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1740),
.A2(n_349),
.B(n_348),
.Y(n_1988)
);

OA21x2_ASAP7_75t_L g1989 ( 
.A1(n_1785),
.A2(n_142),
.B(n_143),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1795),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1735),
.Y(n_1991)
);

INVx5_ASAP7_75t_L g1992 ( 
.A(n_1742),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1813),
.B(n_350),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1829),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1869),
.Y(n_1995)
);

BUFx2_ASAP7_75t_SL g1996 ( 
.A(n_1772),
.Y(n_1996)
);

OAI21x1_ASAP7_75t_L g1997 ( 
.A1(n_1740),
.A2(n_353),
.B(n_352),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1812),
.Y(n_1998)
);

INVx4_ASAP7_75t_L g1999 ( 
.A(n_1795),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1753),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1785),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1804),
.B(n_354),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1910),
.Y(n_2003)
);

BUFx8_ASAP7_75t_L g2004 ( 
.A(n_1901),
.Y(n_2004)
);

AOI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1958),
.A2(n_1834),
.B1(n_1852),
.B2(n_1843),
.Y(n_2005)
);

BUFx2_ASAP7_75t_L g2006 ( 
.A(n_1963),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1952),
.B(n_1817),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1958),
.A2(n_1855),
.B1(n_1873),
.B2(n_1836),
.Y(n_2008)
);

AOI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1965),
.A2(n_1873),
.B1(n_1800),
.B2(n_1805),
.Y(n_2009)
);

BUFx12f_ASAP7_75t_L g2010 ( 
.A(n_1904),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1904),
.Y(n_2011)
);

INVx6_ASAP7_75t_L g2012 ( 
.A(n_1928),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1905),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_SL g2014 ( 
.A1(n_1902),
.A2(n_1831),
.B1(n_1868),
.B2(n_1801),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1946),
.A2(n_1778),
.B1(n_1822),
.B2(n_1857),
.Y(n_2015)
);

OAI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1983),
.A2(n_1831),
.B1(n_1866),
.B2(n_1867),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1983),
.A2(n_1859),
.B1(n_1885),
.B2(n_1822),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1986),
.A2(n_1854),
.B1(n_1833),
.B2(n_1838),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1954),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1908),
.A2(n_1819),
.B1(n_1734),
.B2(n_1882),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1996),
.B(n_1820),
.Y(n_2021)
);

BUFx12f_ASAP7_75t_L g2022 ( 
.A(n_1911),
.Y(n_2022)
);

AOI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_1986),
.A2(n_1840),
.B1(n_1833),
.B2(n_1838),
.Y(n_2023)
);

INVx1_ASAP7_75t_SL g2024 ( 
.A(n_1900),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1952),
.B(n_1759),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1899),
.A2(n_1861),
.B1(n_1856),
.B2(n_1824),
.Y(n_2026)
);

CKINVDCx6p67_ASAP7_75t_R g2027 ( 
.A(n_1972),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1946),
.A2(n_1830),
.B1(n_1854),
.B2(n_1816),
.Y(n_2028)
);

CKINVDCx6p67_ASAP7_75t_R g2029 ( 
.A(n_1966),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1926),
.A2(n_1876),
.B1(n_1893),
.B2(n_1886),
.Y(n_2030)
);

AOI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1907),
.A2(n_1917),
.B1(n_1745),
.B2(n_1936),
.Y(n_2031)
);

AOI22xp33_ASAP7_75t_L g2032 ( 
.A1(n_1917),
.A2(n_1745),
.B1(n_1890),
.B2(n_1776),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1954),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1916),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1938),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_1914),
.A2(n_1776),
.B1(n_1895),
.B2(n_1891),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1970),
.Y(n_2037)
);

BUFx3_ASAP7_75t_L g2038 ( 
.A(n_1944),
.Y(n_2038)
);

INVx1_ASAP7_75t_SL g2039 ( 
.A(n_1900),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1909),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_SL g2041 ( 
.A1(n_1989),
.A2(n_1839),
.B1(n_1826),
.B2(n_1896),
.Y(n_2041)
);

CKINVDCx6p67_ASAP7_75t_R g2042 ( 
.A(n_1898),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1970),
.Y(n_2043)
);

INVx1_ASAP7_75t_SL g2044 ( 
.A(n_1991),
.Y(n_2044)
);

CKINVDCx11_ASAP7_75t_R g2045 ( 
.A(n_1968),
.Y(n_2045)
);

INVx1_ASAP7_75t_SL g2046 ( 
.A(n_1953),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1949),
.Y(n_2047)
);

INVx6_ASAP7_75t_L g2048 ( 
.A(n_1928),
.Y(n_2048)
);

OAI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1937),
.A2(n_1896),
.B1(n_1871),
.B2(n_1863),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1985),
.Y(n_2050)
);

CKINVDCx11_ASAP7_75t_R g2051 ( 
.A(n_1968),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1926),
.A2(n_1871),
.B1(n_1863),
.B2(n_1877),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1987),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1995),
.Y(n_2054)
);

INVx6_ASAP7_75t_L g2055 ( 
.A(n_1928),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_1942),
.B(n_1837),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_SL g2057 ( 
.A1(n_1989),
.A2(n_1864),
.B1(n_1887),
.B2(n_1880),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1908),
.A2(n_1880),
.B1(n_1887),
.B2(n_1864),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_SL g2059 ( 
.A1(n_1943),
.A2(n_1864),
.B1(n_1887),
.B2(n_1880),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1921),
.A2(n_1865),
.B1(n_1823),
.B2(n_1825),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1998),
.Y(n_2061)
);

BUFx3_ASAP7_75t_L g2062 ( 
.A(n_1898),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1898),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_2041),
.B(n_1906),
.Y(n_2064)
);

A2O1A1Ixp33_ASAP7_75t_L g2065 ( 
.A1(n_2008),
.A2(n_1976),
.B(n_1815),
.C(n_1957),
.Y(n_2065)
);

BUFx2_ASAP7_75t_L g2066 ( 
.A(n_2006),
.Y(n_2066)
);

OAI211xp5_ASAP7_75t_L g2067 ( 
.A1(n_2008),
.A2(n_1957),
.B(n_1976),
.C(n_1982),
.Y(n_2067)
);

OA21x2_ASAP7_75t_L g2068 ( 
.A1(n_2031),
.A2(n_1980),
.B(n_1988),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2016),
.A2(n_1736),
.B(n_1862),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2019),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2033),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2037),
.B(n_2000),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_2024),
.B(n_1956),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2039),
.B(n_1921),
.Y(n_2074)
);

AOI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_2016),
.A2(n_1992),
.B(n_1906),
.Y(n_2075)
);

OAI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_2015),
.A2(n_1997),
.B(n_1903),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_2044),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_2032),
.A2(n_1979),
.B(n_1971),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_2018),
.A2(n_1992),
.B(n_1906),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_2009),
.A2(n_2005),
.B1(n_2017),
.B2(n_2014),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2003),
.Y(n_2081)
);

AOI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_2018),
.A2(n_1992),
.B(n_1906),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_2038),
.Y(n_2083)
);

AOI221xp5_ASAP7_75t_L g2084 ( 
.A1(n_2049),
.A2(n_1974),
.B1(n_1982),
.B2(n_1975),
.C(n_1964),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2047),
.Y(n_2085)
);

AOI221xp5_ASAP7_75t_L g2086 ( 
.A1(n_2049),
.A2(n_1974),
.B1(n_1975),
.B2(n_1964),
.C(n_2000),
.Y(n_2086)
);

A2O1A1Ixp33_ASAP7_75t_L g2087 ( 
.A1(n_2009),
.A2(n_1779),
.B(n_1962),
.C(n_1912),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2021),
.B(n_1919),
.Y(n_2088)
);

AO21x2_ASAP7_75t_L g2089 ( 
.A1(n_2043),
.A2(n_1949),
.B(n_1888),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2025),
.B(n_1994),
.Y(n_2090)
);

BUFx8_ASAP7_75t_SL g2091 ( 
.A(n_2010),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2013),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2050),
.Y(n_2093)
);

AOI221x1_ASAP7_75t_SL g2094 ( 
.A1(n_2020),
.A2(n_1945),
.B1(n_2001),
.B2(n_1947),
.C(n_1821),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_2053),
.B(n_1992),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_2034),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_2060),
.B(n_1967),
.Y(n_2097)
);

AND2x2_ASAP7_75t_SL g2098 ( 
.A(n_2052),
.B(n_1934),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2061),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2090),
.B(n_2035),
.Y(n_2100)
);

AOI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_2080),
.A2(n_2014),
.B1(n_2041),
.B2(n_2017),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_L g2102 ( 
.A1(n_2064),
.A2(n_2026),
.B1(n_2036),
.B2(n_2059),
.Y(n_2102)
);

AOI211xp5_ASAP7_75t_L g2103 ( 
.A1(n_2064),
.A2(n_2067),
.B(n_2086),
.C(n_2065),
.Y(n_2103)
);

OAI211xp5_ASAP7_75t_SL g2104 ( 
.A1(n_2084),
.A2(n_2023),
.B(n_2065),
.C(n_2028),
.Y(n_2104)
);

BUFx6f_ASAP7_75t_L g2105 ( 
.A(n_2091),
.Y(n_2105)
);

AOI221x1_ASAP7_75t_L g2106 ( 
.A1(n_2079),
.A2(n_2058),
.B1(n_2007),
.B2(n_2056),
.C(n_1973),
.Y(n_2106)
);

OAI221xp5_ASAP7_75t_L g2107 ( 
.A1(n_2094),
.A2(n_2023),
.B1(n_2026),
.B2(n_2052),
.C(n_2059),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_2095),
.B(n_2066),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_2077),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2073),
.B(n_2040),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_2095),
.Y(n_2111)
);

AOI222xp33_ASAP7_75t_L g2112 ( 
.A1(n_2098),
.A2(n_2030),
.B1(n_2028),
.B2(n_2076),
.C1(n_1925),
.C2(n_1889),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2070),
.B(n_2056),
.Y(n_2113)
);

OAI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_2075),
.A2(n_2030),
.B1(n_2057),
.B2(n_2046),
.C(n_1978),
.Y(n_2114)
);

OAI21x1_ASAP7_75t_L g2115 ( 
.A1(n_2082),
.A2(n_1961),
.B(n_1929),
.Y(n_2115)
);

AOI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_2098),
.A2(n_1914),
.B1(n_1919),
.B2(n_1913),
.Y(n_2116)
);

OAI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_2069),
.A2(n_2057),
.B1(n_1935),
.B2(n_1978),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_2071),
.B(n_2062),
.Y(n_2118)
);

AOI221xp5_ASAP7_75t_L g2119 ( 
.A1(n_2074),
.A2(n_1754),
.B1(n_1796),
.B2(n_1793),
.C(n_1774),
.Y(n_2119)
);

NAND3xp33_ASAP7_75t_L g2120 ( 
.A(n_2087),
.B(n_1994),
.C(n_1945),
.Y(n_2120)
);

OAI221xp5_ASAP7_75t_L g2121 ( 
.A1(n_2103),
.A2(n_2087),
.B1(n_2097),
.B2(n_2083),
.C(n_2011),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_2105),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2108),
.B(n_2088),
.Y(n_2123)
);

AO31x2_ASAP7_75t_L g2124 ( 
.A1(n_2106),
.A2(n_2097),
.A3(n_2085),
.B(n_2093),
.Y(n_2124)
);

BUFx2_ASAP7_75t_L g2125 ( 
.A(n_2111),
.Y(n_2125)
);

INVxp67_ASAP7_75t_SL g2126 ( 
.A(n_2111),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2100),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2108),
.B(n_2096),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2113),
.Y(n_2129)
);

AOI22xp33_ASAP7_75t_L g2130 ( 
.A1(n_2104),
.A2(n_2068),
.B1(n_2078),
.B2(n_1913),
.Y(n_2130)
);

INVxp67_ASAP7_75t_L g2131 ( 
.A(n_2121),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2127),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2127),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_2122),
.Y(n_2134)
);

BUFx3_ASAP7_75t_L g2135 ( 
.A(n_2122),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_2130),
.A2(n_2101),
.B(n_2107),
.Y(n_2136)
);

INVx5_ASAP7_75t_L g2137 ( 
.A(n_2134),
.Y(n_2137)
);

AOI33xp33_ASAP7_75t_L g2138 ( 
.A1(n_2133),
.A2(n_2132),
.A3(n_2102),
.B1(n_2119),
.B2(n_2116),
.B3(n_2136),
.Y(n_2138)
);

INVx5_ASAP7_75t_L g2139 ( 
.A(n_2134),
.Y(n_2139)
);

OAI221xp5_ASAP7_75t_L g2140 ( 
.A1(n_2131),
.A2(n_2112),
.B1(n_2120),
.B2(n_2117),
.C(n_2114),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2135),
.B(n_2129),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_2132),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2135),
.Y(n_2143)
);

AOI21x1_ASAP7_75t_L g2144 ( 
.A1(n_2134),
.A2(n_2125),
.B(n_2128),
.Y(n_2144)
);

INVxp67_ASAP7_75t_SL g2145 ( 
.A(n_2134),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2141),
.B(n_2125),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_2137),
.B(n_2122),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2142),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2143),
.B(n_2129),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2145),
.B(n_2124),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2142),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2145),
.B(n_2122),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2137),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2137),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2137),
.B(n_2128),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2139),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2148),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_2147),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2151),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2152),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2154),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2146),
.B(n_2122),
.Y(n_2162)
);

NAND4xp75_ASAP7_75t_SL g2163 ( 
.A(n_2155),
.B(n_2144),
.C(n_2138),
.D(n_2068),
.Y(n_2163)
);

NAND3xp33_ASAP7_75t_L g2164 ( 
.A(n_2153),
.B(n_2140),
.C(n_2139),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2160),
.B(n_2149),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2162),
.B(n_2149),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2158),
.B(n_2146),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2161),
.B(n_2156),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2167),
.Y(n_2169)
);

AOI22xp33_ASAP7_75t_L g2170 ( 
.A1(n_2166),
.A2(n_2164),
.B1(n_2155),
.B2(n_2159),
.Y(n_2170)
);

OAI21xp33_ASAP7_75t_L g2171 ( 
.A1(n_2165),
.A2(n_2164),
.B(n_2157),
.Y(n_2171)
);

NAND4xp75_ASAP7_75t_L g2172 ( 
.A(n_2168),
.B(n_2154),
.C(n_2163),
.D(n_2147),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2169),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2170),
.B(n_2147),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2171),
.B(n_2105),
.Y(n_2175)
);

A2O1A1Ixp33_ASAP7_75t_L g2176 ( 
.A1(n_2172),
.A2(n_2150),
.B(n_2105),
.C(n_2139),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2169),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_2175),
.Y(n_2178)
);

OAI222xp33_ASAP7_75t_L g2179 ( 
.A1(n_2174),
.A2(n_2139),
.B1(n_1995),
.B2(n_1924),
.C1(n_2126),
.C2(n_2109),
.Y(n_2179)
);

AOI221xp5_ASAP7_75t_L g2180 ( 
.A1(n_2176),
.A2(n_1752),
.B1(n_2054),
.B2(n_2063),
.C(n_2118),
.Y(n_2180)
);

BUFx2_ASAP7_75t_L g2181 ( 
.A(n_2173),
.Y(n_2181)
);

AOI22xp5_ASAP7_75t_L g2182 ( 
.A1(n_2177),
.A2(n_2051),
.B1(n_2045),
.B2(n_2029),
.Y(n_2182)
);

OR2x2_ASAP7_75t_L g2183 ( 
.A(n_2173),
.B(n_2124),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2175),
.B(n_2124),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_L g2185 ( 
.A1(n_2175),
.A2(n_2068),
.B1(n_2042),
.B2(n_2027),
.Y(n_2185)
);

OAI211xp5_ASAP7_75t_SL g2186 ( 
.A1(n_2174),
.A2(n_2004),
.B(n_1897),
.C(n_1875),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2173),
.B(n_2124),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2179),
.B(n_2022),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2178),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_2182),
.B(n_2004),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2181),
.B(n_2124),
.Y(n_2191)
);

NOR2xp67_ASAP7_75t_L g2192 ( 
.A(n_2183),
.B(n_142),
.Y(n_2192)
);

OA22x2_ASAP7_75t_L g2193 ( 
.A1(n_2184),
.A2(n_2118),
.B1(n_2123),
.B2(n_1959),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2180),
.B(n_2123),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2187),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_2185),
.B(n_2113),
.Y(n_2196)
);

OAI322xp33_ASAP7_75t_L g2197 ( 
.A1(n_2186),
.A2(n_1849),
.A3(n_1781),
.B1(n_1888),
.B2(n_1875),
.C1(n_1783),
.C2(n_1897),
.Y(n_2197)
);

AOI211xp5_ASAP7_75t_L g2198 ( 
.A1(n_2179),
.A2(n_2002),
.B(n_1993),
.C(n_1932),
.Y(n_2198)
);

AOI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_2179),
.A2(n_1984),
.B(n_1841),
.Y(n_2199)
);

AOI211xp5_ASAP7_75t_L g2200 ( 
.A1(n_2179),
.A2(n_1993),
.B(n_1932),
.C(n_1849),
.Y(n_2200)
);

AOI211xp5_ASAP7_75t_L g2201 ( 
.A1(n_2190),
.A2(n_146),
.B(n_143),
.C(n_145),
.Y(n_2201)
);

AOI322xp5_ASAP7_75t_L g2202 ( 
.A1(n_2189),
.A2(n_1760),
.A3(n_1939),
.B1(n_2110),
.B2(n_2096),
.C1(n_1756),
.C2(n_1779),
.Y(n_2202)
);

AOI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2188),
.A2(n_1915),
.B1(n_2048),
.B2(n_2012),
.Y(n_2203)
);

AOI221xp5_ASAP7_75t_L g2204 ( 
.A1(n_2191),
.A2(n_1837),
.B1(n_1883),
.B2(n_1860),
.C(n_1827),
.Y(n_2204)
);

OAI322xp33_ASAP7_75t_L g2205 ( 
.A1(n_2193),
.A2(n_145),
.A3(n_146),
.B1(n_147),
.B2(n_148),
.C1(n_149),
.C2(n_150),
.Y(n_2205)
);

AOI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_2200),
.A2(n_1892),
.B1(n_1940),
.B2(n_1930),
.C(n_149),
.Y(n_2206)
);

OAI221xp5_ASAP7_75t_SL g2207 ( 
.A1(n_2198),
.A2(n_2072),
.B1(n_1935),
.B2(n_1927),
.C(n_1894),
.Y(n_2207)
);

NAND4xp25_ASAP7_75t_SL g2208 ( 
.A(n_2194),
.B(n_2199),
.C(n_2196),
.D(n_2192),
.Y(n_2208)
);

AOI211xp5_ASAP7_75t_L g2209 ( 
.A1(n_2195),
.A2(n_150),
.B(n_147),
.C(n_148),
.Y(n_2209)
);

NAND3xp33_ASAP7_75t_L g2210 ( 
.A(n_2197),
.B(n_151),
.C(n_152),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2189),
.B(n_2092),
.Y(n_2211)
);

NAND3xp33_ASAP7_75t_SL g2212 ( 
.A(n_2189),
.B(n_151),
.C(n_152),
.Y(n_2212)
);

OAI21xp33_ASAP7_75t_L g2213 ( 
.A1(n_2188),
.A2(n_1981),
.B(n_2115),
.Y(n_2213)
);

AOI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_2208),
.A2(n_2048),
.B1(n_2055),
.B2(n_2012),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2212),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2211),
.Y(n_2216)
);

A2O1A1Ixp33_ASAP7_75t_SL g2217 ( 
.A1(n_2209),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2205),
.Y(n_2218)
);

AOI211x1_ASAP7_75t_L g2219 ( 
.A1(n_2213),
.A2(n_156),
.B(n_153),
.C(n_154),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2201),
.Y(n_2220)
);

BUFx2_ASAP7_75t_L g2221 ( 
.A(n_2203),
.Y(n_2221)
);

AND4x1_ASAP7_75t_L g2222 ( 
.A(n_2210),
.B(n_158),
.C(n_156),
.D(n_157),
.Y(n_2222)
);

INVxp67_ASAP7_75t_SL g2223 ( 
.A(n_2206),
.Y(n_2223)
);

AOI211x1_ASAP7_75t_SL g2224 ( 
.A1(n_2207),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_2204),
.A2(n_2202),
.B1(n_2048),
.B2(n_2055),
.Y(n_2225)
);

OAI22xp33_ASAP7_75t_L g2226 ( 
.A1(n_2203),
.A2(n_1930),
.B1(n_1934),
.B2(n_1923),
.Y(n_2226)
);

AOI221xp5_ASAP7_75t_L g2227 ( 
.A1(n_2218),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.C(n_162),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2215),
.A2(n_2012),
.B1(n_2055),
.B2(n_1930),
.Y(n_2228)
);

OAI221xp5_ASAP7_75t_L g2229 ( 
.A1(n_2214),
.A2(n_1918),
.B1(n_1941),
.B2(n_1969),
.C(n_1935),
.Y(n_2229)
);

AOI32xp33_ASAP7_75t_L g2230 ( 
.A1(n_2220),
.A2(n_1922),
.A3(n_1955),
.B1(n_1848),
.B2(n_1858),
.Y(n_2230)
);

NAND4xp75_ASAP7_75t_L g2231 ( 
.A(n_2219),
.B(n_164),
.C(n_162),
.D(n_163),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_2222),
.Y(n_2232)
);

AOI221xp5_ASAP7_75t_L g2233 ( 
.A1(n_2226),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_168),
.Y(n_2233)
);

AOI211xp5_ASAP7_75t_L g2234 ( 
.A1(n_2217),
.A2(n_168),
.B(n_165),
.C(n_166),
.Y(n_2234)
);

AOI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2221),
.A2(n_2223),
.B1(n_2225),
.B2(n_2216),
.C(n_2224),
.Y(n_2235)
);

AOI221xp5_ASAP7_75t_L g2236 ( 
.A1(n_2218),
.A2(n_172),
.B1(n_169),
.B2(n_170),
.C(n_173),
.Y(n_2236)
);

OAI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2214),
.A2(n_1918),
.B1(n_1941),
.B2(n_1922),
.C(n_1950),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2218),
.B(n_169),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2218),
.B(n_2099),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2217),
.A2(n_170),
.B(n_172),
.Y(n_2240)
);

AOI221xp5_ASAP7_75t_SL g2241 ( 
.A1(n_2226),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.C(n_177),
.Y(n_2241)
);

NAND4xp25_ASAP7_75t_SL g2242 ( 
.A(n_2225),
.B(n_177),
.C(n_174),
.D(n_175),
.Y(n_2242)
);

AOI221xp5_ASAP7_75t_L g2243 ( 
.A1(n_2218),
.A2(n_181),
.B1(n_178),
.B2(n_180),
.C(n_182),
.Y(n_2243)
);

NOR4xp25_ASAP7_75t_L g2244 ( 
.A(n_2242),
.B(n_182),
.C(n_178),
.D(n_180),
.Y(n_2244)
);

OAI211xp5_ASAP7_75t_SL g2245 ( 
.A1(n_2235),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_2245)
);

NOR3xp33_ASAP7_75t_L g2246 ( 
.A(n_2238),
.B(n_183),
.C(n_184),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2232),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_2239),
.B(n_1889),
.Y(n_2248)
);

A2O1A1Ixp33_ASAP7_75t_L g2249 ( 
.A1(n_2240),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_2249)
);

OAI21xp33_ASAP7_75t_L g2250 ( 
.A1(n_2234),
.A2(n_1923),
.B(n_1933),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2231),
.Y(n_2251)
);

OAI21xp33_ASAP7_75t_L g2252 ( 
.A1(n_2229),
.A2(n_1923),
.B(n_1931),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2227),
.B(n_187),
.Y(n_2253)
);

NAND3xp33_ASAP7_75t_L g2254 ( 
.A(n_2236),
.B(n_188),
.C(n_189),
.Y(n_2254)
);

OAI211xp5_ASAP7_75t_SL g2255 ( 
.A1(n_2243),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_2255)
);

AOI221xp5_ASAP7_75t_L g2256 ( 
.A1(n_2241),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.C(n_193),
.Y(n_2256)
);

NAND5xp2_ASAP7_75t_SL g2257 ( 
.A(n_2233),
.B(n_194),
.C(n_192),
.D(n_193),
.E(n_195),
.Y(n_2257)
);

INVx2_ASAP7_75t_SL g2258 ( 
.A(n_2228),
.Y(n_2258)
);

NOR4xp25_ASAP7_75t_SL g2259 ( 
.A(n_2237),
.B(n_196),
.C(n_194),
.D(n_195),
.Y(n_2259)
);

NAND3xp33_ASAP7_75t_L g2260 ( 
.A(n_2230),
.B(n_196),
.C(n_197),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_SL g2261 ( 
.A1(n_2240),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_2261)
);

OAI211xp5_ASAP7_75t_SL g2262 ( 
.A1(n_2235),
.A2(n_201),
.B(n_198),
.C(n_200),
.Y(n_2262)
);

OAI221xp5_ASAP7_75t_L g2263 ( 
.A1(n_2235),
.A2(n_1941),
.B1(n_203),
.B2(n_201),
.C(n_202),
.Y(n_2263)
);

OAI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2228),
.A2(n_1845),
.B1(n_1842),
.B2(n_1960),
.Y(n_2264)
);

NOR3xp33_ASAP7_75t_L g2265 ( 
.A(n_2238),
.B(n_202),
.C(n_203),
.Y(n_2265)
);

AOI221xp5_ASAP7_75t_L g2266 ( 
.A1(n_2242),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.C(n_208),
.Y(n_2266)
);

OAI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2228),
.A2(n_1999),
.B1(n_2081),
.B2(n_1990),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2231),
.Y(n_2268)
);

AOI222xp33_ASAP7_75t_L g2269 ( 
.A1(n_2235),
.A2(n_1889),
.B1(n_205),
.B2(n_206),
.C1(n_208),
.C2(n_209),
.Y(n_2269)
);

AOI22x1_ASAP7_75t_L g2270 ( 
.A1(n_2240),
.A2(n_211),
.B1(n_204),
.B2(n_210),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_SL g2271 ( 
.A1(n_2232),
.A2(n_1951),
.B1(n_2089),
.B2(n_1990),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2261),
.Y(n_2272)
);

NOR2x1_ASAP7_75t_L g2273 ( 
.A(n_2251),
.B(n_210),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2244),
.B(n_211),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2247),
.B(n_212),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2270),
.Y(n_2276)
);

AOI221xp5_ASAP7_75t_L g2277 ( 
.A1(n_2263),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.C(n_217),
.Y(n_2277)
);

NOR3xp33_ASAP7_75t_L g2278 ( 
.A(n_2245),
.B(n_217),
.C(n_220),
.Y(n_2278)
);

A2O1A1Ixp33_ASAP7_75t_L g2279 ( 
.A1(n_2266),
.A2(n_225),
.B(n_222),
.C(n_223),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2268),
.B(n_225),
.Y(n_2280)
);

NOR3xp33_ASAP7_75t_L g2281 ( 
.A(n_2262),
.B(n_226),
.C(n_227),
.Y(n_2281)
);

AOI221xp5_ASAP7_75t_L g2282 ( 
.A1(n_2256),
.A2(n_226),
.B1(n_227),
.B2(n_229),
.C(n_230),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2249),
.B(n_229),
.Y(n_2283)
);

NOR2x1p5_ASAP7_75t_L g2284 ( 
.A(n_2253),
.B(n_230),
.Y(n_2284)
);

NAND3xp33_ASAP7_75t_SL g2285 ( 
.A(n_2269),
.B(n_231),
.C(n_232),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2254),
.Y(n_2286)
);

AOI222xp33_ASAP7_75t_L g2287 ( 
.A1(n_2260),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.C1(n_236),
.C2(n_237),
.Y(n_2287)
);

AOI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_2257),
.A2(n_237),
.B(n_238),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2246),
.A2(n_1951),
.B1(n_2089),
.B2(n_1999),
.Y(n_2289)
);

OAI221xp5_ASAP7_75t_L g2290 ( 
.A1(n_2250),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.C(n_241),
.Y(n_2290)
);

AOI222xp33_ASAP7_75t_L g2291 ( 
.A1(n_2258),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.C1(n_243),
.C2(n_244),
.Y(n_2291)
);

AOI22xp33_ASAP7_75t_L g2292 ( 
.A1(n_2255),
.A2(n_1977),
.B1(n_1948),
.B2(n_1920),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2265),
.B(n_242),
.Y(n_2293)
);

NOR3xp33_ASAP7_75t_L g2294 ( 
.A(n_2252),
.B(n_243),
.C(n_244),
.Y(n_2294)
);

OAI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2248),
.A2(n_1920),
.B1(n_247),
.B2(n_245),
.Y(n_2295)
);

AOI211xp5_ASAP7_75t_L g2296 ( 
.A1(n_2290),
.A2(n_2285),
.B(n_2277),
.C(n_2282),
.Y(n_2296)
);

BUFx4f_ASAP7_75t_SL g2297 ( 
.A(n_2275),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2288),
.B(n_2259),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2275),
.Y(n_2299)
);

NAND5xp2_ASAP7_75t_L g2300 ( 
.A(n_2272),
.B(n_2271),
.C(n_2248),
.D(n_2267),
.E(n_2264),
.Y(n_2300)
);

NOR2xp67_ASAP7_75t_SL g2301 ( 
.A(n_2280),
.B(n_245),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2274),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2273),
.Y(n_2303)
);

OAI22xp5_ASAP7_75t_L g2304 ( 
.A1(n_2292),
.A2(n_249),
.B1(n_246),
.B2(n_248),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2283),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2278),
.B(n_246),
.Y(n_2306)
);

AOI221x1_ASAP7_75t_L g2307 ( 
.A1(n_2286),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.C(n_252),
.Y(n_2307)
);

NAND3xp33_ASAP7_75t_SL g2308 ( 
.A(n_2287),
.B(n_250),
.C(n_251),
.Y(n_2308)
);

XNOR2x1_ASAP7_75t_L g2309 ( 
.A(n_2284),
.B(n_252),
.Y(n_2309)
);

NOR2x1_ASAP7_75t_L g2310 ( 
.A(n_2276),
.B(n_253),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2293),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2294),
.B(n_255),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2295),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2281),
.B(n_255),
.Y(n_2314)
);

OAI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2279),
.A2(n_256),
.B(n_257),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2291),
.B(n_256),
.Y(n_2316)
);

NAND4xp75_ASAP7_75t_L g2317 ( 
.A(n_2289),
.B(n_260),
.C(n_258),
.D(n_259),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2272),
.B(n_258),
.Y(n_2318)
);

AND2x4_ASAP7_75t_L g2319 ( 
.A(n_2273),
.B(n_259),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2288),
.B(n_260),
.Y(n_2320)
);

BUFx2_ASAP7_75t_L g2321 ( 
.A(n_2273),
.Y(n_2321)
);

NOR4xp25_ASAP7_75t_L g2322 ( 
.A(n_2272),
.B(n_265),
.C(n_261),
.D(n_264),
.Y(n_2322)
);

NAND5xp2_ASAP7_75t_L g2323 ( 
.A(n_2272),
.B(n_261),
.C(n_265),
.D(n_266),
.E(n_267),
.Y(n_2323)
);

AOI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2318),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_2324)
);

AND4x1_ASAP7_75t_L g2325 ( 
.A(n_2322),
.B(n_268),
.C(n_269),
.D(n_270),
.Y(n_2325)
);

NOR3xp33_ASAP7_75t_L g2326 ( 
.A(n_2320),
.B(n_269),
.C(n_270),
.Y(n_2326)
);

AOI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2304),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.C(n_275),
.Y(n_2327)
);

OAI211xp5_ASAP7_75t_SL g2328 ( 
.A1(n_2298),
.A2(n_272),
.B(n_274),
.C(n_275),
.Y(n_2328)
);

OAI211xp5_ASAP7_75t_L g2329 ( 
.A1(n_2315),
.A2(n_276),
.B(n_277),
.C(n_278),
.Y(n_2329)
);

OAI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_2297),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2319),
.B(n_279),
.Y(n_2331)
);

NOR3xp33_ASAP7_75t_SL g2332 ( 
.A(n_2308),
.B(n_279),
.C(n_280),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2319),
.Y(n_2333)
);

O2A1O1Ixp5_ASAP7_75t_L g2334 ( 
.A1(n_2303),
.A2(n_2313),
.B(n_2312),
.C(n_2299),
.Y(n_2334)
);

BUFx2_ASAP7_75t_L g2335 ( 
.A(n_2310),
.Y(n_2335)
);

OAI211xp5_ASAP7_75t_L g2336 ( 
.A1(n_2314),
.A2(n_280),
.B(n_281),
.C(n_282),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_L g2337 ( 
.A(n_2301),
.B(n_281),
.C(n_282),
.Y(n_2337)
);

NOR2x1_ASAP7_75t_L g2338 ( 
.A(n_2321),
.B(n_283),
.Y(n_2338)
);

NAND4xp25_ASAP7_75t_L g2339 ( 
.A(n_2296),
.B(n_283),
.C(n_284),
.D(n_285),
.Y(n_2339)
);

NOR3xp33_ASAP7_75t_L g2340 ( 
.A(n_2302),
.B(n_285),
.C(n_286),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2323),
.B(n_287),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2312),
.B(n_2316),
.Y(n_2342)
);

NAND4xp25_ASAP7_75t_L g2343 ( 
.A(n_2300),
.B(n_287),
.C(n_288),
.D(n_289),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2309),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2306),
.B(n_288),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2341),
.Y(n_2346)
);

OR3x1_ASAP7_75t_L g2347 ( 
.A(n_2343),
.B(n_2305),
.C(n_2311),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2338),
.Y(n_2348)
);

AND2x2_ASAP7_75t_SL g2349 ( 
.A(n_2325),
.B(n_2307),
.Y(n_2349)
);

BUFx2_ASAP7_75t_L g2350 ( 
.A(n_2335),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2340),
.B(n_2317),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2331),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_2333),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2342),
.B(n_290),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2345),
.Y(n_2355)
);

INVx3_ASAP7_75t_L g2356 ( 
.A(n_2342),
.Y(n_2356)
);

AND3x1_ASAP7_75t_L g2357 ( 
.A(n_2326),
.B(n_291),
.C(n_292),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2334),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2339),
.B(n_291),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2337),
.Y(n_2360)
);

INVxp67_ASAP7_75t_L g2361 ( 
.A(n_2330),
.Y(n_2361)
);

NAND4xp75_ASAP7_75t_L g2362 ( 
.A(n_2344),
.B(n_293),
.C(n_294),
.D(n_295),
.Y(n_2362)
);

INVxp67_ASAP7_75t_L g2363 ( 
.A(n_2324),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2332),
.B(n_293),
.Y(n_2364)
);

NOR3xp33_ASAP7_75t_SL g2365 ( 
.A(n_2329),
.B(n_296),
.C(n_297),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2336),
.Y(n_2366)
);

OAI22x1_ASAP7_75t_L g2367 ( 
.A1(n_2358),
.A2(n_2328),
.B1(n_2327),
.B2(n_300),
.Y(n_2367)
);

AOI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_2356),
.A2(n_296),
.B1(n_299),
.B2(n_300),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_2362),
.Y(n_2369)
);

OAI22x1_ASAP7_75t_L g2370 ( 
.A1(n_2350),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_2370)
);

AO22x2_ASAP7_75t_SL g2371 ( 
.A1(n_2346),
.A2(n_301),
.B1(n_355),
.B2(n_356),
.Y(n_2371)
);

AO22x2_ASAP7_75t_L g2372 ( 
.A1(n_2348),
.A2(n_2355),
.B1(n_2366),
.B2(n_2360),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2361),
.A2(n_357),
.B1(n_362),
.B2(n_363),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2357),
.A2(n_2347),
.B1(n_2363),
.B2(n_2353),
.Y(n_2374)
);

BUFx3_ASAP7_75t_L g2375 ( 
.A(n_2353),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2359),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_2376)
);

AOI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_2364),
.A2(n_2349),
.B1(n_2351),
.B2(n_2352),
.Y(n_2377)
);

AOI22xp5_ASAP7_75t_SL g2378 ( 
.A1(n_2354),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_2378)
);

CKINVDCx20_ASAP7_75t_R g2379 ( 
.A(n_2365),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2354),
.Y(n_2380)
);

INVx8_ASAP7_75t_L g2381 ( 
.A(n_2353),
.Y(n_2381)
);

INVx1_ASAP7_75t_SL g2382 ( 
.A(n_2349),
.Y(n_2382)
);

AND4x2_ASAP7_75t_L g2383 ( 
.A(n_2357),
.B(n_371),
.C(n_373),
.D(n_376),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2381),
.B(n_378),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2370),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2381),
.B(n_379),
.Y(n_2386)
);

AOI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_2379),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2383),
.Y(n_2388)
);

AOI31xp33_ASAP7_75t_L g2389 ( 
.A1(n_2369),
.A2(n_384),
.A3(n_388),
.B(n_389),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2380),
.B(n_390),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2382),
.A2(n_391),
.B1(n_393),
.B2(n_394),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2375),
.Y(n_2392)
);

AOI22xp33_ASAP7_75t_L g2393 ( 
.A1(n_2372),
.A2(n_2374),
.B1(n_2367),
.B2(n_2377),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2392),
.A2(n_2376),
.B1(n_2368),
.B2(n_2373),
.Y(n_2394)
);

OAI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2393),
.A2(n_2378),
.B1(n_2371),
.B2(n_397),
.Y(n_2395)
);

NAND4xp25_ASAP7_75t_L g2396 ( 
.A(n_2388),
.B(n_2390),
.C(n_2386),
.D(n_2384),
.Y(n_2396)
);

OAI22xp5_ASAP7_75t_SL g2397 ( 
.A1(n_2385),
.A2(n_395),
.B1(n_396),
.B2(n_398),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2387),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_2398)
);

NAND5xp2_ASAP7_75t_L g2399 ( 
.A(n_2391),
.B(n_402),
.C(n_406),
.D(n_407),
.E(n_408),
.Y(n_2399)
);

AOI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_2389),
.A2(n_409),
.B1(n_412),
.B2(n_413),
.Y(n_2400)
);

AOI22xp33_ASAP7_75t_L g2401 ( 
.A1(n_2392),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_2401)
);

AOI222xp33_ASAP7_75t_L g2402 ( 
.A1(n_2385),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.C1(n_421),
.C2(n_424),
.Y(n_2402)
);

AOI31xp33_ASAP7_75t_L g2403 ( 
.A1(n_2395),
.A2(n_425),
.A3(n_428),
.B(n_429),
.Y(n_2403)
);

AOI31xp33_ASAP7_75t_L g2404 ( 
.A1(n_2394),
.A2(n_430),
.A3(n_431),
.B(n_433),
.Y(n_2404)
);

AOI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2396),
.A2(n_434),
.B1(n_435),
.B2(n_436),
.Y(n_2405)
);

AOI31xp33_ASAP7_75t_L g2406 ( 
.A1(n_2400),
.A2(n_438),
.A3(n_440),
.B(n_445),
.Y(n_2406)
);

AOI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2405),
.A2(n_2398),
.B1(n_2397),
.B2(n_2402),
.Y(n_2407)
);

XNOR2xp5_ASAP7_75t_L g2408 ( 
.A(n_2403),
.B(n_2401),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2408),
.A2(n_2406),
.B(n_2404),
.Y(n_2409)
);

NOR2x1_ASAP7_75t_L g2410 ( 
.A(n_2407),
.B(n_2399),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2410),
.Y(n_2411)
);

XNOR2xp5_ASAP7_75t_L g2412 ( 
.A(n_2411),
.B(n_2409),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2411),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2413),
.B(n_447),
.Y(n_2414)
);

A2O1A1Ixp33_ASAP7_75t_L g2415 ( 
.A1(n_2414),
.A2(n_2412),
.B(n_450),
.C(n_451),
.Y(n_2415)
);

AOI211xp5_ASAP7_75t_L g2416 ( 
.A1(n_2415),
.A2(n_449),
.B(n_453),
.C(n_454),
.Y(n_2416)
);


endmodule