module real_jpeg_25796_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_42),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_2),
.A2(n_25),
.B(n_32),
.C(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_30),
.B1(n_32),
.B2(n_81),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_2),
.B(n_49),
.C(n_67),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_81),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_2),
.A2(n_52),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_2),
.B(n_96),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_5),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_73),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_6),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_73),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_35),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_9),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_12),
.A2(n_53),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_98),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_97),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_87),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_17),
.B(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_61),
.B2(n_86),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_22),
.A2(n_23),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_22),
.A2(n_26),
.B(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_23),
.B(n_105),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_34),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_37),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_52),
.B1(n_56),
.B2(n_58),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_54),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_49),
.B1(n_67),
.B2(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_48),
.B(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_52),
.A2(n_113),
.B(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_85),
.Y(n_84)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_77),
.B2(n_78),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_74),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_64),
.A2(n_74),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_72),
.B1(n_76),
.B2(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_65),
.B(n_75),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_81),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_70),
.A2(n_91),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_111),
.B(n_123),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.C(n_92),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_140),
.B(n_145),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_129),
.B(n_139),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_114),
.B(n_128),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_109),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_124),
.B(n_127),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_138),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_138),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_135),
.C(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_144),
.Y(n_145)
);


endmodule