module fake_jpeg_2289_n_220 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_220);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_24),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_6),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_31),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_41),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_34),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_9),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_84),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_87),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_63),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_70),
.B1(n_63),
.B2(n_68),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_100),
.B1(n_69),
.B2(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_60),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_68),
.B1(n_74),
.B2(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_64),
.B1(n_62),
.B2(n_57),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_74),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_63),
.B1(n_71),
.B2(n_73),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_79),
.B(n_82),
.C(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_119),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_111),
.B1(n_21),
.B2(n_49),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_62),
.B1(n_66),
.B2(n_69),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_66),
.B1(n_77),
.B2(n_76),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_2),
.B(n_3),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_65),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_59),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

OR2x2_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_78),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_0),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_4),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_90),
.B(n_19),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_136),
.B1(n_115),
.B2(n_5),
.Y(n_142)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

CKINVDCx12_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_53),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_1),
.B(n_2),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_51),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_22),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_3),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_7),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_145),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_104),
.B(n_110),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_156),
.B(n_161),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_7),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_164),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_23),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_159),
.C(n_162),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_124),
.B(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_26),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_110),
.B(n_9),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_48),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_11),
.B(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_8),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_10),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_30),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_172),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_128),
.C(n_29),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_175),
.C(n_161),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_130),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

AND2x4_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_144),
.Y(n_188)
);

FAx1_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_180),
.CI(n_172),
.CON(n_202),
.SN(n_202)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_193),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_146),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_167),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_162),
.C(n_151),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_200),
.C(n_192),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_169),
.B1(n_142),
.B2(n_184),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_199),
.B1(n_203),
.B2(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_198),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_181),
.B1(n_180),
.B2(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_202),
.B(n_194),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_195),
.A2(n_182),
.B1(n_163),
.B2(n_14),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_196),
.C(n_185),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_208),
.B1(n_188),
.B2(n_28),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_195),
.B1(n_194),
.B2(n_188),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_46),
.B1(n_43),
.B2(n_40),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_211),
.B(n_207),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_206),
.B(n_37),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_33),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_212),
.B(n_13),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_216),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_SL g218 ( 
.A1(n_217),
.A2(n_15),
.B(n_16),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_17),
.B(n_18),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_18),
.Y(n_220)
);


endmodule