module fake_jpeg_17036_n_360 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_6),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_6),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_46),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_22),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_88)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_28),
.Y(n_87)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_69),
.B(n_89),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_81),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_76),
.A2(n_77),
.B1(n_108),
.B2(n_5),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_27),
.B1(n_22),
.B2(n_34),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_79),
.A2(n_86),
.B1(n_110),
.B2(n_20),
.Y(n_122)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

FAx1_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_19),
.CI(n_28),
.CON(n_84),
.SN(n_84)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_94),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_22),
.B1(n_27),
.B2(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_14),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_15),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_91),
.B(n_93),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_35),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_32),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_21),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_21),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_16),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_47),
.A2(n_16),
.B1(n_14),
.B2(n_36),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_50),
.A2(n_36),
.B1(n_20),
.B2(n_3),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_45),
.B(n_36),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_8),
.Y(n_146)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_20),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_118),
.A2(n_123),
.B(n_132),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_124),
.Y(n_189)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_122),
.A2(n_126),
.B1(n_138),
.B2(n_150),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_7),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_127),
.B(n_143),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_73),
.A2(n_104),
.B1(n_82),
.B2(n_99),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_130),
.A2(n_131),
.B1(n_137),
.B2(n_147),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_73),
.A2(n_7),
.B1(n_2),
.B2(n_4),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_10),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_10),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_142),
.Y(n_169)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_104),
.A2(n_10),
.B1(n_5),
.B2(n_6),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_75),
.B(n_66),
.CI(n_77),
.CON(n_139),
.SN(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_134),
.B(n_141),
.C(n_145),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_72),
.B(n_5),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_82),
.A2(n_0),
.B1(n_8),
.B2(n_11),
.Y(n_147)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_8),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_165),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_163),
.B1(n_68),
.B2(n_80),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_67),
.A2(n_0),
.B1(n_12),
.B2(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_12),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_153),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_70),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_71),
.B(n_109),
.C(n_114),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_160),
.C(n_140),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_97),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_112),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_78),
.B(n_81),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_98),
.B1(n_112),
.B2(n_107),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_107),
.Y(n_165)
);

NOR2xp67_ASAP7_75t_R g166 ( 
.A(n_125),
.B(n_99),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_166),
.A2(n_190),
.B(n_208),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_117),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_168),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_156),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_170),
.A2(n_188),
.B(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_160),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_180),
.Y(n_219)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_154),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_174),
.A2(n_178),
.B1(n_207),
.B2(n_170),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_114),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_179),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_125),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_135),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_135),
.B1(n_128),
.B2(n_159),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_193),
.B1(n_164),
.B2(n_116),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_123),
.B1(n_132),
.B2(n_122),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_186),
.A2(n_147),
.B1(n_151),
.B2(n_120),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_123),
.B(n_132),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_200),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_128),
.A2(n_129),
.B1(n_159),
.B2(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_133),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_206),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_157),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_160),
.B1(n_118),
.B2(n_158),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_139),
.B(n_119),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_124),
.B(n_139),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_134),
.B(n_142),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_118),
.B(n_127),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_133),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_201),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_215),
.C(n_247),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_158),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_220),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_218),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_163),
.B1(n_136),
.B2(n_121),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_224),
.B1(n_226),
.B2(n_233),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_196),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_182),
.A2(n_121),
.B1(n_155),
.B2(n_140),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_185),
.B1(n_200),
.B2(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_179),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_231),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_191),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_199),
.B1(n_186),
.B2(n_197),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_187),
.A2(n_199),
.B1(n_171),
.B2(n_192),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_260)
);

A2O1A1O1Ixp25_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_200),
.B(n_208),
.C(n_169),
.D(n_206),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_243),
.A3(n_175),
.B1(n_184),
.B2(n_198),
.C1(n_203),
.C2(n_232),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_173),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_236),
.B(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_168),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_170),
.B1(n_204),
.B2(n_174),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_190),
.A2(n_169),
.A3(n_202),
.B1(n_176),
.B2(n_180),
.C1(n_189),
.C2(n_167),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_189),
.A2(n_176),
.B1(n_209),
.B2(n_194),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_246),
.Y(n_252)
);

NAND2x1_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_201),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_254),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_237),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_257),
.A2(n_220),
.B(n_225),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_175),
.Y(n_258)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_184),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_259),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_233),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_268),
.C(n_271),
.Y(n_302)
);

AOI221xp5_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_260),
.B1(n_273),
.B2(n_253),
.C(n_267),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_239),
.A2(n_203),
.B1(n_242),
.B2(n_221),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_267),
.B1(n_276),
.B2(n_278),
.Y(n_296)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_213),
.A2(n_241),
.B1(n_231),
.B2(n_210),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_213),
.B(n_212),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_217),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_269),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_240),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_270),
.B(n_274),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_214),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_215),
.C(n_234),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_218),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_224),
.B1(n_210),
.B2(n_211),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_273),
.A2(n_260),
.B1(n_253),
.B2(n_257),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_236),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_275),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_241),
.A2(n_216),
.B1(n_211),
.B2(n_247),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_225),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_248),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_222),
.B(n_219),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_281),
.A2(n_288),
.B(n_292),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_247),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_286),
.C(n_255),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_223),
.Y(n_285)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_290),
.B(n_252),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_250),
.A2(n_229),
.B(n_272),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_229),
.B(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_296),
.B(n_268),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_300),
.B1(n_284),
.B2(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_301),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_262),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_264),
.A2(n_255),
.B1(n_256),
.B2(n_252),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_248),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_291),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_310),
.C(n_311),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_249),
.Y(n_305)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_305),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_316),
.B(n_287),
.Y(n_323)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_309),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_270),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_254),
.C(n_277),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_274),
.B(n_266),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_294),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_318),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_279),
.B1(n_303),
.B2(n_285),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_300),
.C(n_286),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_288),
.C(n_297),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_284),
.A2(n_280),
.B1(n_289),
.B2(n_296),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_315),
.B1(n_308),
.B2(n_314),
.Y(n_326)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_326),
.A2(n_330),
.B(n_323),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_330),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_329),
.C(n_331),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_281),
.C(n_295),
.Y(n_329)
);

AOI31xp33_ASAP7_75t_SL g330 ( 
.A1(n_316),
.A2(n_283),
.A3(n_294),
.B(n_301),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_293),
.C(n_298),
.Y(n_331)
);

NAND4xp25_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_283),
.C(n_289),
.D(n_306),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_332),
.A2(n_333),
.B1(n_313),
.B2(n_322),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_315),
.A2(n_318),
.B(n_312),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_312),
.Y(n_336)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_304),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_338),
.C(n_331),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_310),
.Y(n_338)
);

FAx1_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_307),
.CI(n_322),
.CON(n_340),
.SN(n_340)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_340),
.B(n_327),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_341),
.A2(n_345),
.B(n_329),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_313),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_344),
.B(n_343),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_346),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_342),
.A2(n_333),
.B(n_334),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_347),
.B(n_348),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_349),
.B(n_350),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_339),
.C(n_325),
.Y(n_355)
);

AO21x1_ASAP7_75t_L g357 ( 
.A1(n_355),
.A2(n_356),
.B(n_351),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_352),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_349),
.B(n_353),
.Y(n_358)
);

AOI21x1_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_341),
.B(n_340),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_340),
.Y(n_360)
);


endmodule