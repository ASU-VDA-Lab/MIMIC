module fake_jpeg_18333_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_31),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_36),
.B1(n_14),
.B2(n_26),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_37),
.Y(n_38)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_23),
.B1(n_18),
.B2(n_27),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_27),
.B1(n_25),
.B2(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_46),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_24),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_22),
.C(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_38),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

OA22x2_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_14),
.B1(n_26),
.B2(n_22),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_31),
.B1(n_34),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_31),
.B1(n_34),
.B2(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_58),
.B(n_71),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_24),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_22),
.C(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_25),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_16),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_15),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_12),
.B1(n_8),
.B2(n_7),
.Y(n_86)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_28),
.B(n_1),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_82),
.C(n_71),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_19),
.C(n_6),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_56),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_65),
.B(n_69),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_95),
.B(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_65),
.B1(n_53),
.B2(n_66),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_97),
.B1(n_88),
.B2(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_74),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_73),
.C(n_76),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_74),
.C(n_73),
.Y(n_101)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_70),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_55),
.B(n_56),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_72),
.B1(n_55),
.B2(n_59),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

AO221x1_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_52),
.B1(n_61),
.B2(n_95),
.C(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_102),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_106),
.C(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_80),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_98),
.B1(n_93),
.B2(n_75),
.Y(n_112)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_77),
.B(n_90),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_96),
.B1(n_98),
.B2(n_55),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_112),
.B1(n_106),
.B2(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_117),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_113),
.C(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

XNOR2x1_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_116),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_109),
.B(n_82),
.C(n_78),
.Y(n_124)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_99),
.B(n_75),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_121),
.Y(n_123)
);

AOI222xp33_ASAP7_75t_SL g126 ( 
.A1(n_124),
.A2(n_122),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_81),
.C(n_12),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_0),
.Y(n_129)
);


endmodule