module fake_ibex_126_n_844 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_91, n_54, n_19, n_844);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_844;

wire n_151;
wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_144;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_820;
wire n_805;
wire n_670;
wire n_728;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_794;
wire n_260;
wire n_620;
wire n_683;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_159;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_51),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_14),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_43),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_27),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_65),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_90),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_45),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_59),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_35),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_82),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_54),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_20),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_12),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_31),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_L g167 ( 
.A(n_48),
.B(n_46),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_35),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_29),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_49),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_106),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_109),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_79),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_93),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_76),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_61),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_34),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_53),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_29),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_13),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_122),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_31),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_40),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_56),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_62),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_70),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_96),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_7),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_21),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_10),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_91),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_13),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_32),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_97),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_2),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_1),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_47),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_33),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_50),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_102),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_23),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_28),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_32),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_72),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_80),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_17),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_100),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_41),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_64),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_86),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_38),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_24),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_83),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_41),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_131),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_69),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_99),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_126),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_22),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_38),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_74),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_105),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g243 ( 
.A(n_95),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_139),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_27),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_116),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_55),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_119),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_98),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_14),
.Y(n_250)
);

INVx4_ASAP7_75t_R g251 ( 
.A(n_44),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_18),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_141),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_40),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_104),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_36),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_123),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_147),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_218),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_197),
.B(n_0),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_3),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_158),
.A2(n_71),
.B(n_138),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_173),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_197),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g267 ( 
.A1(n_158),
.A2(n_66),
.B(n_137),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_219),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_147),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_151),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_151),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_193),
.B(n_5),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_183),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_189),
.B(n_6),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_237),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_146),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_237),
.Y(n_282)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_77),
.B(n_132),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_208),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_150),
.B(n_8),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_232),
.A2(n_81),
.B(n_130),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_237),
.B(n_10),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_150),
.B(n_11),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_173),
.Y(n_292)
);

BUFx8_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_219),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_294)
);

XNOR2x2_ASAP7_75t_L g295 ( 
.A(n_145),
.B(n_15),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_239),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_L g297 ( 
.A(n_153),
.B(n_84),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_163),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_223),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_173),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_202),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_191),
.B(n_140),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_142),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_143),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_173),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_149),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_202),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_153),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_144),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_148),
.B(n_16),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_156),
.B(n_18),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_152),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_146),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_202),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_169),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_202),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_154),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_155),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_169),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_160),
.B(n_19),
.Y(n_321)
);

XOR2x2_ASAP7_75t_L g322 ( 
.A(n_162),
.B(n_22),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_164),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_168),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_171),
.Y(n_325)
);

OAI22x1_ASAP7_75t_L g326 ( 
.A1(n_170),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_166),
.B(n_25),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_178),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_170),
.A2(n_213),
.B1(n_225),
.B2(n_209),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_172),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_187),
.B(n_26),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_201),
.B(n_28),
.Y(n_332)
);

BUFx8_ASAP7_75t_SL g333 ( 
.A(n_163),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_174),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_192),
.B(n_195),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_175),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_177),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_179),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g339 ( 
.A(n_157),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_181),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g341 ( 
.A1(n_201),
.A2(n_225),
.B1(n_203),
.B2(n_204),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_182),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_185),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_261),
.B(n_186),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

AND2x6_ASAP7_75t_L g346 ( 
.A(n_261),
.B(n_188),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_209),
.C(n_204),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_198),
.Y(n_348)
);

BUFx4f_ASAP7_75t_L g349 ( 
.A(n_303),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

NAND2x1p5_ASAP7_75t_L g351 ( 
.A(n_285),
.B(n_196),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_213),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_303),
.A2(n_244),
.B1(n_245),
.B2(n_241),
.Y(n_354)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_258),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_276),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_L g357 ( 
.A(n_290),
.B(n_159),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_264),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_303),
.A2(n_220),
.B1(n_256),
.B2(n_254),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_216),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_276),
.B(n_200),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_320),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_245),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_329),
.A2(n_217),
.B1(n_241),
.B2(n_236),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_L g367 ( 
.A(n_290),
.B(n_159),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_307),
.Y(n_368)
);

AND3x1_ASAP7_75t_L g369 ( 
.A(n_272),
.B(n_230),
.C(n_231),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_311),
.A2(n_212),
.B1(n_215),
.B2(n_250),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_335),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_333),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_305),
.B(n_205),
.Y(n_373)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_276),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_341),
.A2(n_217),
.B1(n_236),
.B2(n_234),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_335),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_279),
.B(n_214),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_305),
.B(n_206),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_300),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_311),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_161),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_272),
.Y(n_383)
);

AO22x2_ASAP7_75t_L g384 ( 
.A1(n_260),
.A2(n_316),
.B1(n_311),
.B2(n_312),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_298),
.A2(n_227),
.B1(n_207),
.B2(n_240),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_339),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g387 ( 
.A(n_307),
.B(n_161),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_300),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_318),
.B(n_210),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_324),
.B(n_165),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_211),
.Y(n_394)
);

BUFx10_ASAP7_75t_L g395 ( 
.A(n_331),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_264),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_334),
.B(n_336),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_331),
.B(n_221),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_334),
.B(n_222),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_297),
.B(n_224),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_296),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_299),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_264),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_340),
.B(n_180),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_228),
.Y(n_405)
);

INVx4_ASAP7_75t_SL g406 ( 
.A(n_319),
.Y(n_406)
);

BUFx8_ASAP7_75t_SL g407 ( 
.A(n_332),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_342),
.A2(n_246),
.B1(n_229),
.B2(n_238),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_265),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_293),
.A2(n_235),
.B1(n_253),
.B2(n_180),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_304),
.B(n_194),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_304),
.B(n_194),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_265),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_325),
.B(n_330),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_263),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_325),
.Y(n_418)
);

AND3x2_ASAP7_75t_L g419 ( 
.A(n_295),
.B(n_248),
.C(n_184),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_310),
.B(n_233),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_262),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_325),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_330),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_313),
.B(n_249),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_323),
.B(n_247),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_322),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_323),
.B(n_226),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_337),
.B(n_226),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_330),
.B(n_242),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_327),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_330),
.B(n_242),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_337),
.B(n_243),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_266),
.B(n_167),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_338),
.B(n_343),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_343),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_266),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_322),
.Y(n_437)
);

BUFx4f_ASAP7_75t_L g438 ( 
.A(n_263),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_277),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_268),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_277),
.B(n_257),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_278),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_259),
.B(n_269),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_259),
.B(n_176),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_269),
.A2(n_199),
.B1(n_190),
.B2(n_251),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_270),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_278),
.B(n_92),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_270),
.B(n_30),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_280),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_271),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_271),
.B(n_30),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_273),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_280),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_377),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_371),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_377),
.B(n_274),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_371),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_349),
.A2(n_289),
.B1(n_282),
.B2(n_295),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_430),
.Y(n_462)
);

AND2x2_ASAP7_75t_SL g463 ( 
.A(n_349),
.B(n_263),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_365),
.B(n_275),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_360),
.A2(n_294),
.B1(n_288),
.B2(n_326),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_382),
.B(n_284),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_393),
.B(n_291),
.Y(n_467)
);

AO22x1_ASAP7_75t_L g468 ( 
.A1(n_368),
.A2(n_326),
.B1(n_287),
.B2(n_291),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_347),
.B(n_282),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_404),
.B(n_289),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_428),
.B(n_435),
.Y(n_471)
);

OAI22xp33_ASAP7_75t_L g472 ( 
.A1(n_354),
.A2(n_440),
.B1(n_383),
.B2(n_376),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_348),
.B(n_286),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_364),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_383),
.B(n_352),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_438),
.A2(n_267),
.B(n_283),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

O2A1O1Ixp5_ASAP7_75t_L g478 ( 
.A1(n_417),
.A2(n_302),
.B(n_283),
.C(n_286),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_372),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_351),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_363),
.A2(n_267),
.B1(n_283),
.B2(n_286),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_395),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_378),
.B(n_302),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_361),
.B(n_286),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_428),
.B(n_267),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_413),
.B(n_414),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_420),
.B(n_267),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_361),
.B(n_292),
.Y(n_488)
);

OAI22xp33_ASAP7_75t_L g489 ( 
.A1(n_351),
.A2(n_317),
.B1(n_315),
.B2(n_308),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_427),
.B(n_292),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_443),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_398),
.B(n_317),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_388),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_369),
.A2(n_384),
.B1(n_357),
.B2(n_367),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_384),
.A2(n_317),
.B1(n_315),
.B2(n_308),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_444),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_389),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_344),
.B(n_315),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_SL g500 ( 
.A1(n_384),
.A2(n_315),
.B1(n_308),
.B2(n_306),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_350),
.B(n_306),
.Y(n_504)
);

AO221x2_ASAP7_75t_L g505 ( 
.A1(n_385),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.C(n_39),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_434),
.Y(n_506)
);

AND2x6_ASAP7_75t_SL g507 ( 
.A(n_426),
.B(n_37),
.Y(n_507)
);

NOR2x1p5_ASAP7_75t_L g508 ( 
.A(n_386),
.B(n_39),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_407),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_362),
.B(n_301),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_353),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_359),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_418),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_375),
.B(n_301),
.Y(n_514)
);

BUFx4f_ASAP7_75t_L g515 ( 
.A(n_363),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_380),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_390),
.Y(n_517)
);

AND2x4_ASAP7_75t_SL g518 ( 
.A(n_411),
.B(n_306),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_423),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_356),
.B(n_264),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_363),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_391),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_355),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_391),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_446),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_381),
.B(n_52),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_450),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_355),
.B(n_57),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_370),
.B(n_58),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_387),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_400),
.B(n_345),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_370),
.A2(n_445),
.B1(n_400),
.B2(n_408),
.Y(n_532)
);

BUFx12f_ASAP7_75t_SL g533 ( 
.A(n_425),
.Y(n_533)
);

BUFx4f_ASAP7_75t_L g534 ( 
.A(n_455),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_506),
.Y(n_535)
);

O2A1O1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_532),
.A2(n_397),
.B(n_344),
.C(n_373),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_491),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_480),
.B(n_425),
.Y(n_538)
);

A2O1A1Ixp33_ASAP7_75t_L g539 ( 
.A1(n_464),
.A2(n_405),
.B(n_394),
.C(n_399),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_462),
.B(n_346),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_500),
.A2(n_408),
.B1(n_379),
.B2(n_405),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_494),
.Y(n_542)
);

AND2x2_ASAP7_75t_SL g543 ( 
.A(n_515),
.B(n_445),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_487),
.A2(n_441),
.B(n_431),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_478),
.A2(n_436),
.B(n_453),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_465),
.A2(n_419),
.B(n_432),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_495),
.B(n_441),
.C(n_429),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_419),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_482),
.B(n_415),
.Y(n_549)
);

AO21x1_ASAP7_75t_L g550 ( 
.A1(n_473),
.A2(n_447),
.B(n_433),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_496),
.A2(n_379),
.B1(n_399),
.B2(n_394),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_523),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_485),
.A2(n_473),
.B(n_484),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_457),
.Y(n_554)
);

O2A1O1Ixp33_ASAP7_75t_L g555 ( 
.A1(n_472),
.A2(n_531),
.B(n_475),
.C(n_474),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_454),
.B(n_401),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_SL g557 ( 
.A(n_472),
.B(n_392),
.C(n_424),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_509),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_522),
.Y(n_559)
);

BUFx12f_ASAP7_75t_L g560 ( 
.A(n_479),
.Y(n_560)
);

O2A1O1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_531),
.A2(n_474),
.B(n_501),
.C(n_471),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_454),
.B(n_452),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_SL g563 ( 
.A1(n_456),
.A2(n_448),
.B1(n_402),
.B2(n_449),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_525),
.B(n_442),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_484),
.A2(n_439),
.B(n_429),
.C(n_433),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_524),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_480),
.B(n_406),
.Y(n_567)
);

A2O1A1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_486),
.A2(n_416),
.B(n_422),
.C(n_403),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_463),
.A2(n_403),
.B(n_396),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_530),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_507),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_463),
.A2(n_396),
.B(n_358),
.Y(n_574)
);

AO21x1_ASAP7_75t_L g575 ( 
.A1(n_528),
.A2(n_60),
.B(n_63),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_470),
.A2(n_481),
.B(n_520),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_468),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_520),
.A2(n_477),
.B(n_514),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_514),
.A2(n_358),
.B(n_89),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_466),
.B(n_127),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_483),
.B(n_124),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_459),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_467),
.B(n_118),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_529),
.A2(n_469),
.B1(n_459),
.B2(n_483),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_505),
.A2(n_469),
.B1(n_461),
.B2(n_460),
.Y(n_585)
);

CKINVDCx8_ASAP7_75t_R g586 ( 
.A(n_460),
.Y(n_586)
);

O2A1O1Ixp5_ASAP7_75t_L g587 ( 
.A1(n_489),
.A2(n_499),
.B(n_526),
.C(n_488),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_521),
.A2(n_528),
.B1(n_489),
.B2(n_492),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_504),
.A2(n_510),
.B(n_490),
.Y(n_589)
);

A2O1A1Ixp33_ASAP7_75t_L g590 ( 
.A1(n_499),
.A2(n_488),
.B(n_518),
.C(n_517),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_508),
.B(n_502),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_460),
.A2(n_516),
.B1(n_512),
.B2(n_511),
.Y(n_592)
);

CKINVDCx11_ASAP7_75t_R g593 ( 
.A(n_542),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_538),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_535),
.B(n_505),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_560),
.B(n_493),
.Y(n_596)
);

AO31x2_ASAP7_75t_L g597 ( 
.A1(n_575),
.A2(n_519),
.A3(n_503),
.B(n_513),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_538),
.Y(n_598)
);

AOI221x1_ASAP7_75t_L g599 ( 
.A1(n_582),
.A2(n_503),
.B1(n_513),
.B2(n_519),
.C(n_588),
.Y(n_599)
);

O2A1O1Ixp5_ASAP7_75t_L g600 ( 
.A1(n_587),
.A2(n_588),
.B(n_570),
.C(n_574),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_576),
.A2(n_544),
.B(n_536),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_SL g602 ( 
.A(n_577),
.B(n_573),
.C(n_585),
.Y(n_602)
);

A2O1A1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_539),
.A2(n_557),
.B(n_561),
.C(n_546),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_571),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_538),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_548),
.A2(n_554),
.B1(n_541),
.B2(n_547),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_558),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_569),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_546),
.A2(n_584),
.B1(n_562),
.B2(n_534),
.Y(n_609)
);

NOR2x1_ASAP7_75t_R g610 ( 
.A(n_591),
.B(n_540),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_555),
.B(n_572),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_549),
.B(n_563),
.Y(n_612)
);

AO31x2_ASAP7_75t_L g613 ( 
.A1(n_592),
.A2(n_568),
.A3(n_583),
.B(n_580),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_556),
.B(n_559),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_552),
.Y(n_615)
);

INVx3_ASAP7_75t_SL g616 ( 
.A(n_549),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_566),
.B(n_564),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_545),
.A2(n_589),
.B(n_578),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_586),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_581),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_567),
.Y(n_621)
);

A2O1A1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_579),
.A2(n_536),
.B(n_539),
.C(n_557),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_293),
.C(n_500),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_542),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_542),
.A2(n_498),
.B1(n_494),
.B2(n_349),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_542),
.B(n_494),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_537),
.B(n_497),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_552),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_553),
.A2(n_576),
.B(n_484),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_543),
.A2(n_349),
.B1(n_472),
.B2(n_456),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_542),
.B(n_494),
.Y(n_631)
);

AO31x2_ASAP7_75t_L g632 ( 
.A1(n_550),
.A2(n_553),
.A3(n_575),
.B(n_565),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_537),
.B(n_497),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_542),
.B(n_494),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_539),
.A2(n_546),
.B(n_541),
.C(n_551),
.Y(n_635)
);

OAI221xp5_ASAP7_75t_L g636 ( 
.A1(n_557),
.A2(n_495),
.B1(n_354),
.B2(n_360),
.C(n_546),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_539),
.A2(n_546),
.B(n_541),
.C(n_551),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_537),
.B(n_497),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_542),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_539),
.A2(n_546),
.B(n_541),
.C(n_551),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_536),
.A2(n_539),
.B(n_557),
.C(n_349),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_543),
.A2(n_349),
.B1(n_472),
.B2(n_456),
.Y(n_642)
);

BUFx4f_ASAP7_75t_SL g643 ( 
.A(n_542),
.Y(n_643)
);

AO31x2_ASAP7_75t_L g644 ( 
.A1(n_550),
.A2(n_553),
.A3(n_575),
.B(n_565),
.Y(n_644)
);

OAI221xp5_ASAP7_75t_SL g645 ( 
.A1(n_546),
.A2(n_472),
.B1(n_465),
.B2(n_495),
.C(n_376),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_542),
.B(n_494),
.Y(n_646)
);

INVx6_ASAP7_75t_L g647 ( 
.A(n_560),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_553),
.A2(n_576),
.B(n_484),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_542),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_542),
.A2(n_298),
.B1(n_366),
.B2(n_349),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_542),
.Y(n_651)
);

AOI221xp5_ASAP7_75t_SL g652 ( 
.A1(n_541),
.A2(n_551),
.B1(n_472),
.B2(n_539),
.C(n_532),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_537),
.B(n_497),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_552),
.Y(n_654)
);

O2A1O1Ixp5_ASAP7_75t_L g655 ( 
.A1(n_587),
.A2(n_550),
.B(n_553),
.C(n_588),
.Y(n_655)
);

CKINVDCx11_ASAP7_75t_R g656 ( 
.A(n_542),
.Y(n_656)
);

O2A1O1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_539),
.A2(n_546),
.B(n_541),
.C(n_551),
.Y(n_657)
);

O2A1O1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_539),
.A2(n_546),
.B(n_541),
.C(n_551),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_542),
.A2(n_498),
.B1(n_494),
.B2(n_349),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_542),
.A2(n_298),
.B1(n_426),
.B2(n_437),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_537),
.B(n_535),
.Y(n_661)
);

AOI221x1_ASAP7_75t_L g662 ( 
.A1(n_553),
.A2(n_582),
.B1(n_588),
.B2(n_590),
.C(n_476),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_539),
.A2(n_546),
.B(n_541),
.C(n_551),
.Y(n_663)
);

OAI221xp5_ASAP7_75t_L g664 ( 
.A1(n_557),
.A2(n_495),
.B1(n_354),
.B2(n_360),
.C(n_546),
.Y(n_664)
);

AO31x2_ASAP7_75t_L g665 ( 
.A1(n_550),
.A2(n_553),
.A3(n_575),
.B(n_565),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_537),
.Y(n_666)
);

INVx6_ASAP7_75t_SL g667 ( 
.A(n_538),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_542),
.Y(n_669)
);

AO31x2_ASAP7_75t_L g670 ( 
.A1(n_550),
.A2(n_553),
.A3(n_575),
.B(n_565),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_615),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_652),
.B(n_614),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_617),
.B(n_635),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_643),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_650),
.B(n_645),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_637),
.B(n_640),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_636),
.A2(n_664),
.B1(n_611),
.B2(n_630),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_649),
.Y(n_678)
);

OA21x2_ASAP7_75t_L g679 ( 
.A1(n_662),
.A2(n_599),
.B(n_655),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_642),
.A2(n_609),
.B1(n_612),
.B2(n_634),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_657),
.A2(n_658),
.B1(n_663),
.B2(n_620),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_638),
.B(n_653),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_669),
.B(n_639),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_600),
.A2(n_601),
.B(n_629),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_651),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_646),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_623),
.A2(n_595),
.B1(n_624),
.B2(n_606),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_603),
.B(n_641),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_661),
.A2(n_602),
.B1(n_631),
.B2(n_626),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_627),
.B(n_633),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_593),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_615),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_656),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_666),
.B(n_668),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_607),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_SL g696 ( 
.A1(n_594),
.A2(n_660),
.B1(n_598),
.B2(n_605),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_628),
.B(n_654),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_608),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_661),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_616),
.A2(n_667),
.B1(n_621),
.B2(n_604),
.Y(n_700)
);

BUFx12f_ASAP7_75t_L g701 ( 
.A(n_647),
.Y(n_701)
);

BUFx4f_ASAP7_75t_L g702 ( 
.A(n_647),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_619),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_598),
.B(n_625),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_659),
.B(n_610),
.Y(n_705)
);

BUFx8_ASAP7_75t_SL g706 ( 
.A(n_596),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_610),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_632),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_632),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_644),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_644),
.B(n_665),
.Y(n_711)
);

OA21x2_ASAP7_75t_L g712 ( 
.A1(n_597),
.A2(n_613),
.B(n_670),
.Y(n_712)
);

INVx4_ASAP7_75t_SL g713 ( 
.A(n_613),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_635),
.A2(n_640),
.B(n_657),
.C(n_637),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_638),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_638),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_643),
.Y(n_717)
);

AO21x2_ASAP7_75t_L g718 ( 
.A1(n_601),
.A2(n_648),
.B(n_629),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_634),
.B(n_646),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_638),
.B(n_653),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_636),
.A2(n_664),
.B1(n_349),
.B2(n_611),
.Y(n_721)
);

AO31x2_ASAP7_75t_L g722 ( 
.A1(n_662),
.A2(n_599),
.A3(n_618),
.B(n_622),
.Y(n_722)
);

AO31x2_ASAP7_75t_L g723 ( 
.A1(n_662),
.A2(n_599),
.A3(n_618),
.B(n_622),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_638),
.B(n_653),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_673),
.B(n_676),
.Y(n_725)
);

OAI221xp5_ASAP7_75t_L g726 ( 
.A1(n_675),
.A2(n_677),
.B1(n_680),
.B2(n_721),
.C(n_687),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_697),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_718),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_676),
.B(n_714),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_688),
.B(n_681),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_698),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_684),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_694),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_688),
.B(n_711),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_694),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_711),
.B(n_709),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_710),
.B(n_672),
.Y(n_737)
);

AOI33xp33_ASAP7_75t_L g738 ( 
.A1(n_696),
.A2(n_689),
.A3(n_715),
.B1(n_716),
.B2(n_720),
.B3(n_724),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_713),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_722),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_690),
.B(n_682),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_671),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_682),
.B(n_686),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_722),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_697),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_708),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_692),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_723),
.B(n_699),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_748),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_734),
.B(n_712),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_746),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_732),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_730),
.B(n_725),
.Y(n_753)
);

INVx5_ASAP7_75t_L g754 ( 
.A(n_747),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_739),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_739),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_736),
.B(n_679),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_739),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_729),
.B(n_679),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_736),
.B(n_704),
.Y(n_760)
);

NOR2x1p5_ASAP7_75t_L g761 ( 
.A(n_727),
.B(n_707),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_738),
.A2(n_726),
.B(n_733),
.C(n_735),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_737),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_733),
.B(n_705),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_756),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_750),
.B(n_736),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_752),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_749),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_753),
.B(n_740),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_749),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_754),
.B(n_756),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_751),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_750),
.B(n_737),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_750),
.B(n_737),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_754),
.B(n_738),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_750),
.B(n_744),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_773),
.B(n_763),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_772),
.Y(n_778)
);

NAND2x1_ASAP7_75t_SL g779 ( 
.A(n_772),
.B(n_756),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_773),
.B(n_763),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_766),
.B(n_757),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_769),
.B(n_759),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_774),
.B(n_763),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_768),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_765),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_766),
.B(n_757),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_768),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_771),
.Y(n_788)
);

AO22x1_ASAP7_75t_L g789 ( 
.A1(n_765),
.A2(n_756),
.B1(n_755),
.B2(n_758),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_774),
.B(n_760),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_787),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_787),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_779),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_790),
.B(n_770),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_779),
.A2(n_761),
.B(n_745),
.C(n_727),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_781),
.B(n_776),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_781),
.B(n_776),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_784),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_782),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_789),
.B(n_756),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_788),
.B(n_776),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_782),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_801),
.A2(n_775),
.B1(n_788),
.B2(n_777),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_802),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_795),
.A2(n_762),
.B(n_741),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_802),
.B(n_778),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_796),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_799),
.B(n_786),
.Y(n_808)
);

OA21x2_ASAP7_75t_L g809 ( 
.A1(n_791),
.A2(n_785),
.B(n_767),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_798),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_796),
.B(n_786),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_798),
.B(n_731),
.C(n_762),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_793),
.B(n_756),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_793),
.A2(n_761),
.B(n_745),
.C(n_727),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_810),
.Y(n_815)
);

OAI311xp33_ASAP7_75t_L g816 ( 
.A1(n_805),
.A2(n_726),
.A3(n_764),
.B1(n_731),
.C1(n_700),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_811),
.B(n_797),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_806),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_SL g819 ( 
.A1(n_814),
.A2(n_801),
.B(n_741),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_814),
.A2(n_800),
.B1(n_801),
.B2(n_797),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_807),
.Y(n_821)
);

OAI21xp33_ASAP7_75t_SL g822 ( 
.A1(n_817),
.A2(n_813),
.B(n_811),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_819),
.A2(n_812),
.B1(n_803),
.B2(n_804),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_821),
.A2(n_813),
.B1(n_800),
.B2(n_799),
.Y(n_824)
);

AOI221xp5_ASAP7_75t_L g825 ( 
.A1(n_816),
.A2(n_685),
.B1(n_794),
.B2(n_808),
.C(n_792),
.Y(n_825)
);

AOI222xp33_ASAP7_75t_L g826 ( 
.A1(n_820),
.A2(n_743),
.B1(n_764),
.B2(n_791),
.C1(n_691),
.C2(n_783),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_818),
.A2(n_800),
.B(n_789),
.Y(n_827)
);

OAI221xp5_ASAP7_75t_L g828 ( 
.A1(n_822),
.A2(n_818),
.B1(n_800),
.B2(n_815),
.C(n_809),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_823),
.B(n_817),
.Y(n_829)
);

AOI221xp5_ASAP7_75t_L g830 ( 
.A1(n_827),
.A2(n_678),
.B1(n_743),
.B2(n_719),
.C(n_683),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_824),
.B(n_809),
.Y(n_831)
);

NOR3xp33_ASAP7_75t_L g832 ( 
.A(n_828),
.B(n_830),
.C(n_674),
.Y(n_832)
);

XNOR2xp5_ASAP7_75t_L g833 ( 
.A(n_829),
.B(n_693),
.Y(n_833)
);

NOR3xp33_ASAP7_75t_L g834 ( 
.A(n_831),
.B(n_717),
.C(n_695),
.Y(n_834)
);

NOR5xp2_ASAP7_75t_L g835 ( 
.A(n_828),
.B(n_826),
.C(n_825),
.D(n_742),
.E(n_728),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_833),
.B(n_809),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_834),
.B(n_780),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_836),
.B(n_832),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_837),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_839),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_840),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_838),
.B(n_702),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_842),
.A2(n_701),
.B(n_706),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_843),
.A2(n_835),
.B1(n_702),
.B2(n_703),
.Y(n_844)
);


endmodule