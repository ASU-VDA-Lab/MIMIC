module real_jpeg_2571_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_SL g8 ( 
.A(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_0),
.B(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_0),
.B(n_29),
.Y(n_28)
);

AOI322xp5_ASAP7_75t_L g6 ( 
.A1(n_1),
.A2(n_7),
.A3(n_18),
.B1(n_20),
.B2(n_22),
.C1(n_27),
.C2(n_30),
.Y(n_6)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

OR2x4_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

AO21x2_ASAP7_75t_L g15 ( 
.A1(n_3),
.A2(n_16),
.B(n_17),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_4),
.B(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_12),
.Y(n_11)
);

NAND2x1_ASAP7_75t_SL g13 ( 
.A(n_5),
.B(n_12),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_9),
.B(n_14),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_8),
.B(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_8),
.B(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_13),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_14),
.B(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_19),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);


endmodule