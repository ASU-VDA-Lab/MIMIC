module real_aes_17349_n_361 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_361);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_361;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1893;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_1883;
wire n_608;
wire n_760;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1632;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1638;
wire n_495;
wire n_1078;
wire n_1072;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1457;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1647;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g802 ( .A(n_0), .Y(n_802) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1), .Y(n_1621) );
OAI211xp5_ASAP7_75t_L g1420 ( .A1(n_2), .A2(n_465), .B(n_1417), .C(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1434 ( .A(n_2), .Y(n_1434) );
INVx1_ASAP7_75t_L g377 ( .A(n_3), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_3), .B(n_387), .Y(n_501) );
AND2x2_ASAP7_75t_L g576 ( .A(n_3), .B(n_425), .Y(n_576) );
AND2x2_ASAP7_75t_L g593 ( .A(n_3), .B(n_266), .Y(n_593) );
OAI211xp5_ASAP7_75t_SL g828 ( .A1(n_4), .A2(n_403), .B(n_526), .C(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g843 ( .A(n_4), .Y(n_843) );
INVx1_ASAP7_75t_L g876 ( .A(n_5), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g1622 ( .A1(n_6), .A2(n_276), .B1(n_1623), .B2(n_1624), .Y(n_1622) );
OAI211xp5_ASAP7_75t_L g1626 ( .A1(n_6), .A2(n_1627), .B(n_1628), .C(n_1632), .Y(n_1626) );
INVx1_ASAP7_75t_L g1248 ( .A(n_7), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g1356 ( .A1(n_8), .A2(n_293), .B1(n_784), .B2(n_1306), .Y(n_1356) );
OAI22xp33_ASAP7_75t_L g1363 ( .A1(n_8), .A2(n_293), .B1(n_769), .B2(n_770), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1592 ( .A1(n_9), .A2(n_75), .B1(n_662), .B2(n_663), .Y(n_1592) );
AOI22xp33_ASAP7_75t_L g1603 ( .A1(n_9), .A2(n_231), .B1(n_1313), .B2(n_1327), .Y(n_1603) );
INVx1_ASAP7_75t_L g1884 ( .A(n_10), .Y(n_1884) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_11), .A2(n_79), .B1(n_659), .B2(n_1246), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_11), .A2(n_23), .B1(n_942), .B2(n_1264), .C(n_1266), .Y(n_1263) );
INVx1_ASAP7_75t_L g1485 ( .A(n_12), .Y(n_1485) );
OAI22xp5_ASAP7_75t_L g1904 ( .A1(n_13), .A2(n_48), .B1(n_1302), .B2(n_1905), .Y(n_1904) );
OAI22xp5_ASAP7_75t_L g1913 ( .A1(n_13), .A2(n_48), .B1(n_996), .B2(n_1914), .Y(n_1913) );
AOI22xp33_ASAP7_75t_L g1615 ( .A1(n_14), .A2(n_306), .B1(n_662), .B2(n_1230), .Y(n_1615) );
AOI22xp33_ASAP7_75t_L g1635 ( .A1(n_14), .A2(n_353), .B1(n_942), .B2(n_1636), .Y(n_1635) );
AOI22xp5_ASAP7_75t_L g1669 ( .A1(n_15), .A2(n_222), .B1(n_1656), .B2(n_1670), .Y(n_1669) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_16), .A2(n_28), .B1(n_1110), .B2(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1179 ( .A(n_16), .Y(n_1179) );
OAI211xp5_ASAP7_75t_L g1464 ( .A1(n_17), .A2(n_465), .B(n_1465), .C(n_1466), .Y(n_1464) );
INVx1_ASAP7_75t_L g1473 ( .A(n_17), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g1690 ( .A1(n_18), .A2(n_98), .B1(n_1656), .B2(n_1660), .Y(n_1690) );
AOI22xp33_ASAP7_75t_L g1753 ( .A1(n_19), .A2(n_351), .B1(n_1663), .B2(n_1666), .Y(n_1753) );
INVx1_ASAP7_75t_L g1295 ( .A(n_20), .Y(n_1295) );
OAI22xp33_ASAP7_75t_L g1552 ( .A1(n_21), .A2(n_173), .B1(n_1553), .B2(n_1554), .Y(n_1552) );
OAI22xp33_ASAP7_75t_L g1556 ( .A1(n_21), .A2(n_173), .B1(n_379), .B2(n_756), .Y(n_1556) );
CKINVDCx5p33_ASAP7_75t_R g722 ( .A(n_22), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g1255 ( .A1(n_23), .A2(n_250), .B1(n_660), .B2(n_1143), .Y(n_1255) );
INVx1_ASAP7_75t_L g1451 ( .A(n_24), .Y(n_1451) );
INVx2_ASAP7_75t_L g453 ( .A(n_25), .Y(n_453) );
INVx1_ASAP7_75t_L g639 ( .A(n_26), .Y(n_639) );
INVx1_ASAP7_75t_L g807 ( .A(n_27), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_28), .A2(n_47), .B1(n_1159), .B2(n_1161), .C(n_1162), .Y(n_1158) );
INVx1_ASAP7_75t_L g1379 ( .A(n_29), .Y(n_1379) );
INVx1_ASAP7_75t_L g1252 ( .A(n_30), .Y(n_1252) );
AOI22xp5_ASAP7_75t_L g1662 ( .A1(n_31), .A2(n_229), .B1(n_1663), .B2(n_1666), .Y(n_1662) );
INVx1_ASAP7_75t_L g1495 ( .A(n_32), .Y(n_1495) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_33), .A2(n_297), .B1(n_445), .B2(n_782), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_33), .A2(n_333), .B1(n_421), .B2(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g1574 ( .A(n_34), .Y(n_1574) );
OA222x2_ASAP7_75t_L g1054 ( .A1(n_35), .A2(n_85), .B1(n_260), .B2(n_1055), .C1(n_1057), .C2(n_1061), .Y(n_1054) );
INVx1_ASAP7_75t_L g1108 ( .A(n_35), .Y(n_1108) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_36), .Y(n_372) );
AND2x2_ASAP7_75t_L g1657 ( .A(n_36), .B(n_370), .Y(n_1657) );
AOI22xp33_ASAP7_75t_L g1751 ( .A1(n_37), .A2(n_209), .B1(n_1656), .B2(n_1752), .Y(n_1751) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_38), .A2(n_339), .B1(n_574), .B2(n_943), .Y(n_1201) );
INVxp67_ASAP7_75t_SL g1218 ( .A(n_38), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1704 ( .A1(n_39), .A2(n_219), .B1(n_1656), .B2(n_1660), .Y(n_1704) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_40), .A2(n_225), .B1(n_662), .B2(n_973), .Y(n_1144) );
INVx1_ASAP7_75t_L g1164 ( .A(n_40), .Y(n_1164) );
INVx1_ASAP7_75t_L g1885 ( .A(n_41), .Y(n_1885) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_42), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_43), .A2(n_285), .B1(n_996), .B2(n_1298), .Y(n_1297) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_43), .A2(n_192), .B1(n_445), .B2(n_1306), .Y(n_1305) );
OAI22xp33_ASAP7_75t_L g1349 ( .A1(n_44), .A2(n_191), .B1(n_774), .B2(n_1034), .Y(n_1349) );
OAI22xp33_ASAP7_75t_L g1364 ( .A1(n_44), .A2(n_191), .B1(n_379), .B2(n_433), .Y(n_1364) );
XNOR2xp5_ASAP7_75t_L g1440 ( .A(n_45), .B(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g1003 ( .A(n_46), .Y(n_1003) );
AOI22xp33_ASAP7_75t_SL g1148 ( .A1(n_47), .A2(n_329), .B1(n_676), .B2(n_1143), .Y(n_1148) );
INVxp67_ASAP7_75t_SL g1251 ( .A(n_49), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_49), .A2(n_181), .B1(n_615), .B2(n_1272), .Y(n_1271) );
AOI22xp33_ASAP7_75t_SL g1309 ( .A1(n_50), .A2(n_129), .B1(n_1310), .B2(n_1311), .Y(n_1309) );
AOI22xp33_ASAP7_75t_SL g1338 ( .A1(n_50), .A2(n_265), .B1(n_1220), .B2(n_1333), .Y(n_1338) );
INVx1_ASAP7_75t_L g1491 ( .A(n_51), .Y(n_1491) );
INVx1_ASAP7_75t_L g1010 ( .A(n_52), .Y(n_1010) );
INVx1_ASAP7_75t_L g1534 ( .A(n_53), .Y(n_1534) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_54), .A2(n_399), .B(n_403), .C(n_408), .Y(n_398) );
INVx1_ASAP7_75t_L g474 ( .A(n_54), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g1078 ( .A(n_55), .Y(n_1078) );
INVx1_ASAP7_75t_L g1259 ( .A(n_56), .Y(n_1259) );
INVx1_ASAP7_75t_L g870 ( .A(n_57), .Y(n_870) );
AOI22xp33_ASAP7_75t_SL g1206 ( .A1(n_58), .A2(n_275), .B1(n_943), .B2(n_1207), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_58), .A2(n_254), .B1(n_1099), .B2(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1549 ( .A(n_59), .Y(n_1549) );
AOI22xp5_ASAP7_75t_L g1677 ( .A1(n_60), .A2(n_180), .B1(n_1656), .B2(n_1660), .Y(n_1677) );
CKINVDCx5p33_ASAP7_75t_R g1250 ( .A(n_61), .Y(n_1250) );
INVx1_ASAP7_75t_L g1281 ( .A(n_62), .Y(n_1281) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_63), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_64), .A2(n_76), .B1(n_671), .B2(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1163 ( .A(n_64), .Y(n_1163) );
INVx1_ASAP7_75t_L g513 ( .A(n_65), .Y(n_513) );
INVx1_ASAP7_75t_L g1530 ( .A(n_66), .Y(n_1530) );
OAI22xp33_ASAP7_75t_SL g1197 ( .A1(n_67), .A2(n_263), .B1(n_524), .B2(n_1077), .Y(n_1197) );
INVx1_ASAP7_75t_L g1234 ( .A(n_67), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_68), .A2(n_108), .B1(n_586), .B2(n_590), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_68), .A2(n_243), .B1(n_662), .B2(n_663), .Y(n_661) );
XNOR2xp5_ASAP7_75t_L g1480 ( .A(n_69), .B(n_1481), .Y(n_1480) );
AOI21xp33_ASAP7_75t_L g954 ( .A1(n_70), .A2(n_955), .B(n_956), .Y(n_954) );
AOI221xp5_ASAP7_75t_L g977 ( .A1(n_70), .A2(n_283), .B1(n_973), .B2(n_978), .C(n_980), .Y(n_977) );
CKINVDCx5p33_ASAP7_75t_R g1135 ( .A(n_71), .Y(n_1135) );
XOR2x2_ASAP7_75t_L g568 ( .A(n_72), .B(n_569), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g755 ( .A1(n_73), .A2(n_121), .B1(n_379), .B2(n_756), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g773 ( .A1(n_73), .A2(n_121), .B1(n_445), .B2(n_774), .Y(n_773) );
OAI222xp33_ASAP7_75t_L g916 ( .A1(n_74), .A2(n_83), .B1(n_89), .B2(n_645), .C1(n_917), .C2(n_923), .Y(n_916) );
AOI22xp33_ASAP7_75t_SL g1600 ( .A1(n_75), .A2(n_104), .B1(n_1322), .B2(n_1601), .Y(n_1600) );
INVx1_ASAP7_75t_L g1183 ( .A(n_76), .Y(n_1183) );
INVx1_ASAP7_75t_L g1514 ( .A(n_77), .Y(n_1514) );
OAI211xp5_ASAP7_75t_L g1520 ( .A1(n_77), .A2(n_909), .B(n_1521), .C(n_1523), .Y(n_1520) );
OAI22xp33_ASAP7_75t_L g1607 ( .A1(n_78), .A2(n_316), .B1(n_693), .B2(n_922), .Y(n_1607) );
INVx1_ASAP7_75t_L g1629 ( .A(n_78), .Y(n_1629) );
INVx1_ASAP7_75t_L g1280 ( .A(n_79), .Y(n_1280) );
INVx1_ASAP7_75t_L g873 ( .A(n_80), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g997 ( .A1(n_81), .A2(n_84), .B1(n_998), .B2(n_999), .Y(n_997) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_81), .A2(n_84), .B1(n_484), .B2(n_1044), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g935 ( .A(n_82), .Y(n_935) );
OAI221xp5_ASAP7_75t_L g1092 ( .A1(n_85), .A2(n_204), .B1(n_1093), .B2(n_1095), .C(n_1097), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_86), .A2(n_311), .B1(n_429), .B2(n_615), .Y(n_1172) );
INVx1_ASAP7_75t_L g1185 ( .A(n_86), .Y(n_1185) );
INVx1_ASAP7_75t_L g1068 ( .A(n_87), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_87), .A2(n_141), .B1(n_665), .B2(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1019 ( .A(n_88), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_89), .A2(n_357), .B1(n_967), .B2(n_969), .Y(n_966) );
INVx1_ASAP7_75t_L g1380 ( .A(n_90), .Y(n_1380) );
INVx1_ASAP7_75t_L g795 ( .A(n_91), .Y(n_795) );
INVx1_ASAP7_75t_L g830 ( .A(n_92), .Y(n_830) );
INVx1_ASAP7_75t_L g1573 ( .A(n_93), .Y(n_1573) );
AOI22xp33_ASAP7_75t_SL g1594 ( .A1(n_94), .A2(n_178), .B1(n_1143), .B2(n_1331), .Y(n_1594) );
AOI22xp33_ASAP7_75t_L g1597 ( .A1(n_94), .A2(n_240), .B1(n_1313), .B2(n_1598), .Y(n_1597) );
XOR2x2_ASAP7_75t_L g851 ( .A(n_95), .B(n_852), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_96), .A2(n_170), .B1(n_958), .B2(n_959), .Y(n_957) );
INVx1_ASAP7_75t_L g975 ( .A(n_96), .Y(n_975) );
INVx1_ASAP7_75t_L g1489 ( .A(n_97), .Y(n_1489) );
CKINVDCx5p33_ASAP7_75t_R g1258 ( .A(n_99), .Y(n_1258) );
AOI22xp33_ASAP7_75t_SL g1616 ( .A1(n_100), .A2(n_267), .B1(n_1127), .B2(n_1225), .Y(n_1616) );
AOI221xp5_ASAP7_75t_L g1633 ( .A1(n_100), .A2(n_318), .B1(n_579), .B2(n_584), .C(n_1634), .Y(n_1633) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_101), .A2(n_334), .B1(n_663), .B2(n_1146), .Y(n_1254) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_101), .A2(n_221), .B1(n_943), .B2(n_1161), .C(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1531 ( .A(n_102), .Y(n_1531) );
AOI22xp5_ASAP7_75t_L g1681 ( .A1(n_103), .A2(n_228), .B1(n_1663), .B2(n_1666), .Y(n_1681) );
AOI22xp33_ASAP7_75t_L g1591 ( .A1(n_104), .A2(n_231), .B1(n_662), .B2(n_663), .Y(n_1591) );
OAI22xp33_ASAP7_75t_L g1419 ( .A1(n_105), .A2(n_166), .B1(n_447), .B2(n_774), .Y(n_1419) );
OAI22xp33_ASAP7_75t_L g1429 ( .A1(n_105), .A2(n_166), .B1(n_379), .B2(n_433), .Y(n_1429) );
INVx1_ASAP7_75t_L g1187 ( .A(n_106), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_107), .A2(n_155), .B1(n_995), .B2(n_996), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_107), .A2(n_155), .B1(n_838), .B2(n_1034), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_108), .A2(n_128), .B1(n_668), .B2(n_671), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_109), .A2(n_190), .B1(n_484), .B2(n_774), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g1474 ( .A1(n_109), .A2(n_230), .B1(n_1436), .B2(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1397 ( .A(n_110), .Y(n_1397) );
INVx1_ASAP7_75t_L g370 ( .A(n_111), .Y(n_370) );
INVx1_ASAP7_75t_L g1488 ( .A(n_112), .Y(n_1488) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_113), .A2(n_179), .B1(n_641), .B2(n_645), .Y(n_640) );
XOR2x2_ASAP7_75t_L g1346 ( .A(n_114), .B(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1448 ( .A(n_115), .Y(n_1448) );
INVx1_ASAP7_75t_L g858 ( .A(n_116), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_117), .A2(n_358), .B1(n_421), .B2(n_426), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_117), .A2(n_127), .B1(n_445), .B2(n_454), .Y(n_444) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_118), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_118), .A2(n_290), .B1(n_659), .B2(n_676), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g1196 ( .A1(n_119), .A2(n_159), .B1(n_1069), .B2(n_1070), .Y(n_1196) );
NOR2xp33_ASAP7_75t_L g1238 ( .A(n_119), .B(n_454), .Y(n_1238) );
INVx1_ASAP7_75t_L g813 ( .A(n_120), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_122), .Y(n_1154) );
INVx1_ASAP7_75t_L g809 ( .A(n_123), .Y(n_809) );
INVx1_ASAP7_75t_L g1408 ( .A(n_124), .Y(n_1408) );
INVx1_ASAP7_75t_L g811 ( .A(n_125), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_126), .A2(n_138), .B1(n_423), .B2(n_426), .Y(n_833) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_126), .A2(n_138), .B1(n_782), .B2(n_845), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g432 ( .A1(n_127), .A2(n_332), .B1(n_379), .B2(n_433), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_128), .A2(n_243), .B1(n_582), .B2(n_620), .C(n_622), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_129), .A2(n_245), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
AOI22xp5_ASAP7_75t_L g1686 ( .A1(n_130), .A2(n_330), .B1(n_1663), .B2(n_1666), .Y(n_1686) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_131), .A2(n_353), .B1(n_662), .B2(n_1614), .Y(n_1613) );
AOI21xp33_ASAP7_75t_L g1642 ( .A1(n_131), .A2(n_622), .B(n_1643), .Y(n_1642) );
INVx1_ASAP7_75t_L g1376 ( .A(n_132), .Y(n_1376) );
INVx1_ASAP7_75t_L g832 ( .A(n_133), .Y(n_832) );
OAI211xp5_ASAP7_75t_L g839 ( .A1(n_133), .A2(n_465), .B(n_840), .C(n_842), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_134), .A2(n_333), .B1(n_478), .B2(n_484), .Y(n_897) );
OAI22xp33_ASAP7_75t_L g899 ( .A1(n_134), .A2(n_297), .B1(n_379), .B2(n_756), .Y(n_899) );
INVx1_ASAP7_75t_L g798 ( .A(n_135), .Y(n_798) );
INVx1_ASAP7_75t_L g1533 ( .A(n_136), .Y(n_1533) );
INVx1_ASAP7_75t_L g1571 ( .A(n_137), .Y(n_1571) );
INVx1_ASAP7_75t_L g1910 ( .A(n_139), .Y(n_1910) );
OAI211xp5_ASAP7_75t_L g1916 ( .A1(n_139), .A2(n_520), .B(n_1431), .C(n_1917), .Y(n_1916) );
OAI211xp5_ASAP7_75t_L g1547 ( .A1(n_140), .A2(n_1037), .B(n_1465), .C(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1560 ( .A(n_140), .Y(n_1560) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_141), .A2(n_188), .B1(n_586), .B2(n_590), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g1655 ( .A1(n_142), .A2(n_234), .B1(n_1656), .B2(n_1660), .Y(n_1655) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_143), .A2(n_290), .B1(n_579), .B2(n_580), .C(n_584), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_143), .A2(n_248), .B1(n_657), .B2(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g1540 ( .A(n_144), .Y(n_1540) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_145), .A2(n_204), .B1(n_642), .B2(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1109 ( .A(n_145), .Y(n_1109) );
INVx1_ASAP7_75t_L g1399 ( .A(n_146), .Y(n_1399) );
INVx1_ASAP7_75t_L g1401 ( .A(n_147), .Y(n_1401) );
OAI211xp5_ASAP7_75t_L g757 ( .A1(n_148), .A2(n_403), .B(n_758), .C(n_762), .Y(n_757) );
INVx1_ASAP7_75t_L g780 ( .A(n_148), .Y(n_780) );
INVx1_ASAP7_75t_L g1890 ( .A(n_149), .Y(n_1890) );
OAI22xp33_ASAP7_75t_L g834 ( .A1(n_150), .A2(n_255), .B1(n_433), .B2(n_835), .Y(n_834) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_150), .A2(n_255), .B1(n_447), .B2(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g1013 ( .A(n_151), .Y(n_1013) );
INVx1_ASAP7_75t_L g1455 ( .A(n_152), .Y(n_1455) );
AOI22xp5_ASAP7_75t_L g1671 ( .A1(n_153), .A2(n_244), .B1(n_1663), .B2(n_1666), .Y(n_1671) );
INVx1_ASAP7_75t_L g1619 ( .A(n_154), .Y(n_1619) );
OAI221xp5_ASAP7_75t_L g1637 ( .A1(n_154), .A2(n_206), .B1(n_1638), .B2(n_1639), .C(n_1640), .Y(n_1637) );
OAI221xp5_ASAP7_75t_L g1210 ( .A1(n_156), .A2(n_342), .B1(n_744), .B2(n_1211), .C(n_1213), .Y(n_1210) );
INVx1_ASAP7_75t_L g1231 ( .A(n_156), .Y(n_1231) );
INVx1_ASAP7_75t_L g1199 ( .A(n_157), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_157), .A2(n_275), .B1(n_1099), .B2(n_1225), .Y(n_1224) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_158), .Y(n_1203) );
INVx1_ASAP7_75t_L g1233 ( .A(n_159), .Y(n_1233) );
INVx1_ASAP7_75t_L g1294 ( .A(n_160), .Y(n_1294) );
OAI211xp5_ASAP7_75t_L g1303 ( .A1(n_160), .A2(n_458), .B(n_1037), .C(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1355 ( .A(n_161), .Y(n_1355) );
OAI211xp5_ASAP7_75t_L g1358 ( .A1(n_161), .A2(n_1359), .B(n_1360), .C(n_1361), .Y(n_1358) );
OAI211xp5_ASAP7_75t_L g893 ( .A1(n_162), .A2(n_458), .B(n_465), .C(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g908 ( .A(n_162), .Y(n_908) );
INVx1_ASAP7_75t_L g1468 ( .A(n_163), .Y(n_1468) );
OAI211xp5_ASAP7_75t_SL g1471 ( .A1(n_163), .A2(n_403), .B(n_905), .C(n_1472), .Y(n_1471) );
OAI22xp33_ASAP7_75t_L g1515 ( .A1(n_164), .A2(n_269), .B1(n_445), .B2(n_1516), .Y(n_1515) );
OAI22xp5_ASAP7_75t_L g1518 ( .A1(n_164), .A2(n_269), .B1(n_996), .B2(n_1298), .Y(n_1518) );
OAI22xp5_ASAP7_75t_L g1463 ( .A1(n_165), .A2(n_230), .B1(n_445), .B2(n_782), .Y(n_1463) );
OAI22xp33_ASAP7_75t_L g1476 ( .A1(n_165), .A2(n_190), .B1(n_379), .B2(n_756), .Y(n_1476) );
INVx1_ASAP7_75t_L g1373 ( .A(n_167), .Y(n_1373) );
INVx1_ASAP7_75t_L g1486 ( .A(n_168), .Y(n_1486) );
INVx1_ASAP7_75t_L g1492 ( .A(n_169), .Y(n_1492) );
INVxp67_ASAP7_75t_SL g981 ( .A(n_170), .Y(n_981) );
INVx1_ASAP7_75t_L g1422 ( .A(n_171), .Y(n_1422) );
INVx1_ASAP7_75t_L g1537 ( .A(n_172), .Y(n_1537) );
OAI22xp33_ASAP7_75t_L g1508 ( .A1(n_174), .A2(n_200), .B1(n_484), .B2(n_1509), .Y(n_1508) );
OAI22xp33_ASAP7_75t_L g1519 ( .A1(n_174), .A2(n_200), .B1(n_421), .B2(n_901), .Y(n_1519) );
XNOR2xp5_ASAP7_75t_L g1565 ( .A(n_175), .B(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1377 ( .A(n_176), .Y(n_1377) );
INVx1_ASAP7_75t_L g1403 ( .A(n_177), .Y(n_1403) );
AOI22xp33_ASAP7_75t_SL g1602 ( .A1(n_178), .A2(n_315), .B1(n_1314), .B2(n_1601), .Y(n_1602) );
OAI211xp5_ASAP7_75t_L g571 ( .A1(n_179), .A2(n_572), .B(n_577), .C(n_594), .Y(n_571) );
XOR2x2_ASAP7_75t_L g1879 ( .A(n_180), .B(n_1880), .Y(n_1879) );
AOI22xp33_ASAP7_75t_L g1923 ( .A1(n_180), .A2(n_1924), .B1(n_1927), .B2(n_1930), .Y(n_1923) );
INVxp67_ASAP7_75t_SL g1261 ( .A(n_181), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g1076 ( .A(n_182), .Y(n_1076) );
INVx1_ASAP7_75t_L g1909 ( .A(n_183), .Y(n_1909) );
INVx1_ASAP7_75t_L g1893 ( .A(n_184), .Y(n_1893) );
INVx1_ASAP7_75t_L g1190 ( .A(n_185), .Y(n_1190) );
INVx1_ASAP7_75t_L g507 ( .A(n_186), .Y(n_507) );
INVx1_ASAP7_75t_L g1576 ( .A(n_187), .Y(n_1576) );
OAI22xp5_ASAP7_75t_L g1581 ( .A1(n_187), .A2(n_304), .B1(n_1582), .B2(n_1583), .Y(n_1581) );
INVx1_ASAP7_75t_L g1122 ( .A(n_188), .Y(n_1122) );
INVx1_ASAP7_75t_L g409 ( .A(n_189), .Y(n_409) );
INVx1_ASAP7_75t_L g1292 ( .A(n_192), .Y(n_1292) );
OAI22xp33_ASAP7_75t_L g1551 ( .A1(n_193), .A2(n_349), .B1(n_484), .B2(n_782), .Y(n_1551) );
OAI22xp33_ASAP7_75t_L g1557 ( .A1(n_193), .A2(n_349), .B1(n_421), .B2(n_901), .Y(n_1557) );
INVx1_ASAP7_75t_L g1370 ( .A(n_194), .Y(n_1370) );
INVx1_ASAP7_75t_L g953 ( .A(n_195), .Y(n_953) );
AOI221x1_ASAP7_75t_SL g972 ( .A1(n_195), .A2(n_278), .B1(n_668), .B2(n_973), .C(n_974), .Y(n_972) );
AOI221x1_ASAP7_75t_SL g1063 ( .A1(n_196), .A2(n_272), .B1(n_1064), .B2(n_1065), .C(n_1067), .Y(n_1063) );
AOI21xp33_ASAP7_75t_L g1124 ( .A1(n_196), .A2(n_551), .B(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g595 ( .A(n_197), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_197), .A2(n_317), .B1(n_690), .B2(n_693), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g962 ( .A1(n_198), .A2(n_963), .B(n_964), .Y(n_962) );
INVx1_ASAP7_75t_L g982 ( .A(n_198), .Y(n_982) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_199), .A2(n_273), .B1(n_603), .B2(n_607), .C(n_612), .Y(n_602) );
INVx1_ASAP7_75t_L g679 ( .A(n_199), .Y(n_679) );
INVx2_ASAP7_75t_L g1659 ( .A(n_201), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_201), .B(n_307), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_201), .B(n_1665), .Y(n_1667) );
INVx1_ASAP7_75t_L g519 ( .A(n_202), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g1676 ( .A1(n_203), .A2(n_287), .B1(n_1663), .B2(n_1666), .Y(n_1676) );
OAI22xp33_ASAP7_75t_L g1911 ( .A1(n_205), .A2(n_271), .B1(n_845), .B2(n_1306), .Y(n_1911) );
OAI22xp33_ASAP7_75t_L g1919 ( .A1(n_205), .A2(n_271), .B1(n_999), .B2(n_1436), .Y(n_1919) );
INVx1_ASAP7_75t_L g1618 ( .A(n_206), .Y(n_1618) );
INVx1_ASAP7_75t_L g525 ( .A(n_207), .Y(n_525) );
INVx1_ASAP7_75t_L g1296 ( .A(n_208), .Y(n_1296) );
INVx1_ASAP7_75t_L g992 ( .A(n_210), .Y(n_992) );
INVx1_ASAP7_75t_L g1354 ( .A(n_211), .Y(n_1354) );
INVx1_ASAP7_75t_L g895 ( .A(n_212), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g1687 ( .A1(n_213), .A2(n_322), .B1(n_1656), .B2(n_1670), .Y(n_1687) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_214), .Y(n_1072) );
INVx1_ASAP7_75t_L g535 ( .A(n_215), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_216), .A2(n_348), .B1(n_1313), .B2(n_1314), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_216), .A2(n_220), .B1(n_1336), .B2(n_1337), .Y(n_1335) );
OAI211xp5_ASAP7_75t_L g990 ( .A1(n_217), .A2(n_883), .B(n_909), .C(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g1042 ( .A(n_217), .Y(n_1042) );
INVx1_ASAP7_75t_L g1423 ( .A(n_218), .Y(n_1423) );
OAI211xp5_ASAP7_75t_L g1430 ( .A1(n_218), .A2(n_945), .B(n_1431), .C(n_1433), .Y(n_1430) );
XOR2x2_ASAP7_75t_L g703 ( .A(n_219), .B(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g1326 ( .A1(n_220), .A2(n_344), .B1(n_1313), .B2(n_1327), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_221), .A2(n_319), .B1(n_668), .B2(n_671), .Y(n_1244) );
XNOR2xp5_ASAP7_75t_L g395 ( .A(n_222), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g1887 ( .A(n_223), .Y(n_1887) );
INVx1_ASAP7_75t_L g878 ( .A(n_224), .Y(n_878) );
INVx1_ASAP7_75t_L g1181 ( .A(n_225), .Y(n_1181) );
INVx1_ASAP7_75t_L g1888 ( .A(n_226), .Y(n_1888) );
INVx2_ASAP7_75t_L g491 ( .A(n_227), .Y(n_491) );
INVx1_ASAP7_75t_L g563 ( .A(n_227), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_227), .B(n_453), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_232), .A2(n_241), .B1(n_769), .B2(n_770), .Y(n_768) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_232), .A2(n_241), .B1(n_782), .B2(n_784), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_233), .Y(n_717) );
XNOR2xp5_ASAP7_75t_L g1604 ( .A(n_234), .B(n_1605), .Y(n_1604) );
INVx1_ASAP7_75t_L g1467 ( .A(n_235), .Y(n_1467) );
INVx1_ASAP7_75t_L g914 ( .A(n_236), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g1689 ( .A1(n_237), .A2(n_326), .B1(n_1663), .B2(n_1666), .Y(n_1689) );
INVx1_ASAP7_75t_L g538 ( .A(n_238), .Y(n_538) );
INVx1_ASAP7_75t_L g1454 ( .A(n_239), .Y(n_1454) );
AOI22xp33_ASAP7_75t_SL g1588 ( .A1(n_240), .A2(n_315), .B1(n_660), .B2(n_1589), .Y(n_1588) );
BUFx3_ASAP7_75t_L g449 ( .A(n_242), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g1320 ( .A1(n_245), .A2(n_265), .B1(n_1321), .B2(n_1322), .Y(n_1320) );
INVx1_ASAP7_75t_L g1895 ( .A(n_246), .Y(n_1895) );
INVx1_ASAP7_75t_L g1550 ( .A(n_247), .Y(n_1550) );
OAI211xp5_ASAP7_75t_L g1558 ( .A1(n_247), .A2(n_909), .B(n_1521), .C(n_1559), .Y(n_1558) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_248), .Y(n_616) );
OAI22xp5_ASAP7_75t_SL g937 ( .A1(n_249), .A2(n_291), .B1(n_632), .B2(n_644), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_249), .Y(n_948) );
INVx1_ASAP7_75t_L g1279 ( .A(n_250), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1610 ( .A1(n_251), .A2(n_318), .B1(n_660), .B2(n_1611), .Y(n_1610) );
AOI22xp33_ASAP7_75t_L g1644 ( .A1(n_251), .A2(n_267), .B1(n_942), .B2(n_1161), .Y(n_1644) );
INVx1_ASAP7_75t_L g1368 ( .A(n_252), .Y(n_1368) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_253), .Y(n_713) );
AOI21xp33_ASAP7_75t_L g1200 ( .A1(n_254), .A2(n_963), .B(n_964), .Y(n_1200) );
INVx1_ASAP7_75t_L g865 ( .A(n_256), .Y(n_865) );
INVx1_ASAP7_75t_L g1008 ( .A(n_257), .Y(n_1008) );
INVx1_ASAP7_75t_L g1372 ( .A(n_258), .Y(n_1372) );
INVx1_ASAP7_75t_L g1452 ( .A(n_259), .Y(n_1452) );
INVx1_ASAP7_75t_L g1098 ( .A(n_260), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g1682 ( .A1(n_261), .A2(n_277), .B1(n_1656), .B2(n_1660), .Y(n_1682) );
INVx1_ASAP7_75t_L g1494 ( .A(n_262), .Y(n_1494) );
INVx1_ASAP7_75t_L g1237 ( .A(n_263), .Y(n_1237) );
INVx1_ASAP7_75t_L g503 ( .A(n_264), .Y(n_503) );
BUFx3_ASAP7_75t_L g387 ( .A(n_266), .Y(n_387) );
INVx1_ASAP7_75t_L g425 ( .A(n_266), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g1424 ( .A1(n_268), .A2(n_314), .B1(n_1306), .B2(n_1425), .Y(n_1424) );
OAI22xp5_ASAP7_75t_L g1435 ( .A1(n_268), .A2(n_314), .B1(n_1436), .B2(n_1437), .Y(n_1435) );
XNOR2xp5_ASAP7_75t_L g789 ( .A(n_270), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g1121 ( .A(n_272), .Y(n_1121) );
INVx1_ASAP7_75t_L g684 ( .A(n_273), .Y(n_684) );
INVx1_ASAP7_75t_L g1445 ( .A(n_274), .Y(n_1445) );
INVx1_ASAP7_75t_L g1052 ( .A(n_277), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_278), .A2(n_283), .B1(n_958), .B2(n_959), .Y(n_965) );
INVx1_ASAP7_75t_L g1446 ( .A(n_279), .Y(n_1446) );
INVx1_ASAP7_75t_L g805 ( .A(n_280), .Y(n_805) );
INVx1_ASAP7_75t_L g993 ( .A(n_281), .Y(n_993) );
OAI211xp5_ASAP7_75t_L g1036 ( .A1(n_281), .A2(n_546), .B(n_1037), .C(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g859 ( .A(n_282), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_284), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g1301 ( .A1(n_285), .A2(n_360), .B1(n_845), .B2(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1014 ( .A(n_286), .Y(n_1014) );
INVx1_ASAP7_75t_L g1406 ( .A(n_288), .Y(n_1406) );
CKINVDCx5p33_ASAP7_75t_R g1156 ( .A(n_289), .Y(n_1156) );
INVx1_ASAP7_75t_L g941 ( .A(n_291), .Y(n_941) );
INVx1_ASAP7_75t_L g451 ( .A(n_292), .Y(n_451) );
INVx1_ASAP7_75t_L g463 ( .A(n_292), .Y(n_463) );
INVx1_ASAP7_75t_L g1536 ( .A(n_294), .Y(n_1536) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_295), .Y(n_764) );
INVx1_ASAP7_75t_L g861 ( .A(n_296), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_298), .Y(n_715) );
INVx1_ASAP7_75t_L g961 ( .A(n_299), .Y(n_961) );
INVx1_ASAP7_75t_L g1409 ( .A(n_300), .Y(n_1409) );
INVx1_ASAP7_75t_L g1513 ( .A(n_301), .Y(n_1513) );
INVx1_ASAP7_75t_L g1891 ( .A(n_302), .Y(n_1891) );
AOI22xp5_ASAP7_75t_L g986 ( .A1(n_303), .A2(n_987), .B1(n_988), .B2(n_1045), .Y(n_986) );
INVxp67_ASAP7_75t_SL g1045 ( .A(n_303), .Y(n_1045) );
INVx1_ASAP7_75t_L g1577 ( .A(n_304), .Y(n_1577) );
CKINVDCx5p33_ASAP7_75t_R g1150 ( .A(n_305), .Y(n_1150) );
INVxp67_ASAP7_75t_SL g1641 ( .A(n_306), .Y(n_1641) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_307), .B(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g1665 ( .A(n_307), .Y(n_1665) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_308), .Y(n_730) );
OAI211xp5_ASAP7_75t_SL g1510 ( .A1(n_309), .A2(n_1037), .B(n_1511), .C(n_1512), .Y(n_1510) );
INVx1_ASAP7_75t_L g1524 ( .A(n_309), .Y(n_1524) );
INVx1_ASAP7_75t_L g1578 ( .A(n_310), .Y(n_1578) );
INVx1_ASAP7_75t_L g1138 ( .A(n_311), .Y(n_1138) );
OAI211xp5_ASAP7_75t_L g1907 ( .A1(n_312), .A2(n_465), .B(n_983), .C(n_1908), .Y(n_1907) );
INVx1_ASAP7_75t_L g1918 ( .A(n_312), .Y(n_1918) );
XOR2xp5_ASAP7_75t_L g1928 ( .A(n_313), .B(n_1929), .Y(n_1928) );
INVx1_ASAP7_75t_L g1630 ( .A(n_316), .Y(n_1630) );
INVx1_ASAP7_75t_L g598 ( .A(n_317), .Y(n_598) );
INVx1_ASAP7_75t_L g1268 ( .A(n_319), .Y(n_1268) );
INVx1_ASAP7_75t_L g527 ( .A(n_320), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g1705 ( .A1(n_321), .A2(n_354), .B1(n_1663), .B2(n_1666), .Y(n_1705) );
INVx1_ASAP7_75t_L g414 ( .A(n_323), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g457 ( .A1(n_323), .A2(n_458), .B(n_465), .C(n_469), .Y(n_457) );
INVx1_ASAP7_75t_L g1209 ( .A(n_324), .Y(n_1209) );
INVx1_ASAP7_75t_L g767 ( .A(n_325), .Y(n_767) );
OAI211xp5_ASAP7_75t_L g775 ( .A1(n_325), .A2(n_465), .B(n_776), .C(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g1449 ( .A(n_327), .Y(n_1449) );
OAI22xp5_ASAP7_75t_L g1284 ( .A1(n_328), .A2(n_1285), .B1(n_1339), .B2(n_1340), .Y(n_1284) );
INVxp67_ASAP7_75t_SL g1340 ( .A(n_328), .Y(n_1340) );
AOI211xp5_ASAP7_75t_SL g1176 ( .A1(n_329), .A2(n_1177), .B(n_1178), .C(n_1180), .Y(n_1176) );
AOI21xp5_ASAP7_75t_SL g1204 ( .A1(n_331), .A2(n_963), .B(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1217 ( .A(n_331), .Y(n_1217) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_332), .A2(n_358), .B1(n_478), .B2(n_484), .Y(n_477) );
INVx1_ASAP7_75t_L g1267 ( .A(n_334), .Y(n_1267) );
XNOR2xp5_ASAP7_75t_L g1525 ( .A(n_335), .B(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1539 ( .A(n_336), .Y(n_1539) );
INVx1_ASAP7_75t_L g1394 ( .A(n_337), .Y(n_1394) );
XOR2x2_ASAP7_75t_L g1389 ( .A(n_338), .B(n_1390), .Y(n_1389) );
INVxp67_ASAP7_75t_L g1223 ( .A(n_339), .Y(n_1223) );
OAI211xp5_ASAP7_75t_L g1350 ( .A1(n_340), .A2(n_465), .B(n_1351), .C(n_1352), .Y(n_1350) );
INVx1_ASAP7_75t_L g1362 ( .A(n_340), .Y(n_1362) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_341), .Y(n_709) );
INVxp67_ASAP7_75t_SL g1236 ( .A(n_342), .Y(n_1236) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g1332 ( .A1(n_344), .A2(n_348), .B1(n_663), .B2(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1006 ( .A(n_345), .Y(n_1006) );
INVx1_ASAP7_75t_L g1020 ( .A(n_346), .Y(n_1020) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_347), .Y(n_1089) );
INVx1_ASAP7_75t_L g1570 ( .A(n_350), .Y(n_1570) );
INVx1_ASAP7_75t_L g896 ( .A(n_352), .Y(n_896) );
OAI211xp5_ASAP7_75t_L g904 ( .A1(n_352), .A2(n_905), .B(n_906), .C(n_909), .Y(n_904) );
INVx1_ASAP7_75t_L g442 ( .A(n_355), .Y(n_442) );
INVx2_ASAP7_75t_L g500 ( .A(n_355), .Y(n_500) );
INVx1_ASAP7_75t_L g562 ( .A(n_355), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_356), .Y(n_1090) );
INVx1_ASAP7_75t_L g936 ( .A(n_357), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g1140 ( .A(n_359), .Y(n_1140) );
INVx1_ASAP7_75t_L g1290 ( .A(n_360), .Y(n_1290) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_388), .B(n_1647), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx4f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_373), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g1922 ( .A(n_367), .B(n_376), .Y(n_1922) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g1926 ( .A(n_369), .B(n_372), .Y(n_1926) );
INVx1_ASAP7_75t_L g1933 ( .A(n_369), .Y(n_1933) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g1935 ( .A(n_372), .B(n_1933), .Y(n_1935) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g438 ( .A(n_376), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g533 ( .A(n_377), .B(n_387), .Y(n_533) );
AND2x4_ASAP7_75t_L g623 ( .A(n_377), .B(n_386), .Y(n_623) );
INVx1_ASAP7_75t_L g995 ( .A(n_378), .Y(n_995) );
INVxp67_ASAP7_75t_SL g1298 ( .A(n_378), .Y(n_1298) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_378), .A2(n_434), .B1(n_1573), .B2(n_1574), .Y(n_1572) );
AND2x4_ASAP7_75t_SL g1921 ( .A(n_378), .B(n_1922), .Y(n_1921) );
INVx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x6_ASAP7_75t_L g379 ( .A(n_380), .B(n_385), .Y(n_379) );
OR2x6_ASAP7_75t_L g423 ( .A(n_380), .B(n_424), .Y(n_423) );
BUFx4f_ASAP7_75t_L g826 ( .A(n_380), .Y(n_826) );
INVx1_ASAP7_75t_L g889 ( .A(n_380), .Y(n_889) );
INVxp67_ASAP7_75t_L g1396 ( .A(n_380), .Y(n_1396) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx4f_ASAP7_75t_L g506 ( .A(n_381), .Y(n_506) );
INVx3_ASAP7_75t_L g615 ( .A(n_381), .Y(n_615) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NAND2x1_ASAP7_75t_L g402 ( .A(n_383), .B(n_384), .Y(n_402) );
AND2x2_ASAP7_75t_L g407 ( .A(n_383), .B(n_384), .Y(n_407) );
INVx1_ASAP7_75t_L g419 ( .A(n_383), .Y(n_419) );
INVx2_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
AND2x2_ASAP7_75t_L g435 ( .A(n_383), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g518 ( .A(n_383), .Y(n_518) );
BUFx2_ASAP7_75t_L g413 ( .A(n_384), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_384), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g436 ( .A(n_384), .Y(n_436) );
OR2x2_ASAP7_75t_L g517 ( .A(n_384), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g575 ( .A(n_384), .B(n_431), .Y(n_575) );
INVx1_ASAP7_75t_L g589 ( .A(n_384), .Y(n_589) );
OR2x6_ASAP7_75t_L g835 ( .A(n_385), .B(n_615), .Y(n_835) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g405 ( .A(n_386), .Y(n_405) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g412 ( .A(n_387), .Y(n_412) );
AND2x4_ASAP7_75t_L g417 ( .A(n_387), .B(n_418), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_1341), .B1(n_1342), .B2(n_1646), .Y(n_388) );
INVx1_ASAP7_75t_L g1646 ( .A(n_389), .Y(n_1646) );
XNOR2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_848), .Y(n_389) );
XNOR2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_701), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_568), .B2(n_700), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND3xp33_ASAP7_75t_SL g396 ( .A(n_397), .B(n_443), .C(n_495), .Y(n_396) );
OAI31xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_420), .A3(n_432), .B(n_437), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_399), .A2(n_865), .B1(n_873), .B2(n_886), .Y(n_885) );
OAI211xp5_ASAP7_75t_L g952 ( .A1(n_399), .A2(n_953), .B(n_954), .C(n_957), .Y(n_952) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g526 ( .A(n_400), .Y(n_526) );
INVx2_ASAP7_75t_L g749 ( .A(n_400), .Y(n_749) );
INVx1_ASAP7_75t_L g945 ( .A(n_400), .Y(n_945) );
INVx4_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx4f_ASAP7_75t_L g520 ( .A(n_401), .Y(n_520) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_401), .Y(n_744) );
BUFx4f_ASAP7_75t_L g883 ( .A(n_401), .Y(n_883) );
BUFx4f_ASAP7_75t_L g1077 ( .A(n_401), .Y(n_1077) );
OR2x6_ASAP7_75t_L g1080 ( .A(n_401), .B(n_1081), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1278 ( .A1(n_401), .A2(n_524), .B1(n_533), .B2(n_1279), .C(n_1280), .Y(n_1278) );
BUFx4f_ASAP7_75t_L g1359 ( .A(n_401), .Y(n_1359) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx3_ASAP7_75t_L g761 ( .A(n_402), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g1287 ( .A(n_403), .B(n_1288), .C(n_1293), .Y(n_1287) );
NAND4xp25_ASAP7_75t_L g1568 ( .A(n_403), .B(n_1569), .C(n_1572), .D(n_1575), .Y(n_1568) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g909 ( .A(n_404), .Y(n_909) );
INVx1_ASAP7_75t_L g1360 ( .A(n_404), .Y(n_1360) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_405), .B(n_1316), .Y(n_1432) );
BUFx3_ASAP7_75t_L g579 ( .A(n_406), .Y(n_579) );
AND2x6_ASAP7_75t_L g592 ( .A(n_406), .B(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_SL g606 ( .A(n_406), .B(n_576), .Y(n_606) );
INVx1_ASAP7_75t_L g621 ( .A(n_406), .Y(n_621) );
BUFx6f_ASAP7_75t_L g1066 ( .A(n_406), .Y(n_1066) );
BUFx3_ASAP7_75t_L g1177 ( .A(n_406), .Y(n_1177) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g1317 ( .A(n_407), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_414), .B2(n_415), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_409), .A2(n_470), .B1(n_474), .B2(n_475), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_410), .A2(n_895), .B1(n_907), .B2(n_908), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_410), .A2(n_907), .B1(n_992), .B2(n_993), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_410), .A2(n_907), .B1(n_1467), .B2(n_1473), .Y(n_1472) );
AOI22xp33_ASAP7_75t_L g1523 ( .A1(n_410), .A2(n_765), .B1(n_1513), .B2(n_1524), .Y(n_1523) );
AOI22xp33_ASAP7_75t_L g1559 ( .A1(n_410), .A2(n_765), .B1(n_1549), .B2(n_1560), .Y(n_1559) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI222xp33_ASAP7_75t_L g1575 ( .A1(n_411), .A2(n_831), .B1(n_1177), .B2(n_1576), .C1(n_1577), .C2(n_1578), .Y(n_1575) );
AOI22xp33_ASAP7_75t_L g1917 ( .A1(n_411), .A2(n_417), .B1(n_1909), .B2(n_1918), .Y(n_1917) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
OR2x2_ASAP7_75t_L g428 ( .A(n_412), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g763 ( .A(n_412), .B(n_413), .Y(n_763) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_412), .B(n_943), .Y(n_1289) );
INVx1_ASAP7_75t_L g610 ( .A(n_413), .Y(n_610) );
BUFx2_ASAP7_75t_L g947 ( .A(n_413), .Y(n_947) );
INVx1_ASAP7_75t_L g1087 ( .A(n_413), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_413), .A2(n_949), .B1(n_1135), .B2(n_1154), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1433 ( .A1(n_415), .A2(n_763), .B1(n_1422), .B2(n_1434), .Y(n_1433) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g766 ( .A(n_417), .Y(n_766) );
BUFx3_ASAP7_75t_L g907 ( .A(n_417), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_418), .B(n_593), .Y(n_643) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g769 ( .A(n_423), .Y(n_769) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_423), .Y(n_998) );
BUFx6f_ASAP7_75t_L g1436 ( .A(n_423), .Y(n_1436) );
AND2x4_ASAP7_75t_L g434 ( .A(n_424), .B(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g1291 ( .A(n_426), .Y(n_1291) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g1569 ( .A1(n_427), .A2(n_1289), .B1(n_1570), .B2(n_1571), .Y(n_1569) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g771 ( .A(n_428), .Y(n_771) );
BUFx2_ASAP7_75t_L g903 ( .A(n_428), .Y(n_903) );
INVx8_ASAP7_75t_L g511 ( .A(n_429), .Y(n_511) );
BUFx2_ASAP7_75t_L g617 ( .A(n_429), .Y(n_617) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx4_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g756 ( .A(n_434), .Y(n_756) );
INVx3_ASAP7_75t_SL g996 ( .A(n_434), .Y(n_996) );
INVx2_ASAP7_75t_L g583 ( .A(n_435), .Y(n_583) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_435), .Y(n_601) );
BUFx3_ASAP7_75t_L g955 ( .A(n_435), .Y(n_955) );
OAI31xp33_ASAP7_75t_L g754 ( .A1(n_437), .A2(n_755), .A3(n_757), .B(n_768), .Y(n_754) );
OAI31xp33_ASAP7_75t_L g1428 ( .A1(n_437), .A2(n_1429), .A3(n_1430), .B(n_1435), .Y(n_1428) );
BUFx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI31xp33_ASAP7_75t_L g827 ( .A1(n_438), .A2(n_828), .A3(n_833), .B(n_834), .Y(n_827) );
BUFx2_ASAP7_75t_SL g910 ( .A(n_438), .Y(n_910) );
OAI31xp33_ASAP7_75t_L g989 ( .A1(n_438), .A2(n_990), .A3(n_994), .B(n_997), .Y(n_989) );
BUFx2_ASAP7_75t_L g1299 ( .A(n_438), .Y(n_1299) );
AOI22xp5_ASAP7_75t_L g1567 ( .A1(n_438), .A2(n_786), .B1(n_1568), .B2(n_1579), .Y(n_1567) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g642 ( .A(n_440), .B(n_643), .Y(n_642) );
INVxp67_ASAP7_75t_L g651 ( .A(n_440), .Y(n_651) );
INVx1_ASAP7_75t_L g921 ( .A(n_440), .Y(n_921) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g494 ( .A(n_441), .Y(n_494) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI31xp33_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_457), .A3(n_477), .B(n_488), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g1586 ( .A1(n_446), .A2(n_479), .B1(n_1573), .B2(n_1574), .Y(n_1586) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_447), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g1553 ( .A(n_447), .Y(n_1553) );
INVx1_ASAP7_75t_L g1906 ( .A(n_447), .Y(n_1906) );
OR2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
OR2x4_ASAP7_75t_L g455 ( .A(n_448), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g545 ( .A(n_448), .Y(n_545) );
BUFx4f_ASAP7_75t_L g566 ( .A(n_448), .Y(n_566) );
BUFx3_ASAP7_75t_L g712 ( .A(n_448), .Y(n_712) );
BUFx3_ASAP7_75t_L g1116 ( .A(n_448), .Y(n_1116) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_449), .Y(n_464) );
AND2x4_ASAP7_75t_L g467 ( .A(n_449), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g483 ( .A(n_449), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_449), .B(n_463), .Y(n_487) );
INVx1_ASAP7_75t_L g648 ( .A(n_450), .Y(n_648) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_L g482 ( .A(n_451), .Y(n_482) );
INVx1_ASAP7_75t_L g456 ( .A(n_452), .Y(n_456) );
AND2x4_ASAP7_75t_L g466 ( .A(n_452), .B(n_467), .Y(n_466) );
OR2x6_ASAP7_75t_L g485 ( .A(n_452), .B(n_486), .Y(n_485) );
NAND3x1_ASAP7_75t_L g560 ( .A(n_452), .B(n_561), .C(n_563), .Y(n_560) );
AND2x4_ASAP7_75t_L g649 ( .A(n_452), .B(n_650), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g674 ( .A(n_452), .B(n_563), .Y(n_674) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g472 ( .A(n_453), .Y(n_472) );
NAND2xp33_ASAP7_75t_SL g542 ( .A(n_453), .B(n_491), .Y(n_542) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_SL g783 ( .A(n_455), .Y(n_783) );
BUFx3_ASAP7_75t_L g1306 ( .A(n_455), .Y(n_1306) );
BUFx2_ASAP7_75t_L g1509 ( .A(n_455), .Y(n_1509) );
AND2x4_ASAP7_75t_L g479 ( .A(n_456), .B(n_480), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g1461 ( .A1(n_458), .A2(n_544), .B1(n_1446), .B2(n_1452), .Y(n_1461) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g983 ( .A(n_459), .Y(n_983) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g644 ( .A(n_460), .B(n_634), .Y(n_644) );
INVx4_ASAP7_75t_L g778 ( .A(n_460), .Y(n_778) );
BUFx6f_ASAP7_75t_L g812 ( .A(n_460), .Y(n_812) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g548 ( .A(n_461), .Y(n_548) );
BUFx2_ASAP7_75t_L g733 ( .A(n_461), .Y(n_733) );
NAND2x1p5_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
BUFx2_ASAP7_75t_L g476 ( .A(n_462), .Y(n_476) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g468 ( .A(n_463), .Y(n_468) );
BUFx2_ASAP7_75t_L g473 ( .A(n_464), .Y(n_473) );
AND2x4_ASAP7_75t_L g665 ( .A(n_464), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g682 ( .A(n_464), .Y(n_682) );
CKINVDCx8_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
CKINVDCx8_ASAP7_75t_R g1037 ( .A(n_466), .Y(n_1037) );
OAI31xp33_ASAP7_75t_L g1227 ( .A1(n_466), .A2(n_1228), .A3(n_1238), .B(n_1239), .Y(n_1227) );
AOI211xp5_ASAP7_75t_L g1580 ( .A1(n_466), .A2(n_1246), .B(n_1578), .C(n_1581), .Y(n_1580) );
BUFx2_ASAP7_75t_L g660 ( .A(n_467), .Y(n_660) );
INVx2_ASAP7_75t_L g677 ( .A(n_467), .Y(n_677) );
BUFx2_ASAP7_75t_L g699 ( .A(n_467), .Y(n_699) );
BUFx3_ASAP7_75t_L g1101 ( .A(n_467), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1110 ( .A(n_467), .Y(n_1110) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_467), .Y(n_1225) );
INVx1_ASAP7_75t_L g666 ( .A(n_468), .Y(n_666) );
AOI22xp33_ASAP7_75t_SL g779 ( .A1(n_470), .A2(n_475), .B1(n_764), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_470), .A2(n_475), .B1(n_830), .B2(n_843), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_470), .A2(n_475), .B1(n_895), .B2(n_896), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g1235 ( .A1(n_470), .A2(n_475), .B1(n_1236), .B2(n_1237), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_470), .A2(n_475), .B1(n_1422), .B2(n_1423), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_470), .A2(n_475), .B1(n_1467), .B2(n_1468), .Y(n_1466) );
INVx1_ASAP7_75t_L g1582 ( .A(n_470), .Y(n_1582) );
AOI22xp33_ASAP7_75t_L g1908 ( .A1(n_470), .A2(n_475), .B1(n_1909), .B2(n_1910), .Y(n_1908) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
AND2x4_ASAP7_75t_L g475 ( .A(n_471), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_471), .B(n_473), .Y(n_1040) );
A2O1A1Ixp33_ASAP7_75t_L g1228 ( .A1(n_471), .A2(n_1229), .B(n_1232), .C(n_1235), .Y(n_1228) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND3x4_ASAP7_75t_L g655 ( .A(n_472), .B(n_491), .C(n_628), .Y(n_655) );
BUFx6f_ASAP7_75t_L g1041 ( .A(n_475), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g1352 ( .A1(n_475), .A2(n_1353), .B1(n_1354), .B2(n_1355), .Y(n_1352) );
INVx1_ASAP7_75t_L g1583 ( .A(n_475), .Y(n_1583) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g774 ( .A(n_479), .Y(n_774) );
INVx2_ASAP7_75t_L g838 ( .A(n_479), .Y(n_838) );
INVxp67_ASAP7_75t_L g1302 ( .A(n_479), .Y(n_1302) );
INVx1_ASAP7_75t_L g1516 ( .A(n_479), .Y(n_1516) );
INVx1_ASAP7_75t_L g1554 ( .A(n_479), .Y(n_1554) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_480), .Y(n_662) );
INVx1_ASAP7_75t_L g716 ( .A(n_480), .Y(n_716) );
BUFx6f_ASAP7_75t_L g1120 ( .A(n_480), .Y(n_1120) );
INVx2_ASAP7_75t_L g1902 ( .A(n_480), .Y(n_1902) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx8_ASAP7_75t_L g551 ( .A(n_481), .Y(n_551) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_481), .Y(n_670) );
INVx2_ASAP7_75t_L g804 ( .A(n_481), .Y(n_804) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
AND2x4_ASAP7_75t_L g647 ( .A(n_483), .B(n_648), .Y(n_647) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g785 ( .A(n_485), .Y(n_785) );
INVx2_ASAP7_75t_L g846 ( .A(n_485), .Y(n_846) );
INVx1_ASAP7_75t_L g1426 ( .A(n_485), .Y(n_1426) );
BUFx3_ASAP7_75t_L g552 ( .A(n_486), .Y(n_552) );
INVx1_ASAP7_75t_L g720 ( .A(n_486), .Y(n_720) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g557 ( .A(n_487), .Y(n_557) );
OAI31xp33_ASAP7_75t_SL g891 ( .A1(n_488), .A2(n_892), .A3(n_893), .B(n_897), .Y(n_891) );
OAI31xp33_ASAP7_75t_L g1032 ( .A1(n_488), .A2(n_1033), .A3(n_1036), .B(n_1043), .Y(n_1032) );
AND2x2_ASAP7_75t_SL g488 ( .A(n_489), .B(n_492), .Y(n_488) );
AND2x4_ASAP7_75t_L g786 ( .A(n_489), .B(n_492), .Y(n_786) );
AND2x2_ASAP7_75t_L g847 ( .A(n_489), .B(n_492), .Y(n_847) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_489), .B(n_492), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_489), .B(n_492), .Y(n_1427) );
INVx1_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g650 ( .A(n_491), .Y(n_650) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g532 ( .A(n_494), .Y(n_532) );
OR2x2_ASAP7_75t_L g541 ( .A(n_494), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g634 ( .A(n_494), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_SL g824 ( .A(n_494), .B(n_533), .Y(n_824) );
NOR2xp33_ASAP7_75t_SL g495 ( .A(n_496), .B(n_539), .Y(n_495) );
OAI33xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_502), .A3(n_512), .B1(n_521), .B2(n_528), .B3(n_534), .Y(n_496) );
OAI33xp33_ASAP7_75t_L g1021 ( .A1(n_497), .A2(n_528), .A3(n_1022), .B1(n_1028), .B2(n_1030), .B3(n_1031), .Y(n_1021) );
INVx1_ASAP7_75t_L g1073 ( .A(n_497), .Y(n_1073) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g737 ( .A(n_498), .Y(n_737) );
INVx4_ASAP7_75t_L g817 ( .A(n_498), .Y(n_817) );
INVx2_ASAP7_75t_L g880 ( .A(n_498), .Y(n_880) );
INVx1_ASAP7_75t_L g1497 ( .A(n_498), .Y(n_1497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
OR2x6_ASAP7_75t_L g673 ( .A(n_499), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g1129 ( .A(n_499), .Y(n_1129) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g628 ( .A(n_500), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_500), .B(n_593), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_507), .B2(n_508), .Y(n_502) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_503), .A2(n_525), .B1(n_544), .B2(n_546), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_504), .A2(n_535), .B1(n_536), .B2(n_538), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_504), .A2(n_508), .B1(n_858), .B2(n_876), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g1444 ( .A1(n_504), .A2(n_508), .B1(n_1445), .B2(n_1446), .Y(n_1444) );
OAI22xp5_ASAP7_75t_L g1453 ( .A1(n_504), .A2(n_536), .B1(n_1454), .B2(n_1455), .Y(n_1453) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g1499 ( .A(n_505), .Y(n_1499) );
INVx3_ASAP7_75t_L g1894 ( .A(n_505), .Y(n_1894) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g1025 ( .A(n_506), .Y(n_1025) );
INVx4_ASAP7_75t_L g1182 ( .A(n_506), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g564 ( .A1(n_507), .A2(n_527), .B1(n_565), .B2(n_567), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_508), .A2(n_522), .B1(n_859), .B2(n_878), .Y(n_884) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_510), .A2(n_1394), .B1(n_1395), .B2(n_1397), .Y(n_1393) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g537 ( .A(n_511), .Y(n_537) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_511), .Y(n_740) );
INVx2_ASAP7_75t_L g753 ( .A(n_511), .Y(n_753) );
INVx4_ASAP7_75t_L g819 ( .A(n_511), .Y(n_819) );
INVx2_ASAP7_75t_L g1071 ( .A(n_511), .Y(n_1071) );
INVx2_ASAP7_75t_L g1272 ( .A(n_511), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_519), .B2(n_520), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_513), .A2(n_535), .B1(n_550), .B2(n_552), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_514), .A2(n_861), .B1(n_870), .B2(n_883), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g1447 ( .A1(n_514), .A2(n_883), .B1(n_1448), .B2(n_1449), .Y(n_1447) );
OAI22xp5_ASAP7_75t_L g1544 ( .A1(n_514), .A2(n_1404), .B1(n_1531), .B2(n_1540), .Y(n_1544) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g1375 ( .A(n_515), .Y(n_1375) );
INVx2_ASAP7_75t_L g1400 ( .A(n_515), .Y(n_1400) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g524 ( .A(n_517), .Y(n_524) );
INVx1_ASAP7_75t_L g743 ( .A(n_517), .Y(n_743) );
INVx2_ASAP7_75t_L g748 ( .A(n_517), .Y(n_748) );
BUFx2_ASAP7_75t_L g821 ( .A(n_517), .Y(n_821) );
AND2x2_ASAP7_75t_L g588 ( .A(n_518), .B(n_589), .Y(n_588) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_518), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_519), .A2(n_538), .B1(n_554), .B2(n_555), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_520), .A2(n_1008), .B1(n_1013), .B2(n_1029), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_520), .A2(n_1006), .B1(n_1020), .B2(n_1029), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_525), .B1(n_526), .B2(n_527), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g1371 ( .A1(n_522), .A2(n_1359), .B1(n_1372), .B2(n_1373), .Y(n_1371) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_522), .A2(n_1404), .B1(n_1451), .B2(n_1452), .Y(n_1450) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI21xp33_ASAP7_75t_L g1178 ( .A1(n_524), .A2(n_533), .B(n_1179), .Y(n_1178) );
HB1xp67_ASAP7_75t_L g1505 ( .A(n_524), .Y(n_1505) );
OAI22xp5_ASAP7_75t_L g1543 ( .A1(n_524), .A2(n_883), .B1(n_1533), .B2(n_1536), .Y(n_1543) );
OAI211xp5_ASAP7_75t_SL g1640 ( .A1(n_526), .A2(n_1641), .B(n_1642), .C(n_1644), .Y(n_1640) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI33xp33_ASAP7_75t_L g1443 ( .A1(n_530), .A2(n_817), .A3(n_1444), .B1(n_1447), .B2(n_1450), .B3(n_1453), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x4_ASAP7_75t_L g751 ( .A(n_531), .B(n_533), .Y(n_751) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_SL g584 ( .A(n_533), .Y(n_584) );
INVx4_ASAP7_75t_L g964 ( .A(n_533), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g1506 ( .A1(n_536), .A2(n_886), .B1(n_1489), .B2(n_1492), .Y(n_1506) );
BUFx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI33xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_543), .A3(n_549), .B1(n_553), .B2(n_558), .B3(n_564), .Y(n_539) );
OAI33xp33_ASAP7_75t_L g1456 ( .A1(n_540), .A2(n_1226), .A3(n_1457), .B1(n_1458), .B2(n_1460), .B3(n_1461), .Y(n_1456) );
OAI33xp33_ASAP7_75t_L g1483 ( .A1(n_540), .A2(n_558), .A3(n_1484), .B1(n_1487), .B2(n_1490), .B3(n_1493), .Y(n_1483) );
OAI33xp33_ASAP7_75t_L g1528 ( .A1(n_540), .A2(n_558), .A3(n_1529), .B1(n_1532), .B2(n_1535), .B3(n_1538), .Y(n_1528) );
BUFx4f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx8_ASAP7_75t_L g707 ( .A(n_541), .Y(n_707) );
BUFx2_ASAP7_75t_L g793 ( .A(n_541), .Y(n_793) );
BUFx4f_ASAP7_75t_L g856 ( .A(n_541), .Y(n_856) );
BUFx2_ASAP7_75t_L g1125 ( .A(n_542), .Y(n_1125) );
OR2x2_ASAP7_75t_L g690 ( .A(n_544), .B(n_691), .Y(n_690) );
OR2x6_ASAP7_75t_L g922 ( .A(n_544), .B(n_691), .Y(n_922) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_544), .Y(n_1005) );
OAI22xp33_ASAP7_75t_L g1457 ( .A1(n_544), .A2(n_567), .B1(n_1445), .B2(n_1451), .Y(n_1457) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx3_ASAP7_75t_L g797 ( .A(n_545), .Y(n_797) );
OAI22xp33_ASAP7_75t_L g708 ( .A1(n_546), .A2(n_709), .B1(n_710), .B2(n_713), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_546), .A2(n_1004), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
OAI22xp33_ASAP7_75t_L g1538 ( .A1(n_546), .A2(n_728), .B1(n_1539), .B2(n_1540), .Y(n_1538) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_548), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g1535 ( .A1(n_550), .A2(n_877), .B1(n_1536), .B2(n_1537), .Y(n_1535) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx3_ASAP7_75t_L g554 ( .A(n_551), .Y(n_554) );
AND2x4_ASAP7_75t_L g694 ( .A(n_551), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_SL g979 ( .A(n_551), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_552), .A2(n_1448), .B1(n_1454), .B2(n_1459), .Y(n_1458) );
OAI22xp5_ASAP7_75t_L g1487 ( .A1(n_552), .A2(n_1009), .B1(n_1488), .B2(n_1489), .Y(n_1487) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_552), .A2(n_1009), .B1(n_1533), .B2(n_1534), .Y(n_1532) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_554), .A2(n_1011), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
INVx1_ASAP7_75t_L g1336 ( .A(n_554), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_555), .A2(n_802), .B1(n_803), .B2(n_805), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g1898 ( .A1(n_555), .A2(n_1887), .B1(n_1893), .B2(n_1899), .Y(n_1898) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
CKINVDCx8_ASAP7_75t_R g725 ( .A(n_556), .Y(n_725) );
INVx3_ASAP7_75t_L g877 ( .A(n_556), .Y(n_877) );
INVx3_ASAP7_75t_L g1011 ( .A(n_556), .Y(n_1011) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g633 ( .A(n_557), .Y(n_633) );
OAI33xp33_ASAP7_75t_L g854 ( .A1(n_558), .A2(n_855), .A3(n_857), .B1(n_860), .B2(n_867), .B3(n_874), .Y(n_854) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g726 ( .A(n_559), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g971 ( .A1(n_559), .A2(n_698), .B1(n_972), .B2(n_977), .C(n_984), .Y(n_971) );
INVx2_ASAP7_75t_L g1226 ( .A(n_559), .Y(n_1226) );
NAND3xp33_ASAP7_75t_L g1334 ( .A(n_559), .B(n_1335), .C(n_1338), .Y(n_1334) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g1017 ( .A(n_560), .Y(n_1017) );
OAI33xp33_ASAP7_75t_L g1410 ( .A1(n_560), .A2(n_707), .A3(n_1411), .B1(n_1413), .B2(n_1414), .B3(n_1416), .Y(n_1410) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g637 ( .A(n_562), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_562), .B(n_576), .Y(n_1060) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_565), .A2(n_567), .B1(n_858), .B2(n_859), .Y(n_857) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_566), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_566), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_980) );
OAI22xp33_ASAP7_75t_L g1484 ( .A1(n_567), .A2(n_728), .B1(n_1485), .B2(n_1486), .Y(n_1484) );
OAI22xp33_ASAP7_75t_L g1493 ( .A1(n_567), .A2(n_728), .B1(n_1494), .B2(n_1495), .Y(n_1493) );
OAI22xp33_ASAP7_75t_L g1529 ( .A1(n_567), .A2(n_728), .B1(n_1530), .B2(n_1531), .Y(n_1529) );
INVx1_ASAP7_75t_L g700 ( .A(n_568), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_629), .C(n_652), .Y(n_569) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_602), .B(n_624), .Y(n_570) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
INVx3_ASAP7_75t_L g1627 ( .A(n_573), .Y(n_1627) );
AND2x4_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx1_ASAP7_75t_L g1265 ( .A(n_574), .Y(n_1265) );
BUFx2_ASAP7_75t_L g1327 ( .A(n_574), .Y(n_1327) );
HB1xp67_ASAP7_75t_L g1636 ( .A(n_574), .Y(n_1636) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g591 ( .A(n_575), .Y(n_591) );
BUFx3_ASAP7_75t_L g959 ( .A(n_575), .Y(n_959) );
BUFx3_ASAP7_75t_L g1161 ( .A(n_575), .Y(n_1161) );
AND2x2_ASAP7_75t_L g597 ( .A(n_576), .B(n_588), .Y(n_597) );
AND2x4_ASAP7_75t_L g600 ( .A(n_576), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g930 ( .A(n_576), .B(n_601), .Y(n_930) );
AND2x2_ASAP7_75t_L g968 ( .A(n_576), .B(n_590), .Y(n_968) );
BUFx2_ASAP7_75t_L g1168 ( .A(n_576), .Y(n_1168) );
AOI21xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_585), .B(n_592), .Y(n_577) );
AOI222xp33_ASAP7_75t_L g1293 ( .A1(n_579), .A2(n_763), .B1(n_831), .B2(n_1294), .C1(n_1295), .C2(n_1296), .Y(n_1293) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g1064 ( .A(n_581), .Y(n_1064) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g1321 ( .A(n_582), .Y(n_1321) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g1643 ( .A(n_583), .Y(n_1643) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g958 ( .A(n_587), .Y(n_958) );
INVx1_ASAP7_75t_L g1313 ( .A(n_587), .Y(n_1313) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_588), .B(n_593), .Y(n_638) );
BUFx6f_ASAP7_75t_L g943 ( .A(n_588), .Y(n_943) );
AND2x4_ASAP7_75t_L g1058 ( .A(n_590), .B(n_1059), .Y(n_1058) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g1207 ( .A(n_591), .Y(n_1207) );
AOI21xp5_ASAP7_75t_L g1632 ( .A1(n_592), .A2(n_1633), .B(n_1635), .Y(n_1632) );
INVx1_ASAP7_75t_L g611 ( .A(n_593), .Y(n_611) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_593), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_598), .B2(n_599), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g1628 ( .A1(n_596), .A2(n_1629), .B1(n_1630), .B2(n_1631), .Y(n_1628) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g920 ( .A(n_597), .B(n_921), .Y(n_920) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx6f_ASAP7_75t_L g1631 ( .A(n_600), .Y(n_1631) );
BUFx6f_ASAP7_75t_L g963 ( .A(n_601), .Y(n_963) );
INVx2_ASAP7_75t_L g1171 ( .A(n_601), .Y(n_1171) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g969 ( .A(n_604), .Y(n_969) );
INVx2_ASAP7_75t_L g1638 ( .A(n_604), .Y(n_1638) );
INVx4_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g1639 ( .A(n_609), .Y(n_1639) );
NOR2x1_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g1212 ( .A(n_610), .Y(n_1212) );
INVx1_ASAP7_75t_L g1276 ( .A(n_611), .Y(n_1276) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_616), .B1(n_617), .B2(n_618), .C(n_619), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_613), .A2(n_709), .B1(n_730), .B2(n_739), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_613), .A2(n_717), .B1(n_724), .B2(n_753), .Y(n_752) );
OAI22xp33_ASAP7_75t_L g818 ( .A1(n_613), .A2(n_795), .B1(n_811), .B2(n_819), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_613), .A2(n_739), .B1(n_1408), .B2(n_1409), .Y(n_1407) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
BUFx3_ASAP7_75t_L g1069 ( .A(n_615), .Y(n_1069) );
BUFx3_ASAP7_75t_L g1369 ( .A(n_615), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_617), .A2(n_805), .B1(n_809), .B2(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g956 ( .A(n_623), .Y(n_956) );
OAI221xp5_ASAP7_75t_L g1162 ( .A1(n_623), .A2(n_749), .B1(n_1163), .B2(n_1164), .C(n_1165), .Y(n_1162) );
INVx1_ASAP7_75t_L g1205 ( .A(n_623), .Y(n_1205) );
OAI221xp5_ASAP7_75t_L g1266 ( .A1(n_623), .A2(n_749), .B1(n_1029), .B2(n_1267), .C(n_1268), .Y(n_1266) );
OAI21xp5_ASAP7_75t_SL g1625 ( .A1(n_624), .A2(n_1626), .B(n_1637), .Y(n_1625) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_626), .Y(n_970) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI31xp33_ASAP7_75t_L g1157 ( .A1(n_627), .A2(n_1158), .A3(n_1166), .B(n_1176), .Y(n_1157) );
HB1xp67_ASAP7_75t_L g1193 ( .A(n_627), .Y(n_1193) );
OAI31xp33_ASAP7_75t_L g1262 ( .A1(n_627), .A2(n_1263), .A3(n_1269), .B(n_1277), .Y(n_1262) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI21xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_639), .B(n_640), .Y(n_629) );
AOI21xp33_ASAP7_75t_L g1620 ( .A1(n_630), .A2(n_1621), .B(n_1622), .Y(n_1620) );
INVx8_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
INVx1_ASAP7_75t_L g1139 ( .A(n_632), .Y(n_1139) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
BUFx3_ASAP7_75t_L g808 ( .A(n_633), .Y(n_808) );
INVx1_ASAP7_75t_L g692 ( .A(n_634), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_634), .Y(n_695) );
INVx1_ASAP7_75t_L g1113 ( .A(n_635), .Y(n_1113) );
INVx1_ASAP7_75t_L g1056 ( .A(n_636), .Y(n_1056) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AND2x4_ASAP7_75t_L g683 ( .A(n_637), .B(n_649), .Y(n_683) );
AND2x4_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
AND2x4_ASAP7_75t_L g1623 ( .A(n_642), .B(n_644), .Y(n_1623) );
INVx2_ASAP7_75t_L g1134 ( .A(n_644), .Y(n_1134) );
INVx5_ASAP7_75t_L g1186 ( .A(n_645), .Y(n_1186) );
OR2x6_ASAP7_75t_L g645 ( .A(n_646), .B(n_651), .Y(n_645) );
OR2x2_ASAP7_75t_L g1624 ( .A(n_646), .B(n_651), .Y(n_1624) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
BUFx3_ASAP7_75t_L g659 ( .A(n_647), .Y(n_659) );
INVx8_ASAP7_75t_L g1100 ( .A(n_647), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1106 ( .A(n_647), .Y(n_1106) );
BUFx3_ASAP7_75t_L g1590 ( .A(n_647), .Y(n_1590) );
AND2x6_ASAP7_75t_L g1094 ( .A(n_649), .B(n_681), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_649), .B(n_688), .Y(n_1096) );
INVx1_ASAP7_75t_L g1103 ( .A(n_649), .Y(n_1103) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_689), .C(n_696), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_654), .B(n_678), .Y(n_653) );
AOI33xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .A3(n_661), .B1(n_667), .B2(n_672), .B3(n_675), .Y(n_654) );
BUFx3_ASAP7_75t_L g984 ( .A(n_655), .Y(n_984) );
AOI33xp33_ASAP7_75t_L g1141 ( .A1(n_655), .A2(n_672), .A3(n_1142), .B1(n_1144), .B2(n_1145), .B3(n_1148), .Y(n_1141) );
NAND3xp33_ASAP7_75t_L g1243 ( .A(n_655), .B(n_1244), .C(n_1245), .Y(n_1243) );
AOI33xp33_ASAP7_75t_L g1609 ( .A1(n_655), .A2(n_672), .A3(n_1610), .B1(n_1613), .B2(n_1615), .B3(n_1616), .Y(n_1609) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
BUFx3_ASAP7_75t_L g1333 ( .A(n_659), .Y(n_1333) );
INVx1_ASAP7_75t_L g1612 ( .A(n_659), .Y(n_1612) );
INVx1_ASAP7_75t_L g1415 ( .A(n_662), .Y(n_1415) );
INVx1_ASAP7_75t_L g1899 ( .A(n_662), .Y(n_1899) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g1337 ( .A(n_664), .Y(n_1337) );
INVx2_ASAP7_75t_R g1614 ( .A(n_664), .Y(n_1614) );
INVx5_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx3_ASAP7_75t_L g671 ( .A(n_665), .Y(n_671) );
BUFx3_ASAP7_75t_L g973 ( .A(n_665), .Y(n_973) );
BUFx12f_ASAP7_75t_L g1230 ( .A(n_665), .Y(n_1230) );
INVx1_ASAP7_75t_L g688 ( .A(n_666), .Y(n_688) );
INVx2_ASAP7_75t_L g1009 ( .A(n_668), .Y(n_1009) );
INVx8_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx3_ASAP7_75t_L g723 ( .A(n_669), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_669), .A2(n_718), .B1(n_1373), .B2(n_1380), .Y(n_1385) );
INVx5_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx3_ASAP7_75t_L g864 ( .A(n_670), .Y(n_864) );
INVx2_ASAP7_75t_SL g1147 ( .A(n_670), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_670), .A2(n_1143), .B1(n_1233), .B2(n_1234), .Y(n_1232) );
INVx2_ASAP7_75t_SL g1459 ( .A(n_670), .Y(n_1459) );
NAND3xp33_ASAP7_75t_L g1253 ( .A(n_672), .B(n_1254), .C(n_1255), .Y(n_1253) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI33xp33_ASAP7_75t_L g792 ( .A1(n_673), .A2(n_793), .A3(n_794), .B1(n_801), .B2(n_806), .B3(n_810), .Y(n_792) );
OAI33xp33_ASAP7_75t_L g1896 ( .A1(n_673), .A2(n_707), .A3(n_1897), .B1(n_1898), .B2(n_1900), .B3(n_1901), .Y(n_1896) );
INVx3_ASAP7_75t_L g1117 ( .A(n_674), .Y(n_1117) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g1220 ( .A(n_677), .Y(n_1220) );
INVx1_ASAP7_75t_L g1246 ( .A(n_677), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_684), .B2(n_685), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_680), .A2(n_685), .B1(n_1618), .B2(n_1619), .Y(n_1617) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
NAND2x1_ASAP7_75t_L g934 ( .A(n_681), .B(n_683), .Y(n_934) );
AND2x4_ASAP7_75t_SL g1153 ( .A(n_681), .B(n_683), .Y(n_1153) );
INVx3_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_L g685 ( .A(n_683), .B(n_686), .Y(n_685) );
AND2x4_ASAP7_75t_L g698 ( .A(n_683), .B(n_699), .Y(n_698) );
AND2x4_ASAP7_75t_SL g1155 ( .A(n_683), .B(n_686), .Y(n_1155) );
AOI221xp5_ASAP7_75t_L g932 ( .A1(n_685), .A2(n_933), .B1(n_935), .B2(n_936), .C(n_937), .Y(n_932) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g926 ( .A(n_692), .B(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_694), .B(n_1150), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_694), .B(n_1248), .Y(n_1247) );
AND2x4_ASAP7_75t_L g1136 ( .A(n_695), .B(n_1137), .Y(n_1136) );
NOR3xp33_ASAP7_75t_L g1606 ( .A(n_696), .B(n_1607), .C(n_1608), .Y(n_1606) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_698), .A2(n_1153), .B1(n_1154), .B2(n_1155), .C(n_1156), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1257 ( .A1(n_698), .A2(n_1153), .B1(n_1155), .B2(n_1258), .C(n_1259), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_787), .B2(n_788), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_754), .C(n_772), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_735), .Y(n_705) );
OAI33xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .A3(n_714), .B1(n_721), .B2(n_726), .B3(n_727), .Y(n_706) );
OAI33xp33_ASAP7_75t_L g1381 ( .A1(n_707), .A2(n_1382), .A3(n_1384), .B1(n_1385), .B2(n_1386), .B3(n_1388), .Y(n_1381) );
OAI22xp33_ASAP7_75t_L g1411 ( .A1(n_710), .A2(n_1394), .B1(n_1403), .B2(n_1412), .Y(n_1411) );
OAI22xp33_ASAP7_75t_L g1416 ( .A1(n_710), .A2(n_1397), .B1(n_1406), .B2(n_1417), .Y(n_1416) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g729 ( .A(n_712), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_713), .A2(n_734), .B1(n_746), .B2(n_749), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_714) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_715), .A2(n_722), .B1(n_742), .B2(n_744), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_718), .A2(n_1119), .B1(n_1372), .B2(n_1379), .Y(n_1384) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_718), .A2(n_1401), .B1(n_1409), .B2(n_1415), .Y(n_1414) );
INVx3_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g866 ( .A(n_720), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_725), .A2(n_1119), .B1(n_1121), .B2(n_1122), .Y(n_1118) );
OAI221xp5_ASAP7_75t_L g1215 ( .A1(n_725), .A2(n_1216), .B1(n_1217), .B2(n_1218), .C(n_1219), .Y(n_1215) );
OAI221xp5_ASAP7_75t_L g1221 ( .A1(n_725), .A2(n_1203), .B1(n_1222), .B2(n_1223), .C(n_1224), .Y(n_1221) );
OAI22xp5_ASAP7_75t_L g1413 ( .A1(n_725), .A2(n_1222), .B1(n_1399), .B2(n_1408), .Y(n_1413) );
OAI22xp5_ASAP7_75t_L g1901 ( .A1(n_725), .A2(n_1888), .B1(n_1895), .B2(n_1902), .Y(n_1901) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_730), .B1(n_731), .B2(n_734), .Y(n_727) );
OAI22xp33_ASAP7_75t_L g1382 ( .A1(n_728), .A2(n_1368), .B1(n_1376), .B2(n_1383), .Y(n_1382) );
OAI22xp33_ASAP7_75t_L g1388 ( .A1(n_728), .A2(n_976), .B1(n_1370), .B2(n_1377), .Y(n_1388) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
HB1xp67_ASAP7_75t_L g1465 ( .A(n_731), .Y(n_1465) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g1412 ( .A(n_732), .Y(n_1412) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g800 ( .A(n_733), .Y(n_800) );
OAI33xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .A3(n_741), .B1(n_745), .B2(n_750), .B3(n_752), .Y(n_735) );
OAI33xp33_ASAP7_75t_L g1392 ( .A1(n_736), .A2(n_750), .A3(n_1393), .B1(n_1398), .B2(n_1402), .B3(n_1407), .Y(n_1392) );
INVx1_ASAP7_75t_L g1596 ( .A(n_736), .Y(n_1596) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g1378 ( .A1(n_739), .A2(n_826), .B1(n_1379), .B2(n_1380), .Y(n_1378) );
OAI22xp33_ASAP7_75t_L g1545 ( .A1(n_739), .A2(n_886), .B1(n_1534), .B2(n_1537), .Y(n_1545) );
INVx5_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx6_ASAP7_75t_L g1500 ( .A(n_740), .Y(n_1500) );
OAI221xp5_ASAP7_75t_L g1075 ( .A1(n_742), .A2(n_1076), .B1(n_1077), .B2(n_1078), .C(n_1079), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_742), .A2(n_1403), .B1(n_1404), .B2(n_1406), .Y(n_1402) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx4_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g1029 ( .A(n_748), .Y(n_1029) );
INVx2_ASAP7_75t_L g1165 ( .A(n_748), .Y(n_1165) );
OAI211xp5_ASAP7_75t_L g960 ( .A1(n_749), .A2(n_961), .B(n_962), .C(n_965), .Y(n_960) );
OAI21xp5_ASAP7_75t_L g1074 ( .A1(n_750), .A2(n_1075), .B(n_1080), .Y(n_1074) );
OAI33xp33_ASAP7_75t_L g1366 ( .A1(n_750), .A2(n_815), .A3(n_1367), .B1(n_1371), .B2(n_1374), .B3(n_1378), .Y(n_1366) );
OAI33xp33_ASAP7_75t_L g1882 ( .A1(n_750), .A2(n_815), .A3(n_1883), .B1(n_1886), .B2(n_1889), .B3(n_1892), .Y(n_1882) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g890 ( .A(n_751), .Y(n_890) );
NAND3xp33_ASAP7_75t_L g1319 ( .A(n_751), .B(n_1320), .C(n_1326), .Y(n_1319) );
AOI33xp33_ASAP7_75t_L g1595 ( .A1(n_751), .A2(n_1596), .A3(n_1597), .B1(n_1600), .B2(n_1602), .B3(n_1603), .Y(n_1595) );
OAI22xp33_ASAP7_75t_L g1367 ( .A1(n_753), .A2(n_1368), .B1(n_1369), .B2(n_1370), .Y(n_1367) );
OAI22xp5_ASAP7_75t_L g1892 ( .A1(n_753), .A2(n_1893), .B1(n_1894), .B2(n_1895), .Y(n_1892) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_760), .A2(n_802), .B1(n_807), .B2(n_821), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_760), .A2(n_798), .B1(n_813), .B2(n_821), .Y(n_822) );
BUFx2_ASAP7_75t_L g905 ( .A(n_760), .Y(n_905) );
BUFx3_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_761), .B(n_1060), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_761), .B(n_1175), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_761), .B(n_1275), .Y(n_1274) );
INVx2_ASAP7_75t_SL g1405 ( .A(n_761), .Y(n_1405) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_765), .B2(n_767), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_763), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_763), .A2(n_765), .B1(n_1354), .B2(n_1362), .Y(n_1361) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g831 ( .A(n_766), .Y(n_831) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g999 ( .A(n_771), .Y(n_999) );
INVx2_ASAP7_75t_L g1437 ( .A(n_771), .Y(n_1437) );
OAI31xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_775), .A3(n_781), .B(n_786), .Y(n_772) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OAI22xp33_ASAP7_75t_L g1897 ( .A1(n_777), .A2(n_797), .B1(n_1884), .B2(n_1890), .Y(n_1897) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g841 ( .A(n_778), .Y(n_841) );
INVx2_ASAP7_75t_L g976 ( .A(n_778), .Y(n_976) );
INVx1_ASAP7_75t_L g1383 ( .A(n_778), .Y(n_1383) );
INVx1_ASAP7_75t_L g1417 ( .A(n_778), .Y(n_1417) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g1044 ( .A(n_783), .Y(n_1044) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OAI31xp33_ASAP7_75t_L g1300 ( .A1(n_786), .A2(n_1301), .A3(n_1303), .B(n_1305), .Y(n_1300) );
OAI31xp33_ASAP7_75t_L g1348 ( .A1(n_786), .A2(n_1349), .A3(n_1350), .B(n_1356), .Y(n_1348) );
OAI31xp33_ASAP7_75t_L g1462 ( .A1(n_786), .A2(n_1463), .A3(n_1464), .B(n_1469), .Y(n_1462) );
OAI31xp33_ASAP7_75t_L g1546 ( .A1(n_786), .A2(n_1547), .A3(n_1551), .B(n_1552), .Y(n_1546) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_827), .C(n_836), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_814), .Y(n_791) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_796), .B1(n_798), .B2(n_799), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_796), .A2(n_961), .B1(n_975), .B2(n_976), .Y(n_974) );
BUFx4f_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
OAI22xp33_ASAP7_75t_L g810 ( .A1(n_797), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
OAI22xp33_ASAP7_75t_L g1900 ( .A1(n_797), .A2(n_799), .B1(n_1885), .B2(n_1891), .Y(n_1900) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVxp67_ASAP7_75t_L g1511 ( .A(n_800), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_803), .A2(n_807), .B1(n_808), .B2(n_809), .Y(n_806) );
INVx2_ASAP7_75t_L g1330 ( .A(n_803), .Y(n_1330) );
BUFx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g869 ( .A(n_804), .Y(n_869) );
INVx3_ASAP7_75t_L g927 ( .A(n_804), .Y(n_927) );
INVx1_ASAP7_75t_L g872 ( .A(n_812), .Y(n_872) );
OAI33xp33_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_818), .A3(n_820), .B1(n_822), .B2(n_823), .B3(n_825), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_SL g1318 ( .A(n_817), .Y(n_1318) );
INVx2_ASAP7_75t_L g1027 ( .A(n_819), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1180 ( .A1(n_819), .A2(n_1181), .B1(n_1182), .B2(n_1183), .Y(n_1180) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OAI22xp33_ASAP7_75t_L g1883 ( .A1(n_826), .A2(n_1070), .B1(n_1884), .B2(n_1885), .Y(n_1883) );
INVx1_ASAP7_75t_L g1915 ( .A(n_835), .Y(n_1915) );
OAI31xp33_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_839), .A3(n_844), .B(n_847), .Y(n_836) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g1115 ( .A1(n_841), .A2(n_1072), .B1(n_1078), .B2(n_1116), .C(n_1117), .Y(n_1115) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g1584 ( .A1(n_846), .A2(n_1570), .B1(n_1571), .B2(n_1585), .Y(n_1584) );
OAI31xp33_ASAP7_75t_L g1903 ( .A1(n_847), .A2(n_1904), .A3(n_1907), .B(n_1911), .Y(n_1903) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
XNOR2x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_1047), .Y(n_849) );
XNOR2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_911), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_891), .C(n_898), .Y(n_852) );
NOR2xp33_ASAP7_75t_SL g853 ( .A(n_854), .B(n_879), .Y(n_853) );
OAI33xp33_ASAP7_75t_L g1001 ( .A1(n_855), .A2(n_1002), .A3(n_1007), .B1(n_1012), .B2(n_1015), .B3(n_1018), .Y(n_1001) );
OAI22xp33_ASAP7_75t_L g1214 ( .A1(n_855), .A2(n_1215), .B1(n_1221), .B2(n_1226), .Y(n_1214) );
BUFx3_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OAI22xp33_ASAP7_75t_SL g860 ( .A1(n_861), .A2(n_862), .B1(n_865), .B2(n_866), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g1490 ( .A1(n_862), .A2(n_877), .B1(n_1491), .B2(n_1492), .Y(n_1490) );
INVx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_863), .A2(n_1089), .B1(n_1090), .B2(n_1106), .Y(n_1105) );
INVx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_866), .A2(n_1009), .B1(n_1449), .B2(n_1455), .Y(n_1460) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_870), .B1(n_871), .B2(n_873), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_871), .A2(n_1003), .B1(n_1004), .B2(n_1006), .Y(n_1002) );
INVx2_ASAP7_75t_SL g871 ( .A(n_872), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_876), .B1(n_877), .B2(n_878), .Y(n_874) );
OAI33xp33_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .A3(n_882), .B1(n_884), .B2(n_885), .B3(n_890), .Y(n_879) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
OAI33xp33_ASAP7_75t_L g1496 ( .A1(n_890), .A2(n_1497), .A3(n_1498), .B1(n_1501), .B2(n_1504), .B3(n_1506), .Y(n_1496) );
OAI33xp33_ASAP7_75t_L g1541 ( .A1(n_890), .A2(n_1497), .A3(n_1542), .B1(n_1543), .B2(n_1544), .B3(n_1545), .Y(n_1541) );
OAI31xp33_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_900), .A3(n_904), .B(n_910), .Y(n_898) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx2_ASAP7_75t_SL g902 ( .A(n_903), .Y(n_902) );
HB1xp67_ASAP7_75t_L g1475 ( .A(n_903), .Y(n_1475) );
OAI31xp33_ASAP7_75t_L g1357 ( .A1(n_910), .A2(n_1358), .A3(n_1363), .B(n_1364), .Y(n_1357) );
OAI31xp33_ASAP7_75t_L g1470 ( .A1(n_910), .A2(n_1471), .A3(n_1474), .B(n_1476), .Y(n_1470) );
OAI31xp33_ASAP7_75t_SL g1517 ( .A1(n_910), .A2(n_1518), .A3(n_1519), .B(n_1520), .Y(n_1517) );
OAI31xp33_ASAP7_75t_L g1555 ( .A1(n_910), .A2(n_1556), .A3(n_1557), .B(n_1558), .Y(n_1555) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
AO22x2_ASAP7_75t_L g912 ( .A1(n_913), .A2(n_985), .B1(n_986), .B2(n_1046), .Y(n_912) );
INVx1_ASAP7_75t_SL g1046 ( .A(n_913), .Y(n_1046) );
XNOR2x1_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
NOR2x1_ASAP7_75t_L g915 ( .A(n_916), .B(n_931), .Y(n_915) );
INVxp67_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_922), .Y(n_918) );
INVx3_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
AOI22xp5_ASAP7_75t_L g1088 ( .A1(n_920), .A2(n_929), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
AND2x4_ASAP7_75t_L g929 ( .A(n_921), .B(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
NAND2x1_ASAP7_75t_L g924 ( .A(n_925), .B(n_928), .Y(n_924) );
INVx2_ASAP7_75t_SL g925 ( .A(n_926), .Y(n_925) );
INVx2_ASAP7_75t_L g1222 ( .A(n_927), .Y(n_1222) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
NAND3xp33_ASAP7_75t_SL g931 ( .A(n_932), .B(n_938), .C(n_971), .Y(n_931) );
INVx2_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_935), .A2(n_947), .B1(n_948), .B2(n_949), .Y(n_946) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_966), .B(n_970), .Y(n_938) );
NAND3xp33_ASAP7_75t_L g939 ( .A(n_940), .B(n_952), .C(n_960), .Y(n_939) );
A2O1A1Ixp33_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_942), .B(n_944), .C(n_951), .Y(n_940) );
A2O1A1Ixp33_ASAP7_75t_SL g1208 ( .A1(n_942), .A2(n_951), .B(n_1209), .C(n_1210), .Y(n_1208) );
BUFx6f_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx3_ASAP7_75t_L g1160 ( .A(n_943), .Y(n_1160) );
A2O1A1Ixp33_ASAP7_75t_L g1173 ( .A1(n_943), .A2(n_951), .B(n_1140), .C(n_1174), .Y(n_1173) );
A2O1A1Ixp33_ASAP7_75t_L g1273 ( .A1(n_943), .A2(n_1252), .B(n_1274), .C(n_1276), .Y(n_1273) );
NAND2xp5_ASAP7_75t_SL g944 ( .A(n_945), .B(n_946), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g1275 ( .A1(n_947), .A2(n_949), .B1(n_1250), .B2(n_1258), .Y(n_1275) );
INVx1_ASAP7_75t_L g1213 ( .A(n_949), .Y(n_1213) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
BUFx2_ASAP7_75t_L g1310 ( .A(n_955), .Y(n_1310) );
HB1xp67_ASAP7_75t_L g1634 ( .A(n_955), .Y(n_1634) );
BUFx3_ASAP7_75t_L g1311 ( .A(n_959), .Y(n_1311) );
INVx1_ASAP7_75t_SL g1599 ( .A(n_959), .Y(n_1599) );
BUFx3_ASAP7_75t_L g1601 ( .A(n_963), .Y(n_1601) );
INVx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_973), .A2(n_1108), .B1(n_1109), .B2(n_1110), .Y(n_1107) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
OAI211xp5_ASAP7_75t_L g1123 ( .A1(n_983), .A2(n_1076), .B(n_1124), .C(n_1126), .Y(n_1123) );
HB1xp67_ASAP7_75t_L g1351 ( .A(n_983), .Y(n_1351) );
NAND3xp33_ASAP7_75t_L g1328 ( .A(n_984), .B(n_1329), .C(n_1332), .Y(n_1328) );
AOI33xp33_ASAP7_75t_L g1587 ( .A1(n_984), .A2(n_1588), .A3(n_1591), .B1(n_1592), .B2(n_1593), .B3(n_1594), .Y(n_1587) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
NAND3xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_1000), .C(n_1032), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_992), .A2(n_1039), .B1(n_1041), .B2(n_1042), .Y(n_1038) );
NOR2xp33_ASAP7_75t_SL g1000 ( .A(n_1001), .B(n_1021), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_1003), .A2(n_1019), .B1(n_1023), .B2(n_1026), .Y(n_1022) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1009), .B1(n_1010), .B2(n_1011), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_1010), .A2(n_1014), .B1(n_1023), .B2(n_1026), .Y(n_1031) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
BUFx2_ASAP7_75t_L g1387 ( .A(n_1017), .Y(n_1387) );
BUFx2_ASAP7_75t_L g1593 ( .A(n_1017), .Y(n_1593) );
INVx2_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_1025), .Y(n_1024) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1029), .Y(n_1503) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_1035), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_1039), .A2(n_1041), .B1(n_1295), .B2(n_1296), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_1039), .A2(n_1041), .B1(n_1513), .B2(n_1514), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1548 ( .A1(n_1039), .A2(n_1041), .B1(n_1549), .B2(n_1550), .Y(n_1548) );
BUFx3_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
BUFx3_ASAP7_75t_L g1353 ( .A(n_1040), .Y(n_1353) );
XNOR2x1_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1283), .Y(n_1047) );
OA22x2_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1050), .B1(n_1188), .B2(n_1282), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
XOR2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1130), .Y(n_1050) );
XNOR2x1_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1053), .Y(n_1051) );
NAND4xp75_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1062), .C(n_1088), .D(n_1091), .Y(n_1053) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
AOI211x1_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1073), .B(n_1074), .C(n_1084), .Y(n_1062) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
AOI221xp5_ASAP7_75t_L g1169 ( .A1(n_1066), .A2(n_1150), .B1(n_1156), .B2(n_1170), .C(n_1172), .Y(n_1169) );
AOI221xp5_ASAP7_75t_L g1270 ( .A1(n_1066), .A2(n_1170), .B1(n_1248), .B2(n_1259), .C(n_1271), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1069), .B1(n_1070), .B2(n_1072), .Y(n_1067) );
BUFx6f_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
OAI211xp5_ASAP7_75t_SL g1198 ( .A1(n_1077), .A2(n_1199), .B(n_1200), .C(n_1201), .Y(n_1198) );
OAI211xp5_ASAP7_75t_SL g1202 ( .A1(n_1077), .A2(n_1203), .B(n_1204), .C(n_1206), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_1077), .A2(n_1375), .B1(n_1376), .B2(n_1377), .Y(n_1374) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
NAND2x2_ASAP7_75t_L g1085 ( .A(n_1082), .B(n_1086), .Y(n_1085) );
INVx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx2_ASAP7_75t_SL g1086 ( .A(n_1087), .Y(n_1086) );
OAI31xp67_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1104), .A3(n_1114), .B(n_1128), .Y(n_1091) );
INVx4_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
A2O1A1Ixp33_ASAP7_75t_L g1097 ( .A1(n_1098), .A2(n_1099), .B(n_1101), .C(n_1102), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g1099 ( .A(n_1100), .Y(n_1099) );
INVx3_ASAP7_75t_L g1127 ( .A(n_1100), .Y(n_1127) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1100), .Y(n_1137) );
INVx8_ASAP7_75t_L g1143 ( .A(n_1100), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_1101), .A2(n_1209), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
AOI21xp33_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1107), .B(n_1111), .Y(n_1104) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
OAI21xp5_ASAP7_75t_SL g1114 ( .A1(n_1115), .A2(n_1118), .B(n_1123), .Y(n_1114) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx2_ASAP7_75t_SL g1216 ( .A(n_1120), .Y(n_1216) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
XNOR2x1_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1187), .Y(n_1130) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1151), .Y(n_1131) );
NAND3xp33_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1141), .C(n_1149), .Y(n_1132) );
AOI222xp33_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1135), .B1(n_1136), .B2(n_1138), .C1(n_1139), .C2(n_1140), .Y(n_1133) );
AOI222xp33_ASAP7_75t_L g1249 ( .A1(n_1134), .A2(n_1136), .B1(n_1139), .B2(n_1250), .C1(n_1251), .C2(n_1252), .Y(n_1249) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
NAND3xp33_ASAP7_75t_SL g1151 ( .A(n_1152), .B(n_1157), .C(n_1184), .Y(n_1151) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
OAI21xp33_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1169), .B(n_1173), .Y(n_1166) );
OAI21xp5_ASAP7_75t_SL g1269 ( .A1(n_1167), .A2(n_1270), .B(n_1273), .Y(n_1269) );
INVxp67_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
OAI21xp5_ASAP7_75t_L g1195 ( .A1(n_1168), .A2(n_1196), .B(n_1197), .Y(n_1195) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1186), .B(n_1261), .Y(n_1260) );
XNOR2xp5_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1240), .Y(n_1188) );
XOR2xp5_ASAP7_75t_L g1282 ( .A(n_1189), .B(n_1240), .Y(n_1282) );
XNOR2x1_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1191), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1227), .Y(n_1191) );
AOI21xp5_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1194), .B(n_1214), .Y(n_1192) );
NAND4xp25_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1198), .C(n_1202), .D(n_1208), .Y(n_1194) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
HB1xp67_ASAP7_75t_L g1331 ( .A(n_1225), .Y(n_1331) );
XNOR2x1_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1281), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1256), .Y(n_1241) );
NAND4xp25_ASAP7_75t_SL g1242 ( .A(n_1243), .B(n_1247), .C(n_1249), .D(n_1253), .Y(n_1242) );
NAND3xp33_ASAP7_75t_SL g1256 ( .A(n_1257), .B(n_1260), .C(n_1262), .Y(n_1256) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1285), .Y(n_1339) );
NAND3xp33_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1300), .C(n_1307), .Y(n_1285) );
OAI21xp5_ASAP7_75t_L g1286 ( .A1(n_1287), .A2(n_1297), .B(n_1299), .Y(n_1286) );
AOI22xp5_ASAP7_75t_L g1288 ( .A1(n_1289), .A2(n_1290), .B1(n_1291), .B2(n_1292), .Y(n_1288) );
OAI31xp33_ASAP7_75t_SL g1912 ( .A1(n_1299), .A2(n_1913), .A3(n_1916), .B(n_1919), .Y(n_1912) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1306), .Y(n_1585) );
AND4x1_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1319), .C(n_1328), .D(n_1334), .Y(n_1307) );
NAND3xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1312), .C(n_1318), .Y(n_1308) );
INVx2_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1316), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
BUFx2_ASAP7_75t_L g1325 ( .A(n_1317), .Y(n_1325) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
XNOR2xp5_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1477), .Y(n_1342) );
OAI22xp5_ASAP7_75t_L g1343 ( .A1(n_1344), .A2(n_1345), .B1(n_1438), .B2(n_1439), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
XNOR2x1_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1389), .Y(n_1345) );
NAND3xp33_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1357), .C(n_1365), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g1398 ( .A1(n_1359), .A2(n_1399), .B1(n_1400), .B2(n_1401), .Y(n_1398) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1359), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1889 ( .A1(n_1359), .A2(n_1400), .B1(n_1890), .B2(n_1891), .Y(n_1889) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1381), .Y(n_1365) );
OAI22xp5_ASAP7_75t_L g1886 ( .A1(n_1375), .A2(n_1404), .B1(n_1887), .B2(n_1888), .Y(n_1886) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
NAND3xp33_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1418), .C(n_1428), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1410), .Y(n_1391) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_1404), .A2(n_1488), .B1(n_1491), .B2(n_1502), .Y(n_1501) );
OAI22xp33_ASAP7_75t_L g1504 ( .A1(n_1404), .A2(n_1486), .B1(n_1495), .B2(n_1505), .Y(n_1504) );
INVx5_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
OAI31xp33_ASAP7_75t_L g1418 ( .A1(n_1419), .A2(n_1420), .A3(n_1424), .B(n_1427), .Y(n_1418) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
OAI31xp33_ASAP7_75t_L g1507 ( .A1(n_1427), .A2(n_1508), .A3(n_1510), .B(n_1515), .Y(n_1507) );
INVx2_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
BUFx2_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
NAND3xp33_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1462), .C(n_1470), .Y(n_1441) );
NOR2xp33_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1456), .Y(n_1442) );
AOI22xp5_ASAP7_75t_L g1477 ( .A1(n_1478), .A2(n_1561), .B1(n_1562), .B2(n_1645), .Y(n_1477) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1478), .Y(n_1645) );
HB1xp67_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
XOR2xp5_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1525), .Y(n_1479) );
AND3x1_ASAP7_75t_L g1481 ( .A(n_1482), .B(n_1507), .C(n_1517), .Y(n_1481) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1496), .Y(n_1482) );
OAI22xp33_ASAP7_75t_L g1498 ( .A1(n_1485), .A2(n_1494), .B1(n_1499), .B2(n_1500), .Y(n_1498) );
OAI22xp33_ASAP7_75t_L g1542 ( .A1(n_1499), .A2(n_1500), .B1(n_1530), .B2(n_1539), .Y(n_1542) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
AND3x1_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1546), .C(n_1555), .Y(n_1526) );
NOR2xp33_ASAP7_75t_L g1527 ( .A(n_1528), .B(n_1541), .Y(n_1527) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
XNOR2x1_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1604), .Y(n_1564) );
NAND3x1_ASAP7_75t_L g1566 ( .A(n_1567), .B(n_1587), .C(n_1595), .Y(n_1566) );
NAND3xp33_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1584), .C(n_1586), .Y(n_1579) );
BUFx2_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_SL g1598 ( .A(n_1599), .Y(n_1598) );
AND3x1_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1620), .C(n_1625), .Y(n_1605) );
NAND2xp5_ASAP7_75t_SL g1608 ( .A(n_1609), .B(n_1617), .Y(n_1608) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
OAI221xp5_ASAP7_75t_L g1647 ( .A1(n_1648), .A2(n_1877), .B1(n_1879), .B2(n_1920), .C(n_1923), .Y(n_1647) );
AOI21xp5_ASAP7_75t_L g1648 ( .A1(n_1649), .A2(n_1791), .B(n_1844), .Y(n_1648) );
NAND4xp25_ASAP7_75t_L g1649 ( .A(n_1650), .B(n_1761), .C(n_1777), .D(n_1783), .Y(n_1649) );
NOR5xp2_ASAP7_75t_L g1650 ( .A(n_1651), .B(n_1715), .C(n_1728), .D(n_1735), .E(n_1758), .Y(n_1650) );
OAI21xp5_ASAP7_75t_SL g1651 ( .A1(n_1652), .A2(n_1672), .B(n_1691), .Y(n_1651) );
NOR2xp33_ASAP7_75t_L g1692 ( .A(n_1652), .B(n_1673), .Y(n_1692) );
OAI31xp33_ASAP7_75t_L g1869 ( .A1(n_1652), .A2(n_1870), .A3(n_1871), .B(n_1872), .Y(n_1869) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1790 ( .A(n_1653), .B(n_1748), .Y(n_1790) );
AOI221xp5_ASAP7_75t_L g1807 ( .A1(n_1653), .A2(n_1731), .B1(n_1808), .B2(n_1809), .C(n_1811), .Y(n_1807) );
AND2x2_ASAP7_75t_L g1653 ( .A(n_1654), .B(n_1668), .Y(n_1653) );
INVx1_ASAP7_75t_L g1718 ( .A(n_1654), .Y(n_1718) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1654), .Y(n_1730) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1654), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1654), .B(n_1706), .Y(n_1780) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1662), .Y(n_1654) );
AND2x6_ASAP7_75t_L g1656 ( .A(n_1657), .B(n_1658), .Y(n_1656) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1657), .B(n_1661), .Y(n_1660) );
AND2x4_ASAP7_75t_L g1663 ( .A(n_1657), .B(n_1664), .Y(n_1663) );
AND2x6_ASAP7_75t_L g1666 ( .A(n_1657), .B(n_1667), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1670 ( .A(n_1657), .B(n_1661), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1752 ( .A(n_1657), .B(n_1661), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1664 ( .A(n_1659), .B(n_1665), .Y(n_1664) );
OAI21xp5_ASAP7_75t_L g1932 ( .A1(n_1661), .A2(n_1933), .B(n_1934), .Y(n_1932) );
CKINVDCx5p33_ASAP7_75t_R g1706 ( .A(n_1668), .Y(n_1706) );
OR2x2_ASAP7_75t_L g1727 ( .A(n_1668), .B(n_1703), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1755 ( .A(n_1668), .B(n_1718), .Y(n_1755) );
HB1xp67_ASAP7_75t_SL g1773 ( .A(n_1668), .Y(n_1773) );
NAND2xp5_ASAP7_75t_L g1837 ( .A(n_1668), .B(n_1748), .Y(n_1837) );
NAND2xp5_ASAP7_75t_L g1849 ( .A(n_1668), .B(n_1675), .Y(n_1849) );
AND2x4_ASAP7_75t_L g1668 ( .A(n_1669), .B(n_1671), .Y(n_1668) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1672), .Y(n_1860) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1673), .B(n_1678), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1784 ( .A(n_1673), .B(n_1710), .Y(n_1784) );
NAND2xp5_ASAP7_75t_L g1867 ( .A(n_1673), .B(n_1756), .Y(n_1867) );
CKINVDCx14_ASAP7_75t_R g1673 ( .A(n_1674), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1674), .B(n_1726), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1674), .B(n_1703), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1741 ( .A(n_1674), .B(n_1695), .Y(n_1741) );
NAND2xp5_ASAP7_75t_L g1787 ( .A(n_1674), .B(n_1723), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1801 ( .A(n_1674), .B(n_1802), .Y(n_1801) );
NOR2xp33_ASAP7_75t_L g1813 ( .A(n_1674), .B(n_1727), .Y(n_1813) );
NOR2xp33_ASAP7_75t_L g1833 ( .A(n_1674), .B(n_1769), .Y(n_1833) );
NOR2xp33_ASAP7_75t_L g1843 ( .A(n_1674), .B(n_1736), .Y(n_1843) );
INVx3_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
CKINVDCx5p33_ASAP7_75t_R g1707 ( .A(n_1675), .Y(n_1707) );
NOR2xp33_ASAP7_75t_L g1744 ( .A(n_1675), .B(n_1712), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1675), .B(n_1680), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1782 ( .A(n_1675), .B(n_1696), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1817 ( .A(n_1675), .B(n_1789), .Y(n_1817) );
NAND2xp5_ASAP7_75t_L g1839 ( .A(n_1675), .B(n_1798), .Y(n_1839) );
NAND2xp5_ASAP7_75t_L g1841 ( .A(n_1675), .B(n_1723), .Y(n_1841) );
NAND2xp5_ASAP7_75t_L g1871 ( .A(n_1675), .B(n_1769), .Y(n_1871) );
AND2x4_ASAP7_75t_SL g1675 ( .A(n_1676), .B(n_1677), .Y(n_1675) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
OR2x2_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1683), .Y(n_1679) );
INVx2_ASAP7_75t_L g1695 ( .A(n_1680), .Y(n_1695) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1680), .B(n_1688), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_1680), .B(n_1697), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1772 ( .A(n_1680), .B(n_1696), .Y(n_1772) );
AND2x2_ASAP7_75t_L g1795 ( .A(n_1680), .B(n_1796), .Y(n_1795) );
NAND2xp5_ASAP7_75t_L g1810 ( .A(n_1680), .B(n_1685), .Y(n_1810) );
OAI322xp33_ASAP7_75t_L g1811 ( .A1(n_1680), .A2(n_1694), .A3(n_1789), .B1(n_1812), .B2(n_1814), .C1(n_1818), .C2(n_1820), .Y(n_1811) );
OR2x2_ASAP7_75t_L g1847 ( .A(n_1680), .B(n_1782), .Y(n_1847) );
OR2x2_ASAP7_75t_L g1858 ( .A(n_1680), .B(n_1685), .Y(n_1858) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1682), .Y(n_1680) );
OR2x2_ASAP7_75t_L g1757 ( .A(n_1683), .B(n_1695), .Y(n_1757) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1683), .Y(n_1798) );
OR2x2_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1688), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_1684), .B(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
OR2x2_ASAP7_75t_L g1712 ( .A(n_1685), .B(n_1713), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1685), .B(n_1688), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1775 ( .A(n_1685), .B(n_1695), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1686), .B(n_1687), .Y(n_1685) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1688), .Y(n_1697) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1688), .Y(n_1713) );
NAND2xp5_ASAP7_75t_L g1830 ( .A(n_1688), .B(n_1695), .Y(n_1830) );
NAND2x1_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1690), .Y(n_1688) );
AOI22xp33_ASAP7_75t_L g1691 ( .A1(n_1692), .A2(n_1693), .B1(n_1699), .B2(n_1708), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1693 ( .A(n_1694), .B(n_1698), .Y(n_1693) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_1695), .B(n_1696), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1710 ( .A(n_1695), .B(n_1711), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1695), .B(n_1723), .Y(n_1722) );
OR2x2_ASAP7_75t_L g1767 ( .A(n_1695), .B(n_1768), .Y(n_1767) );
OR2x2_ASAP7_75t_L g1803 ( .A(n_1695), .B(n_1712), .Y(n_1803) );
NOR2xp33_ASAP7_75t_L g1815 ( .A(n_1695), .B(n_1816), .Y(n_1815) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1696), .B(n_1740), .Y(n_1739) );
NAND2xp5_ASAP7_75t_L g1746 ( .A(n_1696), .B(n_1747), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1696), .B(n_1707), .Y(n_1796) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1698), .Y(n_1760) );
OAI21xp5_ASAP7_75t_L g1848 ( .A1(n_1698), .A2(n_1849), .B(n_1850), .Y(n_1848) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
NAND2xp5_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1707), .Y(n_1700) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1701), .Y(n_1876) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
OR2x2_ASAP7_75t_L g1716 ( .A(n_1702), .B(n_1717), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1703), .B(n_1706), .Y(n_1702) );
INVx2_ASAP7_75t_SL g1737 ( .A(n_1703), .Y(n_1737) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1703), .Y(n_1748) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1705), .Y(n_1703) );
OR2x2_ASAP7_75t_L g1736 ( .A(n_1706), .B(n_1737), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1706), .B(n_1730), .Y(n_1743) );
NOR2xp33_ASAP7_75t_L g1762 ( .A(n_1706), .B(n_1763), .Y(n_1762) );
OAI22xp5_ASAP7_75t_L g1793 ( .A1(n_1706), .A2(n_1773), .B1(n_1794), .B2(n_1797), .Y(n_1793) );
NAND3xp33_ASAP7_75t_L g1832 ( .A(n_1706), .B(n_1723), .C(n_1833), .Y(n_1832) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1707), .Y(n_1721) );
NAND2xp5_ASAP7_75t_L g1828 ( .A(n_1707), .B(n_1829), .Y(n_1828) );
INVxp33_ASAP7_75t_SL g1708 ( .A(n_1709), .Y(n_1708) );
NOR2xp33_ASAP7_75t_SL g1709 ( .A(n_1710), .B(n_1714), .Y(n_1709) );
INVx2_ASAP7_75t_L g1734 ( .A(n_1710), .Y(n_1734) );
AOI222xp33_ASAP7_75t_L g1783 ( .A1(n_1711), .A2(n_1784), .B1(n_1785), .B2(n_1786), .C1(n_1788), .C2(n_1790), .Y(n_1783) );
NOR2xp33_ASAP7_75t_L g1819 ( .A(n_1711), .B(n_1798), .Y(n_1819) );
A2O1A1Ixp33_ASAP7_75t_L g1872 ( .A1(n_1711), .A2(n_1721), .B(n_1790), .C(n_1802), .Y(n_1872) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
A2O1A1Ixp33_ASAP7_75t_L g1873 ( .A1(n_1714), .A2(n_1785), .B(n_1813), .C(n_1874), .Y(n_1873) );
OAI21xp5_ASAP7_75t_SL g1715 ( .A1(n_1716), .A2(n_1719), .B(n_1724), .Y(n_1715) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1716), .Y(n_1868) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1718), .Y(n_1789) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1718), .B(n_1765), .Y(n_1806) );
AND2x2_ASAP7_75t_L g1808 ( .A(n_1718), .B(n_1726), .Y(n_1808) );
NAND2xp5_ASAP7_75t_L g1855 ( .A(n_1718), .B(n_1856), .Y(n_1855) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1722), .Y(n_1720) );
AOI221xp5_ASAP7_75t_L g1859 ( .A1(n_1722), .A2(n_1825), .B1(n_1860), .B2(n_1861), .C(n_1862), .Y(n_1859) );
NAND2xp5_ASAP7_75t_L g1724 ( .A(n_1723), .B(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1723), .Y(n_1768) );
AND2x2_ASAP7_75t_L g1852 ( .A(n_1723), .B(n_1747), .Y(n_1852) );
NAND2xp5_ASAP7_75t_L g1759 ( .A(n_1725), .B(n_1760), .Y(n_1759) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1725), .B(n_1775), .Y(n_1774) );
NAND2xp5_ASAP7_75t_L g1826 ( .A(n_1726), .B(n_1785), .Y(n_1826) );
INVx2_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
AOI21xp33_ASAP7_75t_L g1792 ( .A1(n_1727), .A2(n_1793), .B(n_1799), .Y(n_1792) );
INVxp67_ASAP7_75t_SL g1728 ( .A(n_1729), .Y(n_1728) );
NAND2xp5_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1731), .Y(n_1729) );
NOR2xp33_ASAP7_75t_L g1731 ( .A(n_1732), .B(n_1734), .Y(n_1731) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
OAI21xp33_ASAP7_75t_L g1754 ( .A1(n_1733), .A2(n_1755), .B(n_1756), .Y(n_1754) );
OAI211xp5_ASAP7_75t_SL g1735 ( .A1(n_1736), .A2(n_1738), .B(n_1742), .C(n_1754), .Y(n_1735) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1736), .Y(n_1861) );
INVx2_ASAP7_75t_L g1769 ( .A(n_1737), .Y(n_1769) );
AND2x2_ASAP7_75t_L g1851 ( .A(n_1737), .B(n_1852), .Y(n_1851) );
O2A1O1Ixp33_ASAP7_75t_SL g1862 ( .A1(n_1737), .A2(n_1804), .B(n_1863), .C(n_1864), .Y(n_1862) );
CKINVDCx14_ASAP7_75t_R g1738 ( .A(n_1739), .Y(n_1738) );
NAND2xp5_ASAP7_75t_L g1797 ( .A(n_1740), .B(n_1798), .Y(n_1797) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
OR2x2_ASAP7_75t_L g1804 ( .A(n_1741), .B(n_1768), .Y(n_1804) );
AOI211xp5_ASAP7_75t_L g1853 ( .A1(n_1741), .A2(n_1854), .B(n_1855), .C(n_1857), .Y(n_1853) );
AOI221xp5_ASAP7_75t_L g1742 ( .A1(n_1743), .A2(n_1744), .B1(n_1745), .B2(n_1748), .C(n_1749), .Y(n_1742) );
NOR2xp33_ASAP7_75t_L g1766 ( .A(n_1743), .B(n_1767), .Y(n_1766) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1743), .Y(n_1820) );
O2A1O1Ixp33_ASAP7_75t_L g1865 ( .A1(n_1744), .A2(n_1866), .B(n_1868), .C(n_1869), .Y(n_1865) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1746), .B(n_1765), .Y(n_1764) );
INVx2_ASAP7_75t_L g1765 ( .A(n_1748), .Y(n_1765) );
NAND2xp5_ASAP7_75t_L g1831 ( .A(n_1749), .B(n_1832), .Y(n_1831) );
INVx3_ASAP7_75t_L g1749 ( .A(n_1750), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1750 ( .A(n_1751), .B(n_1753), .Y(n_1750) );
HB1xp67_ASAP7_75t_L g1878 ( .A(n_1752), .Y(n_1878) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1755), .Y(n_1864) );
INVx2_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
INVxp67_ASAP7_75t_SL g1758 ( .A(n_1759), .Y(n_1758) );
O2A1O1Ixp33_ASAP7_75t_L g1761 ( .A1(n_1762), .A2(n_1766), .B(n_1769), .C(n_1770), .Y(n_1761) );
OAI31xp33_ASAP7_75t_L g1777 ( .A1(n_1762), .A2(n_1766), .A3(n_1778), .B(n_1781), .Y(n_1777) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1764), .Y(n_1763) );
AND2x2_ASAP7_75t_L g1788 ( .A(n_1765), .B(n_1789), .Y(n_1788) );
OR2x2_ASAP7_75t_L g1824 ( .A(n_1765), .B(n_1789), .Y(n_1824) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1767), .Y(n_1822) );
NAND2xp5_ASAP7_75t_L g1779 ( .A(n_1769), .B(n_1780), .Y(n_1779) );
O2A1O1Ixp33_ASAP7_75t_L g1770 ( .A1(n_1771), .A2(n_1773), .B(n_1774), .C(n_1776), .Y(n_1770) );
AOI21xp33_ASAP7_75t_L g1874 ( .A1(n_1771), .A2(n_1875), .B(n_1876), .Y(n_1874) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
NAND2xp5_ASAP7_75t_L g1842 ( .A(n_1775), .B(n_1843), .Y(n_1842) );
CKINVDCx14_ASAP7_75t_R g1870 ( .A(n_1775), .Y(n_1870) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1776), .Y(n_1785) );
AOI221xp5_ASAP7_75t_L g1845 ( .A1(n_1776), .A2(n_1808), .B1(n_1846), .B2(n_1848), .C(n_1853), .Y(n_1845) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
INVx1_ASAP7_75t_L g1863 ( .A(n_1781), .Y(n_1863) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1784), .Y(n_1875) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
AOI222xp33_ASAP7_75t_L g1834 ( .A1(n_1788), .A2(n_1823), .B1(n_1835), .B2(n_1836), .C1(n_1838), .C2(n_1840), .Y(n_1834) );
NAND5xp2_ASAP7_75t_L g1791 ( .A(n_1792), .B(n_1807), .C(n_1821), .D(n_1834), .E(n_1842), .Y(n_1791) );
INVx1_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
INVxp67_ASAP7_75t_SL g1854 ( .A(n_1796), .Y(n_1854) );
AOI21xp33_ASAP7_75t_L g1799 ( .A1(n_1800), .A2(n_1804), .B(n_1805), .Y(n_1799) );
INVx1_ASAP7_75t_L g1800 ( .A(n_1801), .Y(n_1800) );
INVx1_ASAP7_75t_L g1802 ( .A(n_1803), .Y(n_1802) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1804), .Y(n_1835) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
INVxp67_ASAP7_75t_SL g1812 ( .A(n_1813), .Y(n_1812) );
INVxp67_ASAP7_75t_L g1814 ( .A(n_1815), .Y(n_1814) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
HB1xp67_ASAP7_75t_L g1818 ( .A(n_1819), .Y(n_1818) );
AOI221xp5_ASAP7_75t_L g1821 ( .A1(n_1822), .A2(n_1823), .B1(n_1825), .B2(n_1827), .C(n_1831), .Y(n_1821) );
INVx1_ASAP7_75t_L g1823 ( .A(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1826), .Y(n_1825) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
INVx1_ASAP7_75t_L g1829 ( .A(n_1830), .Y(n_1829) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1837), .Y(n_1856) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1839), .Y(n_1838) );
INVxp67_ASAP7_75t_SL g1840 ( .A(n_1841), .Y(n_1840) );
NAND4xp25_ASAP7_75t_L g1844 ( .A(n_1845), .B(n_1859), .C(n_1865), .D(n_1873), .Y(n_1844) );
INVxp67_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1851), .Y(n_1850) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVx4_ASAP7_75t_L g1877 ( .A(n_1878), .Y(n_1877) );
HB1xp67_ASAP7_75t_L g1929 ( .A(n_1880), .Y(n_1929) );
NAND3xp33_ASAP7_75t_L g1880 ( .A(n_1881), .B(n_1903), .C(n_1912), .Y(n_1880) );
NOR2xp33_ASAP7_75t_L g1881 ( .A(n_1882), .B(n_1896), .Y(n_1881) );
INVx1_ASAP7_75t_L g1905 ( .A(n_1906), .Y(n_1905) );
INVx1_ASAP7_75t_L g1914 ( .A(n_1915), .Y(n_1914) );
CKINVDCx5p33_ASAP7_75t_R g1920 ( .A(n_1921), .Y(n_1920) );
BUFx3_ASAP7_75t_L g1924 ( .A(n_1925), .Y(n_1924) );
BUFx3_ASAP7_75t_L g1925 ( .A(n_1926), .Y(n_1925) );
INVxp33_ASAP7_75t_SL g1927 ( .A(n_1928), .Y(n_1927) );
INVx1_ASAP7_75t_L g1930 ( .A(n_1931), .Y(n_1930) );
INVx1_ASAP7_75t_L g1931 ( .A(n_1932), .Y(n_1931) );
INVx1_ASAP7_75t_L g1934 ( .A(n_1935), .Y(n_1934) );
endmodule