module real_jpeg_4940_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_0),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_0),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_1),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_1),
.Y(n_144)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_1),
.Y(n_363)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_1),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g460 ( 
.A(n_1),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_2),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_2),
.A2(n_53),
.B1(n_230),
.B2(n_313),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_2),
.A2(n_53),
.B1(n_290),
.B2(n_390),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_2),
.A2(n_53),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_3),
.Y(n_332)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_3),
.Y(n_336)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_5),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_6),
.A2(n_60),
.B1(n_348),
.B2(n_350),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_6),
.A2(n_60),
.B1(n_393),
.B2(n_395),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_6),
.A2(n_60),
.B1(n_440),
.B2(n_442),
.Y(n_439)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_9),
.A2(n_117),
.B1(n_277),
.B2(n_280),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_9),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_9),
.A2(n_255),
.B1(n_280),
.B2(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_9),
.A2(n_280),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_L g456 ( 
.A1(n_9),
.A2(n_280),
.B1(n_457),
.B2(n_459),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_10),
.Y(n_196)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_12),
.A2(n_86),
.B1(n_88),
.B2(n_91),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_12),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_12),
.A2(n_91),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_12),
.A2(n_91),
.B1(n_203),
.B2(n_222),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_12),
.A2(n_91),
.B1(n_287),
.B2(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_13),
.A2(n_162),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_13),
.A2(n_166),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_13),
.A2(n_43),
.B1(n_166),
.B2(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_13),
.A2(n_166),
.B1(n_362),
.B2(n_364),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_14),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_180)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_14),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_14),
.A2(n_124),
.B1(n_187),
.B2(n_254),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_14),
.A2(n_187),
.B1(n_368),
.B2(n_370),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_14),
.A2(n_57),
.B1(n_187),
.B2(n_408),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_15),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_15),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_15),
.A2(n_181),
.B1(n_210),
.B2(n_230),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_15),
.A2(n_69),
.B1(n_210),
.B2(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_15),
.A2(n_58),
.B1(n_132),
.B2(n_210),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_16),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_16),
.A2(n_98),
.B1(n_124),
.B2(n_127),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_16),
.A2(n_98),
.B1(n_130),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_16),
.A2(n_98),
.B1(n_119),
.B2(n_222),
.Y(n_387)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_18),
.A2(n_127),
.B1(n_156),
.B2(n_159),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_18),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_18),
.B(n_174),
.C(n_177),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_18),
.B(n_77),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_18),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_18),
.B(n_122),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_18),
.B(n_268),
.Y(n_267)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_536),
.B(n_539),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_145),
.B(n_535),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_137),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_27),
.B(n_137),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_128),
.C(n_134),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_28),
.A2(n_29),
.B1(n_531),
.B2(n_532),
.Y(n_530)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_61),
.C(n_99),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_30),
.B(n_523),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_47),
.B1(n_54),
.B2(n_56),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_31),
.A2(n_54),
.B1(n_56),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_31),
.A2(n_54),
.B1(n_129),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_31),
.A2(n_360),
.B(n_407),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_31),
.A2(n_54),
.B1(n_407),
.B2(n_428),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_31),
.A2(n_47),
.B1(n_54),
.B2(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_32),
.A2(n_358),
.B(n_359),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_32),
.B(n_361),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_32),
.A2(n_55),
.B(n_538),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_40),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.Y(n_40)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_42),
.Y(n_265)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_42),
.Y(n_272)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_44),
.Y(n_402)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_54),
.B(n_159),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_54),
.A2(n_428),
.B(n_461),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_55),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_55),
.B(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_61),
.A2(n_99),
.B1(n_100),
.B2(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_61),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_61)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_62),
.A2(n_92),
.B1(n_304),
.B2(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_62),
.A2(n_92),
.B1(n_400),
.B2(n_403),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_62),
.A2(n_85),
.B1(n_92),
.B2(n_512),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_77),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_72),
.B2(n_74),
.Y(n_63)
);

AOI32xp33_ASAP7_75t_L g283 ( 
.A1(n_64),
.A2(n_267),
.A3(n_284),
.B1(n_287),
.B2(n_289),
.Y(n_283)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_69),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_71),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_73),
.Y(n_293)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_76),
.Y(n_444)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_77),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g429 ( 
.A1(n_77),
.A2(n_135),
.B1(n_308),
.B2(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_77),
.A2(n_135),
.B1(n_438),
.B2(n_439),
.Y(n_437)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_81),
.Y(n_258)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_86),
.Y(n_370)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_92),
.B(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_92),
.A2(n_304),
.B(n_307),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_99),
.A2(n_100),
.B1(n_510),
.B2(n_511),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_99),
.B(n_507),
.C(n_510),
.Y(n_518)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_121),
.B(n_123),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_101),
.A2(n_155),
.B(n_160),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_101),
.A2(n_121),
.B1(n_207),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_101),
.A2(n_160),
.B(n_253),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_101),
.A2(n_121),
.B1(n_372),
.B2(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_102),
.B(n_161),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_102),
.A2(n_122),
.B1(n_389),
.B2(n_392),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_102),
.A2(n_122),
.B1(n_392),
.B2(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_102),
.A2(n_122),
.B1(n_413),
.B2(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_113),
.Y(n_291)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_114),
.A2(n_207),
.B(n_214),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_121),
.A2(n_214),
.B(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_123),
.Y(n_447)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_126),
.Y(n_373)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_126),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_128),
.B(n_134),
.Y(n_532)
);

OAI21xp33_ASAP7_75t_SL g358 ( 
.A1(n_131),
.A2(n_159),
.B(n_339),
.Y(n_358)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_135),
.A2(n_261),
.B(n_269),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_135),
.B(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_135),
.A2(n_269),
.B(n_474),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_137),
.B(n_537),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_137),
.B(n_537),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_138),
.Y(n_538)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_144),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_529),
.B(n_534),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_500),
.B(n_526),
.Y(n_146)
);

OAI311xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_376),
.A3(n_476),
.B1(n_494),
.C1(n_495),
.Y(n_147)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_318),
.B(n_375),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_295),
.B(n_317),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_247),
.B(n_294),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_217),
.B(n_246),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_178),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_153),
.B(n_178),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_169),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_154),
.A2(n_169),
.B1(n_170),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_154),
.Y(n_244)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_158),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_159),
.A2(n_191),
.B(n_197),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_SL g261 ( 
.A1(n_159),
.A2(n_262),
.B(n_266),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_159),
.B(n_330),
.Y(n_339)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_165),
.Y(n_416)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_204),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_205),
.C(n_216),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_191),
.B(n_197),
.Y(n_179)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_185),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_190),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_191),
.A2(n_342),
.B1(n_343),
.B2(n_346),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_191),
.A2(n_382),
.B1(n_383),
.B2(n_387),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_191),
.A2(n_385),
.B(n_387),
.Y(n_417)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_201),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_192),
.A2(n_235),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_192),
.A2(n_276),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_192),
.A2(n_347),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_200),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_200),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_215),
.B2(n_216),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_239),
.B(n_245),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_227),
.B(n_238),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_223),
.Y(n_351)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_237),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_237),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_234),
.B(n_236),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_232),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_275),
.B(n_281),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_243),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_249),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_273),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_259),
.B2(n_260),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_259),
.C(n_273),
.Y(n_296)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx5_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_257),
.Y(n_391)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_262),
.Y(n_404)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_265),
.Y(n_306)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_296),
.B(n_297),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_302),
.B2(n_316),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_301),
.C(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_309),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_310),
.C(n_311),
.Y(n_352)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_319),
.B(n_320),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_355),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_321)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_340),
.B2(n_341),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_324),
.B(n_340),
.Y(n_472)
);

OAI32xp33_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_328),
.A3(n_331),
.B1(n_333),
.B2(n_339),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_352),
.B(n_353),
.C(n_355),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_365),
.B2(n_374),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_356),
.B(n_366),
.C(n_371),
.Y(n_485)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_365),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_371),
.Y(n_365)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_367),
.Y(n_474)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

INVx11_ASAP7_75t_L g394 ( 
.A(n_373),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_462),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_SL g495 ( 
.A1(n_377),
.A2(n_462),
.B(n_496),
.C(n_499),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_431),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_378),
.B(n_431),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_410),
.C(n_419),
.Y(n_378)
);

FAx1_ASAP7_75t_SL g475 ( 
.A(n_379),
.B(n_410),
.CI(n_419),
.CON(n_475),
.SN(n_475)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_398),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_399),
.C(n_406),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_388),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_381),
.B(n_388),
.Y(n_468)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx8_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

INVx8_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_406),
.Y(n_398)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_400),
.Y(n_430)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_417),
.B2(n_418),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_417),
.Y(n_451)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_417),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_417),
.A2(n_418),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_417),
.A2(n_451),
.B(n_454),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_426),
.C(n_429),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_420),
.B(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_421),
.B(n_423),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_426),
.A2(n_427),
.B1(n_429),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_429),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_432),
.B(n_435),
.C(n_449),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_449),
.B2(n_450),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_445),
.B(n_448),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_446),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_439),
.Y(n_512)
);

INVx4_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_448),
.B(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_448),
.B(n_503),
.C(n_505),
.Y(n_525)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_461),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_456),
.Y(n_508)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_475),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_475),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_468),
.C(n_469),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_464),
.A2(n_465),
.B1(n_468),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_487),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_472),
.C(n_473),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_470),
.A2(n_471),
.B1(n_473),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_475),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_489),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_478),
.A2(n_497),
.B(n_498),
.Y(n_496)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_486),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_486),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_483),
.C(n_485),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_492),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_483),
.A2(n_484),
.B1(n_485),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_485),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_491),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_515),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_514),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_502),
.B(n_514),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_507),
.B1(n_509),
.B2(n_513),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_506),
.A2(n_507),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_506),
.B(n_517),
.C(n_521),
.Y(n_533)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_509),
.Y(n_513)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_515),
.A2(n_527),
.B(n_528),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_516),
.B(n_525),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_525),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_518),
.B1(n_519),
.B2(n_520),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_533),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_533),
.Y(n_534)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);


endmodule