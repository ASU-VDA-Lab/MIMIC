module fake_jpeg_16582_n_204 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_1),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_42),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_0),
.CON(n_36),
.SN(n_36)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_40),
.B(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_18),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_53),
.B1(n_55),
.B2(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_50),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_3),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_5),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_21),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_31),
.B1(n_30),
.B2(n_20),
.Y(n_82)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_57),
.Y(n_64)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_17),
.B(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_28),
.B(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_71),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_R g115 ( 
.A(n_69),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_15),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_15),
.Y(n_77)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_83),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_20),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_31),
.B1(n_30),
.B2(n_24),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_80),
.B1(n_66),
.B2(n_75),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_16),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_42),
.B(n_29),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_94),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_87),
.B1(n_82),
.B2(n_66),
.Y(n_119)
);

NOR2xp67_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_14),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_76),
.Y(n_131)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_8),
.B(n_50),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_102),
.B(n_68),
.Y(n_134)
);

AO21x2_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_37),
.B(n_47),
.Y(n_102)
);

OAI22x1_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_34),
.B1(n_61),
.B2(n_71),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_102),
.B1(n_99),
.B2(n_109),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_34),
.C(n_72),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_112),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_34),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_62),
.B(n_75),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_83),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_61),
.CI(n_89),
.CON(n_113),
.SN(n_113)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_112),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_70),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_127),
.B1(n_136),
.B2(n_137),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_129),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_126),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_64),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_139),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_106),
.B(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_68),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_141),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_68),
.B1(n_76),
.B2(n_104),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_102),
.B1(n_106),
.B2(n_95),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_93),
.B(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_103),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_113),
.C(n_108),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_148),
.C(n_144),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_106),
.B(n_92),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_152),
.B1(n_120),
.B2(n_149),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_107),
.C(n_100),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_96),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_139),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_101),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_138),
.B1(n_130),
.B2(n_120),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_116),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_134),
.B1(n_131),
.B2(n_138),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_142),
.A3(n_140),
.B1(n_119),
.B2(n_132),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_165),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_143),
.C(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_128),
.C(n_137),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_121),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_170),
.B(n_147),
.Y(n_184)
);

OAI322xp33_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_154),
.A3(n_155),
.B1(n_149),
.B2(n_161),
.C1(n_122),
.C2(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_169),
.B(n_172),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_134),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_181),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_161),
.B1(n_160),
.B2(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_182),
.Y(n_187)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_165),
.B(n_166),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_180),
.Y(n_194)
);

OAI321xp33_ASAP7_75t_L g188 ( 
.A1(n_179),
.A2(n_172),
.A3(n_167),
.B1(n_170),
.B2(n_153),
.C(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_190),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_180),
.C(n_184),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_185),
.B(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_192),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_189),
.A2(n_178),
.B1(n_183),
.B2(n_187),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_197),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_195),
.A2(n_193),
.B(n_196),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.C(n_198),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_194),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule