module fake_aes_5721_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_5), .B(n_6), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_1), .B(n_8), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_SL g17 ( .A(n_13), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_18), .B(n_12), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
INVx2_ASAP7_75t_SL g21 ( .A(n_20), .Y(n_21) );
AO31x2_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_15), .A3(n_16), .B(n_11), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
AOI211xp5_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_17), .B(n_14), .C(n_16), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OAI21xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_24), .B(n_18), .Y(n_27) );
AOI221xp5_ASAP7_75t_SL g28 ( .A1(n_25), .A2(n_18), .B1(n_12), .B2(n_22), .C(n_14), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
NOR2xp33_ASAP7_75t_L g30 ( .A(n_28), .B(n_0), .Y(n_30) );
AND3x4_ASAP7_75t_L g31 ( .A(n_30), .B(n_2), .C(n_3), .Y(n_31) );
AOI21xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_12), .B(n_22), .Y(n_32) );
CKINVDCx20_ASAP7_75t_R g33 ( .A(n_31), .Y(n_33) );
AOI322xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_2), .A3(n_3), .B1(n_32), .B2(n_7), .C1(n_9), .C2(n_4), .Y(n_34) );
endmodule