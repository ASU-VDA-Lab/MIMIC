module fake_jpeg_26393_n_285 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_285);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_32),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_26),
.Y(n_48)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_25),
.B1(n_18),
.B2(n_13),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_35),
.B1(n_33),
.B2(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_48),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_57),
.Y(n_79)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_35),
.B1(n_33),
.B2(n_25),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_59),
.B1(n_62),
.B2(n_36),
.Y(n_77)
);

OAI22x1_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_30),
.B1(n_39),
.B2(n_23),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_27),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_35),
.B1(n_25),
.B2(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_18),
.B1(n_13),
.B2(n_20),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_34),
.B1(n_36),
.B2(n_28),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_67),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_68),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_75),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_77),
.B1(n_80),
.B2(n_45),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_49),
.B1(n_34),
.B2(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_32),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_49),
.B1(n_40),
.B2(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_87),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_30),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_30),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_41),
.B1(n_45),
.B2(n_28),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_56),
.A3(n_66),
.B1(n_58),
.B2(n_65),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_97),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_68),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_66),
.C(n_62),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_98),
.C(n_102),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_55),
.C(n_59),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_41),
.C(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_89),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_12),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_108),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_64),
.B(n_67),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_74),
.B(n_70),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_16),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_85),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_22),
.C(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_16),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_112),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_87),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_119),
.B(n_101),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_105),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_120),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_77),
.B(n_85),
.C(n_89),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_126),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_50),
.B1(n_71),
.B2(n_75),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_99),
.B1(n_50),
.B2(n_82),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_64),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_107),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_140),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_51),
.B(n_19),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_19),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_108),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_125),
.B(n_119),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_149),
.B1(n_127),
.B2(n_116),
.Y(n_165)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_153),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_151),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_98),
.C(n_90),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_156),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_111),
.B1(n_118),
.B2(n_128),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_104),
.C(n_11),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_155),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_97),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_97),
.B1(n_82),
.B2(n_83),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_121),
.B1(n_63),
.B2(n_86),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_83),
.C(n_60),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_63),
.B1(n_86),
.B2(n_21),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_110),
.B1(n_113),
.B2(n_112),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_158),
.B(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_174),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_119),
.B(n_111),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_168),
.B(n_170),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_144),
.B1(n_149),
.B2(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_53),
.B1(n_14),
.B2(n_20),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_176),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_115),
.B(n_131),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_131),
.B(n_121),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_171),
.A2(n_53),
.B1(n_45),
.B2(n_26),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_21),
.B(n_11),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_10),
.C(n_9),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_156),
.B(n_17),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_167),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_141),
.B1(n_138),
.B2(n_139),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_199),
.B1(n_22),
.B2(n_19),
.Y(n_214)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_168),
.C(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_194),
.C(n_196),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_138),
.C(n_51),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_195),
.A2(n_166),
.B1(n_173),
.B2(n_172),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_26),
.C(n_14),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_14),
.B(n_15),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_202),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_14),
.C(n_31),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_161),
.C(n_182),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_169),
.B1(n_176),
.B2(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_215),
.C(n_217),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_193),
.B(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_158),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_211),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_16),
.B1(n_20),
.B2(n_17),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_212),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_216),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_14),
.C(n_31),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_16),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_31),
.C(n_19),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_31),
.C(n_19),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_39),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_23),
.B1(n_15),
.B2(n_3),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_23),
.B1(n_15),
.B2(n_3),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_227),
.B(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_209),
.B(n_213),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_230),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_197),
.CI(n_207),
.CON(n_224),
.SN(n_224)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_200),
.B(n_196),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_200),
.B(n_199),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_229),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_183),
.B(n_185),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_197),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_233),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_201),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_226),
.A2(n_215),
.B1(n_217),
.B2(n_219),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_225),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_218),
.B(n_15),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_30),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_31),
.C(n_23),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_244),
.C(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_1),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_23),
.C(n_30),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_1),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_258),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_252),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_228),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_227),
.C(n_225),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.C(n_4),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_224),
.C(n_231),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_1),
.B(n_2),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_247),
.B(n_248),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_264),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_268),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_237),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_251),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_4),
.C2(n_30),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_4),
.C(n_5),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_269),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_256),
.B1(n_253),
.B2(n_254),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_274),
.B(n_265),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_6),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_270),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_272),
.A2(n_267),
.B(n_7),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_278),
.A2(n_275),
.B(n_7),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_279),
.A2(n_280),
.B(n_276),
.C(n_7),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_281),
.B(n_6),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_6),
.C(n_8),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_8),
.B(n_276),
.Y(n_285)
);


endmodule