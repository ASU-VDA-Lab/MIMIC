module fake_jpeg_30478_n_29 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

OR2x2_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_7),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_8),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_0),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.C(n_21),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_14),
.B1(n_18),
.B2(n_10),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_23),
.C(n_24),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_11),
.A2(n_9),
.B1(n_18),
.B2(n_16),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_9),
.A2(n_15),
.B(n_13),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_26),
.C(n_22),
.Y(n_29)
);


endmodule