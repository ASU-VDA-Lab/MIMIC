module fake_jpeg_6788_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_38),
.B(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_45),
.B(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_13),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_12),
.B(n_1),
.C(n_3),
.Y(n_103)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_54),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_55),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_60),
.Y(n_107)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_20),
.B1(n_22),
.B2(n_36),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_63),
.A2(n_67),
.B1(n_90),
.B2(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_22),
.B1(n_20),
.B2(n_28),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_92),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_20),
.B1(n_36),
.B2(n_18),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_20),
.B1(n_18),
.B2(n_34),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_78),
.B1(n_87),
.B2(n_97),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_70),
.Y(n_109)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_73),
.Y(n_122)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_18),
.B1(n_35),
.B2(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_93),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_34),
.Y(n_84)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_35),
.B1(n_17),
.B2(n_29),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_55),
.A2(n_17),
.B1(n_31),
.B2(n_34),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_94),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_43),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_43),
.A2(n_31),
.B1(n_21),
.B2(n_32),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_41),
.B(n_0),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_32),
.B1(n_23),
.B2(n_30),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_41),
.B(n_32),
.C(n_23),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_0),
.C(n_1),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_24),
.B1(n_30),
.B2(n_32),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_30),
.B1(n_23),
.B2(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_0),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_33),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_119),
.Y(n_145)
);

OR2x4_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_33),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_125),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_58),
.A2(n_23),
.B1(n_25),
.B2(n_33),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_92),
.B1(n_99),
.B2(n_66),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_123),
.Y(n_163)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_25),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_127),
.Y(n_148)
);

OR2x2_ASAP7_75t_SL g125 ( 
.A(n_65),
.B(n_12),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_132),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_19),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_87),
.C(n_93),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_131),
.B1(n_61),
.B2(n_7),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_60),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_103),
.B1(n_83),
.B2(n_98),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_82),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

OR2x2_ASAP7_75t_SL g134 ( 
.A(n_65),
.B(n_5),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_134),
.B(n_135),
.Y(n_174)
);

OR2x2_ASAP7_75t_SL g135 ( 
.A(n_82),
.B(n_102),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_117),
.C(n_137),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_78),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_144),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_141),
.B1(n_146),
.B2(n_147),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_95),
.B1(n_91),
.B2(n_59),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_124),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_99),
.B1(n_76),
.B2(n_72),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_105),
.A2(n_86),
.B1(n_62),
.B2(n_71),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_158),
.B(n_161),
.C(n_133),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_77),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_157),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

INVx4_ASAP7_75t_SL g208 ( 
.A(n_155),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_81),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_75),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_105),
.A2(n_68),
.B1(n_73),
.B2(n_61),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_75),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_112),
.A2(n_100),
.B1(n_96),
.B2(n_89),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_121),
.B(n_6),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_6),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_117),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_112),
.A2(n_89),
.B1(n_9),
.B2(n_10),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_173),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_8),
.Y(n_171)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_8),
.Y(n_172)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_9),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_128),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_191),
.C(n_199),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_141),
.B1(n_161),
.B2(n_154),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_108),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_183),
.B(n_171),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_108),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_151),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_159),
.A2(n_120),
.B(n_115),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_190),
.B(n_198),
.Y(n_221)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_194),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_137),
.B(n_119),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_196),
.Y(n_230)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_9),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_139),
.A2(n_110),
.B(n_119),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_126),
.C(n_110),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_142),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_126),
.C(n_109),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_146),
.C(n_170),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_148),
.B(n_9),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_209),
.B(n_143),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_214),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_190),
.B1(n_187),
.B2(n_182),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_232),
.B1(n_180),
.B2(n_182),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_140),
.C(n_166),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_152),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_235),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_223),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_203),
.B1(n_198),
.B2(n_179),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_176),
.B(n_192),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_226),
.C(n_236),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_SL g225 ( 
.A1(n_181),
.A2(n_157),
.B(n_166),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_207),
.B(n_184),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_148),
.C(n_174),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_228),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_150),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_185),
.A2(n_174),
.B1(n_167),
.B2(n_123),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_177),
.A2(n_186),
.B(n_188),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_186),
.B(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_172),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_178),
.B(n_181),
.C(n_199),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_237),
.A2(n_242),
.B(n_251),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_212),
.A2(n_179),
.B1(n_205),
.B2(n_227),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_250),
.B1(n_254),
.B2(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

OAI32xp33_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_233),
.A3(n_221),
.B1(n_222),
.B2(n_210),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_230),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_184),
.B(n_195),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_212),
.Y(n_246)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_209),
.B1(n_206),
.B2(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_257),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_217),
.A2(n_193),
.B(n_195),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_256),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_189),
.B1(n_194),
.B2(n_106),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_217),
.A2(n_168),
.B(n_175),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_236),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_270),
.Y(n_286)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_269),
.B1(n_273),
.B2(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_265),
.Y(n_276)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_216),
.C(n_226),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_248),
.C(n_256),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_239),
.A2(n_230),
.B1(n_211),
.B2(n_235),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_244),
.A2(n_211),
.B1(n_231),
.B2(n_162),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_197),
.C(n_10),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_274),
.A2(n_245),
.B(n_258),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_250),
.B1(n_237),
.B2(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_283),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_249),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_287),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_251),
.B(n_247),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_265),
.B(n_263),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_243),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_248),
.C(n_253),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_284),
.B(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_272),
.B(n_271),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_296),
.B(n_276),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_288),
.A2(n_260),
.B1(n_271),
.B2(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_276),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_299),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_287),
.C(n_289),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_277),
.A3(n_285),
.B1(n_281),
.B2(n_286),
.C1(n_279),
.C2(n_280),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_304),
.C(n_306),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_281),
.C(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

AOI31xp33_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_269),
.A3(n_286),
.B(n_278),
.Y(n_308)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_310),
.A3(n_290),
.B1(n_243),
.B2(n_245),
.C(n_297),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_290),
.A3(n_298),
.B1(n_293),
.B2(n_294),
.C1(n_299),
.C2(n_280),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_261),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_284),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_312),
.A2(n_313),
.B(n_315),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_267),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_252),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_306),
.C(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_257),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_321),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_313),
.A3(n_318),
.B1(n_317),
.B2(n_297),
.C1(n_304),
.C2(n_262),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_322),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_323),
.Y(n_325)
);


endmodule