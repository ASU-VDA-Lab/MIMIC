module fake_jpeg_8028_n_95 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_1),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_3),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_43),
.B1(n_37),
.B2(n_47),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_43),
.B1(n_37),
.B2(n_45),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_33),
.B1(n_5),
.B2(n_4),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_4),
.CON(n_66),
.SN(n_66)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_69),
.A3(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_10),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_24),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_70),
.B1(n_67),
.B2(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_83),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_72),
.B(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_85),
.B(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_73),
.B(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_82),
.B(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_80),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_90),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_78),
.B1(n_79),
.B2(n_60),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_26),
.B(n_27),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_29),
.Y(n_95)
);


endmodule