module fake_jpeg_8051_n_226 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_26),
.B1(n_27),
.B2(n_25),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_53),
.B1(n_38),
.B2(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_30),
.B1(n_17),
.B2(n_29),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_33),
.B(n_27),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_51),
.B(n_20),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_26),
.B1(n_27),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_56),
.B1(n_20),
.B2(n_17),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_26),
.B1(n_20),
.B2(n_29),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_26),
.B1(n_15),
.B2(n_24),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_29),
.B1(n_14),
.B2(n_17),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_63),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_75),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_2),
.Y(n_62)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_2),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_72),
.Y(n_86)
);

INVxp67_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_36),
.B1(n_40),
.B2(n_57),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_63),
.B(n_59),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_65),
.B(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_38),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_80),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_101),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_36),
.B(n_48),
.C(n_46),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_83),
.A2(n_88),
.B(n_90),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_76),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_45),
.C(n_31),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_14),
.C(n_19),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_45),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_57),
.B1(n_55),
.B2(n_31),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_55),
.B1(n_31),
.B2(n_34),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_28),
.B(n_21),
.C(n_16),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_70),
.B(n_28),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_79),
.Y(n_108)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_77),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_67),
.B1(n_14),
.B2(n_19),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_107),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_79),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_67),
.B1(n_64),
.B2(n_24),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_116),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_82),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_88),
.C(n_84),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_123),
.B(n_103),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_21),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_124),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_121),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_19),
.B1(n_23),
.B2(n_15),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_24),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_16),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_2),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_98),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_119),
.B(n_116),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_90),
.B(n_105),
.Y(n_130)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_136),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_124),
.C(n_117),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_103),
.B(n_98),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_23),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_150),
.C(n_154),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_115),
.C(n_112),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_114),
.C(n_106),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_110),
.B1(n_91),
.B2(n_111),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_133),
.B1(n_135),
.B2(n_147),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_138),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_91),
.B1(n_110),
.B2(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_158),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_107),
.B1(n_120),
.B2(n_81),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_123),
.B1(n_92),
.B2(n_87),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_99),
.C(n_104),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_131),
.C(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_162),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_127),
.B(n_93),
.C(n_99),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_134),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_137),
.B(n_133),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_156),
.B(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_168),
.B1(n_178),
.B2(n_150),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_145),
.A3(n_137),
.B1(n_144),
.B2(n_139),
.C1(n_134),
.C2(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_176),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_174),
.C(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_164),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_149),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_162),
.B1(n_155),
.B2(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_184),
.B1(n_175),
.B2(n_167),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_177),
.B(n_152),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_186),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_190),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_163),
.B1(n_138),
.B2(n_143),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_174),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_131),
.B(n_102),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_191),
.B(n_196),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_23),
.B1(n_15),
.B2(n_5),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_23),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_172),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_171),
.C(n_186),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_189),
.C(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_101),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_199),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_171),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_3),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_206),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_190),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_193),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_207),
.B(n_6),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_6),
.B(n_7),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_213),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_212),
.B(n_202),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_197),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_193),
.B1(n_8),
.B2(n_9),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_205),
.C(n_208),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_214),
.B(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_12),
.C(n_8),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_212),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_10),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_220),
.Y(n_226)
);


endmodule