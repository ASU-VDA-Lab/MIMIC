module fake_netlist_6_1776_n_788 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_788);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_788;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_736;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_97),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_37),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_18),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_106),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_75),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_65),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_1),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_10),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_99),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_35),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_118),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_33),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_41),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_10),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_30),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_72),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_42),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_67),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_55),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_121),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_112),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_85),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_61),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_14),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_49),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_48),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_138),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_44),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_63),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_113),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_93),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_19),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_77),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_31),
.B(n_54),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_12),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_71),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_8),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_89),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_78),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

OAI22x1_ASAP7_75t_SL g212 ( 
.A1(n_163),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

BUFx8_ASAP7_75t_SL g213 ( 
.A(n_174),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_189),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_4),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_5),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_179),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_6),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_17),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_159),
.B(n_6),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_179),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_171),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_167),
.Y(n_240)
);

OAI21x1_ASAP7_75t_L g241 ( 
.A1(n_169),
.A2(n_178),
.B(n_176),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

INVxp33_ASAP7_75t_SL g243 ( 
.A(n_156),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_160),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_161),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_242),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_213),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_252),
.Y(n_258)
);

NOR2x1p5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_168),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_244),
.Y(n_264)
);

BUFx16f_ASAP7_75t_R g265 ( 
.A(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_233),
.B(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_R g268 ( 
.A(n_249),
.B(n_157),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_R g269 ( 
.A(n_249),
.B(n_183),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_243),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_250),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_250),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_250),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_250),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_228),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_R g279 ( 
.A(n_249),
.B(n_170),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_239),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_233),
.B(n_172),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_239),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_216),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_196),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_251),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_217),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_173),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_251),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_222),
.A2(n_202),
.B(n_204),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_221),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_251),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_248),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_219),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_284),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_220),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_231),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_287),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_241),
.B(n_231),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_287),
.B(n_298),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_224),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_SL g313 ( 
.A(n_266),
.B(n_268),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_269),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_274),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_286),
.B(n_231),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_293),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_262),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_281),
.B(n_224),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_290),
.B(n_231),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_235),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_295),
.B(n_223),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_296),
.B(n_263),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_283),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_259),
.B(n_224),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_260),
.B(n_223),
.C(n_230),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_L g333 ( 
.A(n_279),
.B(n_180),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_270),
.B(n_248),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_254),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_264),
.B(n_225),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_256),
.B(n_238),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

NAND3xp33_ASAP7_75t_L g342 ( 
.A(n_278),
.B(n_248),
.C(n_225),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_225),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_257),
.B(n_181),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_255),
.Y(n_348)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_257),
.A2(n_241),
.B(n_226),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_256),
.B(n_184),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_L g352 ( 
.A(n_301),
.B(n_186),
.Y(n_352)
);

BUFx6f_ASAP7_75t_SL g353 ( 
.A(n_265),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_253),
.B(n_235),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_258),
.B(n_247),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_258),
.B(n_247),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_284),
.B(n_210),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_258),
.B(n_247),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_258),
.B(n_246),
.Y(n_361)
);

NOR3xp33_ASAP7_75t_L g362 ( 
.A(n_266),
.B(n_219),
.C(n_214),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_284),
.B(n_210),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_287),
.B(n_188),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_258),
.B(n_246),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_258),
.B(n_246),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_361),
.A2(n_211),
.B(n_234),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_362),
.A2(n_246),
.B1(n_200),
.B2(n_236),
.Y(n_368)
);

NAND2xp33_ASAP7_75t_L g369 ( 
.A(n_306),
.B(n_190),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_304),
.B(n_246),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_359),
.Y(n_371)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_316),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_362),
.A2(n_236),
.B1(n_214),
.B2(n_226),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_7),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_236),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_312),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_303),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_191),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_360),
.A2(n_212),
.B1(n_195),
.B2(n_198),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_355),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_192),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_199),
.Y(n_383)
);

AND2x6_ASAP7_75t_SL g384 ( 
.A(n_330),
.B(n_344),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_303),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

BUFx12f_ASAP7_75t_SL g387 ( 
.A(n_363),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_316),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

BUFx2_ASAP7_75t_SL g391 ( 
.A(n_307),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_212),
.Y(n_392)
);

INVx8_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_356),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_R g395 ( 
.A(n_313),
.B(n_20),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_211),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_345),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_322),
.B(n_211),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_211),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_334),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_305),
.B(n_9),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_302),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_322),
.B(n_21),
.Y(n_407)
);

NOR3xp33_ASAP7_75t_SL g408 ( 
.A(n_332),
.B(n_11),
.C(n_12),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_315),
.B(n_211),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_349),
.A2(n_234),
.B1(n_232),
.B2(n_227),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_305),
.B(n_13),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_344),
.B(n_227),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_323),
.B(n_311),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_346),
.B(n_13),
.Y(n_414)
);

BUFx4f_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_317),
.A2(n_234),
.B1(n_232),
.B2(n_227),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_316),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_330),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_311),
.B(n_227),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_342),
.B(n_22),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_323),
.B(n_227),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_324),
.B(n_232),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_327),
.A2(n_234),
.B1(n_232),
.B2(n_16),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_328),
.B(n_23),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_349),
.A2(n_234),
.B1(n_232),
.B2(n_16),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_314),
.B(n_14),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_320),
.B(n_24),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_310),
.B(n_15),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_340),
.A2(n_15),
.B1(n_152),
.B2(n_26),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_343),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_321),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_329),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_339),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_339),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_387),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_436),
.B(n_335),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_309),
.B(n_333),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_381),
.A2(n_352),
.B1(n_337),
.B2(n_364),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_419),
.B(n_347),
.Y(n_442)
);

NAND2x1p5_ASAP7_75t_L g443 ( 
.A(n_371),
.B(n_351),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_372),
.A2(n_309),
.B(n_32),
.Y(n_444)
);

AND2x6_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_29),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_381),
.A2(n_353),
.B1(n_36),
.B2(n_38),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_375),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_376),
.B(n_34),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_353),
.B1(n_40),
.B2(n_43),
.Y(n_451)
);

NOR2x1_ASAP7_75t_L g452 ( 
.A(n_391),
.B(n_39),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_372),
.A2(n_45),
.B(n_46),
.Y(n_453)
);

NOR2x1_ASAP7_75t_R g454 ( 
.A(n_403),
.B(n_47),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_377),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_379),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_SL g457 ( 
.A1(n_429),
.A2(n_53),
.B(n_56),
.C(n_57),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_388),
.B(n_58),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_370),
.A2(n_59),
.B(n_60),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_423),
.B(n_62),
.Y(n_461)
);

OAI21xp33_ASAP7_75t_L g462 ( 
.A1(n_374),
.A2(n_64),
.B(n_66),
.Y(n_462)
);

O2A1O1Ixp33_ASAP7_75t_SL g463 ( 
.A1(n_431),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_421),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_397),
.B(n_412),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_79),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_410),
.A2(n_402),
.B(n_396),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_80),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_426),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_SL g471 ( 
.A(n_417),
.B(n_86),
.Y(n_471)
);

AOI21xp33_ASAP7_75t_L g472 ( 
.A1(n_406),
.A2(n_87),
.B(n_88),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_418),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_426),
.B(n_90),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_R g475 ( 
.A(n_384),
.B(n_91),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_386),
.Y(n_476)
);

AOI21x1_ASAP7_75t_L g477 ( 
.A1(n_409),
.A2(n_92),
.B(n_94),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_382),
.B(n_95),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_384),
.B(n_96),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_422),
.A2(n_98),
.B(n_100),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_383),
.B(n_101),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_417),
.A2(n_102),
.B(n_104),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_405),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_415),
.B(n_105),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_SL g486 ( 
.A(n_417),
.B(n_111),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_415),
.B(n_115),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_433),
.A2(n_368),
.B1(n_407),
.B2(n_378),
.Y(n_488)
);

OR2x2_ASAP7_75t_SL g489 ( 
.A(n_411),
.B(n_117),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_378),
.B(n_119),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_434),
.B(n_120),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_393),
.B(n_435),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_393),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_450),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_440),
.A2(n_430),
.B(n_389),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_465),
.Y(n_496)
);

AO21x2_ASAP7_75t_L g497 ( 
.A1(n_468),
.A2(n_424),
.B(n_420),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_473),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_438),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_455),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_476),
.Y(n_501)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_475),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_437),
.A2(n_400),
.B(n_428),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_444),
.A2(n_404),
.B(n_389),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_447),
.Y(n_507)
);

AO21x2_ASAP7_75t_L g508 ( 
.A1(n_488),
.A2(n_401),
.B(n_395),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_491),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_448),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_484),
.B(n_380),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_439),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_491),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_458),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_467),
.Y(n_516)
);

CKINVDCx12_ASAP7_75t_R g517 ( 
.A(n_454),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_485),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_490),
.A2(n_404),
.B(n_385),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_460),
.B(n_385),
.Y(n_520)
);

INVx5_ASAP7_75t_SL g521 ( 
.A(n_493),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_449),
.A2(n_416),
.B(n_367),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_445),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_478),
.A2(n_425),
.B(n_369),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_471),
.B(n_380),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_482),
.A2(n_408),
.B(n_123),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_459),
.A2(n_122),
.B(n_124),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_489),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_481),
.A2(n_126),
.B(n_127),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_445),
.Y(n_530)
);

AO21x2_ASAP7_75t_L g531 ( 
.A1(n_457),
.A2(n_392),
.B(n_130),
.Y(n_531)
);

AOI22x1_ASAP7_75t_L g532 ( 
.A1(n_487),
.A2(n_432),
.B1(n_132),
.B2(n_133),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_445),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_466),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_474),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_462),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_453),
.A2(n_129),
.B(n_135),
.Y(n_538)
);

INVx6_ASAP7_75t_L g539 ( 
.A(n_492),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_443),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_486),
.B(n_136),
.Y(n_541)
);

AOI22x1_ASAP7_75t_L g542 ( 
.A1(n_483),
.A2(n_432),
.B1(n_140),
.B2(n_141),
.Y(n_542)
);

INVx6_ASAP7_75t_L g543 ( 
.A(n_509),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_533),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_507),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_441),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_511),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_530),
.B(n_464),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_498),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_528),
.A2(n_451),
.B1(n_479),
.B2(n_469),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_509),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_506),
.A2(n_461),
.B(n_456),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_494),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_SL g554 ( 
.A(n_509),
.B(n_442),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_498),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_509),
.Y(n_556)
);

OA21x2_ASAP7_75t_L g557 ( 
.A1(n_519),
.A2(n_472),
.B(n_464),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_500),
.Y(n_558)
);

BUFx12f_ASAP7_75t_L g559 ( 
.A(n_499),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_535),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_501),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_510),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_519),
.A2(n_452),
.B(n_470),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_532),
.A2(n_446),
.B1(n_463),
.B2(n_144),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_512),
.A2(n_139),
.B1(n_143),
.B2(n_146),
.Y(n_565)
);

OAI21x1_ASAP7_75t_SL g566 ( 
.A1(n_530),
.A2(n_147),
.B(n_148),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_513),
.B(n_496),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_514),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_503),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_514),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_510),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

OAI22xp33_ASAP7_75t_L g573 ( 
.A1(n_515),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_520),
.Y(n_574)
);

OAI21x1_ASAP7_75t_SL g575 ( 
.A1(n_523),
.A2(n_534),
.B(n_504),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_539),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_505),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_537),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_512),
.A2(n_542),
.B1(n_525),
.B2(n_539),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_539),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_520),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_516),
.B(n_536),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_504),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_536),
.B(n_540),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_538),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_558),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_567),
.B(n_502),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_550),
.A2(n_524),
.B(n_526),
.Y(n_589)
);

OAI21xp33_ASAP7_75t_SL g590 ( 
.A1(n_567),
.A2(n_526),
.B(n_524),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_547),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_SL g592 ( 
.A(n_579),
.B(n_525),
.C(n_499),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_502),
.Y(n_593)
);

NOR2x1p5_ASAP7_75t_L g594 ( 
.A(n_559),
.B(n_536),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_558),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_547),
.B(n_536),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_576),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_546),
.A2(n_521),
.B1(n_541),
.B2(n_518),
.Y(n_598)
);

NOR3xp33_ASAP7_75t_SL g599 ( 
.A(n_573),
.B(n_517),
.C(n_518),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_R g600 ( 
.A(n_545),
.B(n_517),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_582),
.B(n_521),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_553),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_546),
.B(n_518),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_559),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_577),
.A2(n_495),
.B(n_527),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_R g606 ( 
.A(n_545),
.B(n_521),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_583),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_R g608 ( 
.A(n_576),
.B(n_508),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_580),
.Y(n_609)
);

OAI21xp33_ASAP7_75t_L g610 ( 
.A1(n_564),
.A2(n_541),
.B(n_527),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_580),
.B(n_508),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_553),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_R g613 ( 
.A(n_546),
.B(n_495),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_SL g614 ( 
.A(n_565),
.B(n_531),
.C(n_508),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_R g615 ( 
.A(n_544),
.B(n_531),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_583),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_560),
.B(n_529),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_SL g618 ( 
.A1(n_578),
.A2(n_529),
.B(n_538),
.C(n_497),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_585),
.B(n_522),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_551),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_551),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_543),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_R g623 ( 
.A(n_544),
.B(n_522),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_561),
.Y(n_624)
);

AO21x1_ASAP7_75t_L g625 ( 
.A1(n_548),
.A2(n_578),
.B(n_572),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_568),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_569),
.B(n_570),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_548),
.A2(n_569),
.B1(n_544),
.B2(n_568),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_570),
.B(n_555),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_543),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_543),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_549),
.B(n_555),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_R g633 ( 
.A(n_557),
.B(n_581),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_575),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_634),
.B(n_581),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_611),
.B(n_584),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_602),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_619),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_612),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_627),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_624),
.B(n_571),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_587),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_629),
.B(n_571),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_595),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_592),
.A2(n_554),
.B1(n_548),
.B2(n_566),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_614),
.A2(n_556),
.B(n_574),
.Y(n_646)
);

AOI21xp33_ASAP7_75t_SL g647 ( 
.A1(n_604),
.A2(n_566),
.B(n_581),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_625),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_591),
.B(n_554),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_617),
.B(n_586),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_609),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_598),
.B(n_574),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_603),
.B(n_628),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_607),
.B(n_616),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_626),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_626),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_616),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_589),
.B(n_586),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_632),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_605),
.B(n_586),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_596),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_608),
.B(n_557),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_599),
.A2(n_562),
.B1(n_543),
.B2(n_574),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_601),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_594),
.B(n_562),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_588),
.B(n_557),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_590),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_593),
.B(n_620),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_599),
.B(n_562),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_618),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_623),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_623),
.B(n_563),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_637),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_657),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_661),
.B(n_597),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_645),
.B(n_615),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_655),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_661),
.B(n_621),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_656),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_666),
.B(n_610),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_659),
.B(n_622),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_637),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_639),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_664),
.B(n_631),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_652),
.A2(n_663),
.B(n_647),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_639),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_655),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_657),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_653),
.B(n_630),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_666),
.B(n_638),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_642),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_659),
.B(n_606),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_640),
.B(n_606),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_642),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_650),
.B(n_556),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_638),
.B(n_563),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_644),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_636),
.B(n_650),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_636),
.B(n_615),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_653),
.B(n_662),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_SL g701 ( 
.A(n_649),
.B(n_600),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_651),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_644),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_640),
.B(n_575),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_673),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_690),
.B(n_680),
.Y(n_706)
);

NAND2x1p5_ASAP7_75t_L g707 ( 
.A(n_676),
.B(n_671),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_698),
.B(n_700),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_698),
.B(n_650),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_674),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_677),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_673),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_679),
.B(n_650),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_685),
.B(n_669),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_683),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_683),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_682),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_686),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_700),
.B(n_654),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_691),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_684),
.B(n_654),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_674),
.B(n_648),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_697),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_688),
.B(n_648),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_714),
.A2(n_701),
.B1(n_676),
.B2(n_669),
.Y(n_725)
);

NAND2x1_ASAP7_75t_L g726 ( 
.A(n_711),
.B(n_677),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_708),
.B(n_699),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_710),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_710),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_722),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_714),
.A2(n_701),
.B1(n_669),
.B2(n_689),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_707),
.A2(n_689),
.B1(n_692),
.B2(n_693),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_709),
.B(n_702),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_724),
.Y(n_734)
);

NOR2x1_ASAP7_75t_R g735 ( 
.A(n_719),
.B(n_668),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_L g736 ( 
.A1(n_725),
.A2(n_707),
.B1(n_706),
.B2(n_713),
.Y(n_736)
);

OAI21xp33_ASAP7_75t_SL g737 ( 
.A1(n_727),
.A2(n_722),
.B(n_724),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_728),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_726),
.Y(n_739)
);

AOI211xp5_ASAP7_75t_L g740 ( 
.A1(n_732),
.A2(n_678),
.B(n_675),
.C(n_681),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_731),
.A2(n_671),
.B1(n_704),
.B2(n_696),
.Y(n_741)
);

OAI21xp33_ASAP7_75t_SL g742 ( 
.A1(n_734),
.A2(n_721),
.B(n_723),
.Y(n_742)
);

AOI221xp5_ASAP7_75t_L g743 ( 
.A1(n_736),
.A2(n_732),
.B1(n_730),
.B2(n_729),
.C(n_733),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_737),
.B(n_735),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_740),
.B(n_720),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_741),
.A2(n_669),
.B1(n_695),
.B2(n_658),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_738),
.Y(n_747)
);

OAI31xp33_ASAP7_75t_L g748 ( 
.A1(n_739),
.A2(n_718),
.A3(n_717),
.B(n_716),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_744),
.B(n_742),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_747),
.Y(n_750)
);

XNOR2xp5_ASAP7_75t_L g751 ( 
.A(n_743),
.B(n_695),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_745),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_748),
.B(n_715),
.Y(n_753)
);

AO22x2_ASAP7_75t_L g754 ( 
.A1(n_752),
.A2(n_687),
.B1(n_712),
.B2(n_705),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_750),
.Y(n_755)
);

AOI221xp5_ASAP7_75t_L g756 ( 
.A1(n_749),
.A2(n_753),
.B1(n_751),
.B2(n_746),
.C(n_667),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_756),
.A2(n_755),
.B1(n_754),
.B2(n_695),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_756),
.A2(n_665),
.B(n_667),
.C(n_658),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_755),
.B(n_665),
.C(n_556),
.Y(n_759)
);

NOR2x1_ASAP7_75t_L g760 ( 
.A(n_757),
.B(n_646),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_759),
.A2(n_665),
.B1(n_703),
.B2(n_672),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_758),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_759),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_759),
.Y(n_764)
);

NOR2x1_ASAP7_75t_L g765 ( 
.A(n_757),
.B(n_646),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_762),
.A2(n_670),
.B1(n_665),
.B2(n_658),
.C(n_635),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_763),
.A2(n_670),
.B(n_694),
.Y(n_767)
);

XOR2x1_ASAP7_75t_L g768 ( 
.A(n_764),
.B(n_635),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_760),
.A2(n_658),
.B1(n_660),
.B2(n_672),
.Y(n_769)
);

OR3x2_ASAP7_75t_L g770 ( 
.A(n_765),
.B(n_613),
.C(n_633),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_761),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_768),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_771),
.Y(n_773)
);

NOR4xp25_ASAP7_75t_SL g774 ( 
.A(n_766),
.B(n_633),
.C(n_613),
.D(n_552),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_767),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_773),
.Y(n_776)
);

XOR2x1_ASAP7_75t_L g777 ( 
.A(n_772),
.B(n_770),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_775),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_776),
.A2(n_769),
.B1(n_774),
.B2(n_635),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_777),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_778),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_780),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_781),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_782),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_784),
.B(n_783),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_785),
.A2(n_779),
.B1(n_635),
.B2(n_660),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_786),
.B(n_694),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_787),
.A2(n_660),
.B1(n_641),
.B2(n_643),
.Y(n_788)
);


endmodule