module fake_jpeg_29841_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_2),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx4f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_20),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_9),
.Y(n_20)
);

INVxp33_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_7),
.A2(n_10),
.B1(n_6),
.B2(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

XOR2x2_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_20),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_32),
.B(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_19),
.B1(n_24),
.B2(n_27),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_35),
.B1(n_20),
.B2(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

AOI322xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_36),
.A3(n_37),
.B1(n_23),
.B2(n_18),
.C1(n_24),
.C2(n_31),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_23),
.B1(n_10),
.B2(n_11),
.Y(n_41)
);


endmodule