module real_jpeg_25559_n_17 (n_108, n_8, n_0, n_111, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_106, n_11, n_14, n_110, n_112, n_7, n_3, n_5, n_4, n_105, n_109, n_1, n_16, n_15, n_13, n_113, n_103, n_17);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_106;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_3;
input n_5;
input n_4;
input n_105;
input n_109;
input n_1;
input n_16;
input n_15;
input n_13;
input n_113;
input n_103;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_1),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_1),
.B(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_2),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_3),
.B(n_57),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_5),
.B(n_29),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_6),
.B(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_7),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_8),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_12),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_12),
.B(n_86),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g17 ( 
.A(n_14),
.B(n_18),
.CI(n_27),
.CON(n_17),
.SN(n_17)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_15),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_23),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_23),
.B(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_26),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_100),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_94),
.B(n_99),
.Y(n_31)
);

OAI321xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_85),
.A3(n_89),
.B1(n_92),
.B2(n_93),
.C(n_103),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_79),
.B(n_84),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_74),
.B(n_78),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_68),
.B(n_73),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_67),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_60),
.B(n_66),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_56),
.B(n_59),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B(n_55),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_62),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_70),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_98),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_104),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_105),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_106),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_107),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_108),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_109),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_110),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_111),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_112),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_113),
.Y(n_91)
);


endmodule