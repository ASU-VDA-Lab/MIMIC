module real_aes_7381_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_726;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_693;
wire n_496;
wire n_281;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_725;
wire n_455;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_817;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_749;
wire n_385;
wire n_275;
wire n_358;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_692;
wire n_789;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_753;
wire n_283;
wire n_314;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_0), .A2(n_246), .B1(n_648), .B2(n_649), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_1), .A2(n_257), .B1(n_623), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_2), .A2(n_248), .B1(n_480), .B2(n_765), .Y(n_764) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_3), .A2(n_42), .B1(n_287), .B2(n_303), .C(n_308), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_4), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_5), .B(n_347), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_6), .Y(n_576) );
AOI22xp5_ASAP7_75t_SL g740 ( .A1(n_7), .A2(n_70), .B1(n_513), .B2(n_741), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_8), .A2(n_23), .B1(n_454), .B2(n_496), .Y(n_677) );
AOI222xp33_ASAP7_75t_L g835 ( .A1(n_9), .A2(n_38), .B1(n_122), .B2(n_363), .C1(n_523), .C2(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_10), .A2(n_83), .B1(n_578), .B2(n_580), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_11), .A2(n_267), .B1(n_516), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_12), .A2(n_133), .B1(n_343), .B2(n_516), .Y(n_515) );
XOR2x2_ASAP7_75t_L g610 ( .A(n_13), .B(n_611), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_14), .A2(n_184), .B1(n_311), .B2(n_581), .Y(n_613) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_15), .A2(n_129), .B1(n_411), .B2(n_493), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_16), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_17), .A2(n_222), .B1(n_342), .B2(n_346), .C(n_348), .Y(n_341) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_18), .A2(n_143), .B1(n_471), .B2(n_472), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_19), .A2(n_148), .B1(n_366), .B2(n_637), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g694 ( .A1(n_20), .A2(n_117), .B1(n_139), .B2(n_440), .C1(n_541), .C2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_21), .A2(n_191), .B1(n_471), .B2(n_710), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_22), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_24), .Y(n_829) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_25), .A2(n_54), .B1(n_346), .B2(n_831), .C(n_832), .Y(n_830) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_26), .A2(n_230), .B1(n_327), .B2(n_578), .C(n_819), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_27), .A2(n_570), .B1(n_606), .B2(n_607), .Y(n_569) );
INVx1_ASAP7_75t_L g607 ( .A(n_27), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_28), .A2(n_179), .B1(n_507), .B2(n_508), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_29), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_30), .Y(n_403) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_31), .A2(n_96), .B1(n_292), .B2(n_297), .Y(n_300) );
INVx1_ASAP7_75t_L g790 ( .A(n_31), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_32), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_33), .A2(n_43), .B1(n_399), .B2(n_695), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_34), .A2(n_73), .B1(n_654), .B2(n_655), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_35), .Y(n_309) );
AOI22xp5_ASAP7_75t_SL g739 ( .A1(n_36), .A2(n_264), .B1(n_417), .B2(n_649), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g824 ( .A1(n_37), .A2(n_81), .B1(n_303), .B2(n_825), .C(n_827), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_39), .A2(n_164), .B1(n_495), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_40), .A2(n_89), .B1(n_504), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_41), .A2(n_195), .B1(n_337), .B2(n_452), .Y(n_554) );
AOI22xp5_ASAP7_75t_SL g734 ( .A1(n_44), .A2(n_149), .B1(n_409), .B2(n_735), .Y(n_734) );
AO22x1_ASAP7_75t_L g527 ( .A1(n_45), .A2(n_528), .B1(n_559), .B2(n_560), .Y(n_527) );
INVx1_ASAP7_75t_L g559 ( .A(n_45), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_46), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_47), .A2(n_65), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_48), .A2(n_261), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_49), .A2(n_225), .B1(n_449), .B2(n_557), .Y(n_556) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_50), .A2(n_135), .B1(n_199), .B2(n_439), .C1(n_440), .C2(n_541), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_51), .A2(n_255), .B1(n_420), .B2(n_493), .Y(n_809) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_52), .A2(n_99), .B1(n_292), .B2(n_293), .Y(n_302) );
INVx1_ASAP7_75t_L g791 ( .A(n_52), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_53), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_55), .A2(n_76), .B1(n_480), .B2(n_519), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_56), .A2(n_206), .B1(n_481), .B2(n_519), .Y(n_802) );
AOI222xp33_ASAP7_75t_L g521 ( .A1(n_57), .A2(n_163), .B1(n_218), .B2(n_401), .C1(n_522), .C2(n_523), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_58), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_59), .A2(n_167), .B1(n_454), .B2(n_474), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_60), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_61), .A2(n_269), .B1(n_327), .B2(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_62), .A2(n_91), .B1(n_643), .B2(n_644), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_63), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_64), .Y(n_443) );
XOR2xp5_ASAP7_75t_L g682 ( .A(n_66), .B(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_67), .A2(n_239), .B1(n_409), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_68), .A2(n_251), .B1(n_551), .B2(n_552), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_69), .A2(n_630), .B1(n_631), .B2(n_657), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_69), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_71), .A2(n_142), .B1(n_480), .B2(n_488), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_72), .A2(n_240), .B1(n_287), .B2(n_420), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_74), .A2(n_201), .B1(n_421), .B2(n_507), .Y(n_757) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_75), .A2(n_136), .B1(n_407), .B2(n_409), .Y(n_406) );
AOI222xp33_ASAP7_75t_L g362 ( .A1(n_77), .A2(n_102), .B1(n_158), .B2(n_363), .C1(n_366), .C2(n_372), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_78), .A2(n_124), .B1(n_411), .B2(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g625 ( .A(n_79), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_80), .A2(n_138), .B1(n_471), .B2(n_808), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_82), .A2(n_131), .B1(n_322), .B2(n_327), .C(n_331), .Y(n_321) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_84), .A2(n_247), .B1(n_623), .B2(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_85), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_86), .A2(n_165), .B1(n_305), .B2(n_472), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_87), .A2(n_252), .B1(n_374), .B2(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_88), .A2(n_97), .B1(n_346), .B2(n_484), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_90), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_92), .A2(n_216), .B1(n_578), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_93), .A2(n_154), .B1(n_651), .B2(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_94), .A2(n_214), .B1(n_481), .B2(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_95), .A2(n_134), .B1(n_327), .B2(n_619), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_98), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_100), .A2(n_817), .B1(n_837), .B2(n_838), .Y(n_816) );
INVx1_ASAP7_75t_L g837 ( .A(n_100), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_101), .B(n_342), .Y(n_730) );
INVx1_ASAP7_75t_L g278 ( .A(n_103), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_104), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_105), .A2(n_119), .B1(n_502), .B2(n_581), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_106), .A2(n_145), .B1(n_368), .B2(n_399), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_107), .A2(n_121), .B1(n_449), .B2(n_502), .Y(n_666) );
INVx1_ASAP7_75t_L g276 ( .A(n_108), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_109), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_110), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_111), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_112), .A2(n_130), .B1(n_502), .B2(n_508), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_113), .Y(n_828) );
OA22x2_ASAP7_75t_L g384 ( .A1(n_114), .A2(n_385), .B1(n_386), .B2(n_387), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_114), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_115), .A2(n_150), .B1(n_496), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_116), .A2(n_118), .B1(n_586), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_120), .A2(n_140), .B1(n_488), .B2(n_627), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_123), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_125), .A2(n_217), .B1(n_407), .B2(n_449), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_126), .A2(n_132), .B1(n_303), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g726 ( .A1(n_127), .A2(n_173), .B1(n_366), .B2(n_399), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_128), .A2(n_169), .B1(n_471), .B2(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_137), .Y(n_354) );
XNOR2x2_ASAP7_75t_L g498 ( .A(n_141), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g279 ( .A(n_144), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_146), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_147), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_151), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_152), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_153), .Y(n_834) );
INVx1_ASAP7_75t_L g715 ( .A(n_155), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_156), .B(n_401), .Y(n_400) );
XOR2xp5_ASAP7_75t_L g793 ( .A(n_157), .B(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_159), .A2(n_263), .B1(n_452), .B2(n_454), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_160), .B(n_484), .Y(n_483) );
AND2x6_ASAP7_75t_L g275 ( .A(n_161), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_161), .Y(n_784) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_162), .A2(n_231), .B1(n_292), .B2(n_293), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_166), .A2(n_249), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp5_ASAP7_75t_SL g736 ( .A1(n_168), .A2(n_229), .B1(n_414), .B2(n_737), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_170), .A2(n_238), .B1(n_327), .B2(n_417), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_171), .Y(n_799) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_172), .B(n_342), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_174), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_175), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_176), .B(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_177), .A2(n_223), .B1(n_449), .B2(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_178), .Y(n_833) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_180), .A2(n_186), .B1(n_420), .B2(n_421), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_181), .A2(n_268), .B1(n_346), .B2(n_484), .Y(n_621) );
AO22x2_ASAP7_75t_L g296 ( .A1(n_182), .A2(n_241), .B1(n_292), .B2(n_297), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_183), .A2(n_266), .B1(n_495), .B2(n_496), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_185), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_187), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_188), .A2(n_250), .B1(n_414), .B2(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_189), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_190), .A2(n_226), .B1(n_495), .B2(n_693), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_192), .A2(n_745), .B1(n_773), .B2(n_774), .Y(n_744) );
INVx1_ASAP7_75t_L g773 ( .A(n_192), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_193), .A2(n_211), .B1(n_372), .B2(n_522), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_194), .A2(n_219), .B1(n_512), .B2(n_513), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_196), .Y(n_600) );
AO22x1_ASAP7_75t_L g284 ( .A1(n_197), .A2(n_285), .B1(n_376), .B2(n_377), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_197), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_198), .Y(n_670) );
INVx1_ASAP7_75t_L g742 ( .A(n_200), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_202), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_203), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_204), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_205), .A2(n_258), .B1(n_496), .B2(n_651), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_207), .A2(n_265), .B1(n_492), .B2(n_493), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_208), .A2(n_210), .B1(n_420), .B2(n_513), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_209), .A2(n_271), .B(n_280), .C(n_792), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_212), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_213), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_215), .B(n_347), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_220), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_221), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_224), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_227), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_228), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_231), .B(n_789), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_232), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_233), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_234), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_235), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_236), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_237), .Y(n_820) );
INVx1_ASAP7_75t_L g787 ( .A(n_241), .Y(n_787) );
OA22x2_ASAP7_75t_L g423 ( .A1(n_242), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_242), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_243), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_244), .B(n_342), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_245), .Y(n_456) );
INVx1_ASAP7_75t_L g292 ( .A(n_253), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_253), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_254), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_256), .A2(n_260), .B1(n_421), .B2(n_496), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_259), .B(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_262), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_276), .Y(n_783) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_277), .A2(n_782), .B(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_563), .B1(n_777), .B2(n_778), .C(n_779), .Y(n_280) );
INVx1_ASAP7_75t_L g777 ( .A(n_281), .Y(n_777) );
AOI22xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_527), .B1(n_561), .B2(n_562), .Y(n_281) );
INVx1_ASAP7_75t_L g561 ( .A(n_282), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_378), .B2(n_526), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g377 ( .A(n_285), .Y(n_377) );
AND4x1_ASAP7_75t_L g285 ( .A(n_286), .B(n_321), .C(n_341), .D(n_362), .Y(n_285) );
BUFx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g408 ( .A(n_288), .Y(n_408) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_288), .Y(n_495) );
BUFx2_ASAP7_75t_SL g735 ( .A(n_288), .Y(n_735) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_298), .Y(n_288) );
AND2x4_ASAP7_75t_L g313 ( .A(n_289), .B(n_314), .Y(n_313) );
AND2x6_ASAP7_75t_L g324 ( .A(n_289), .B(n_325), .Y(n_324) );
AND2x6_ASAP7_75t_L g365 ( .A(n_289), .B(n_359), .Y(n_365) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_295), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_290), .B(n_296), .Y(n_307) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_291), .B(n_296), .Y(n_330) );
AND2x2_ASAP7_75t_L g352 ( .A(n_291), .B(n_300), .Y(n_352) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_294), .Y(n_297) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
INVx1_ASAP7_75t_L g371 ( .A(n_296), .Y(n_371) );
AND2x4_ASAP7_75t_L g306 ( .A(n_298), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_298), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g328 ( .A(n_298), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g418 ( .A(n_298), .B(n_319), .Y(n_418) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g314 ( .A(n_299), .B(n_302), .Y(n_314) );
OR2x2_ASAP7_75t_L g326 ( .A(n_299), .B(n_302), .Y(n_326) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g359 ( .A(n_300), .B(n_302), .Y(n_359) );
INVx1_ASAP7_75t_L g353 ( .A(n_301), .Y(n_353) );
AND2x2_ASAP7_75t_L g370 ( .A(n_301), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g340 ( .A(n_302), .Y(n_340) );
INVx4_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g648 ( .A(n_304), .Y(n_648) );
INVx4_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g409 ( .A(n_306), .Y(n_409) );
BUFx3_ASAP7_75t_L g474 ( .A(n_306), .Y(n_474) );
INVx2_ASAP7_75t_L g553 ( .A(n_306), .Y(n_553) );
BUFx3_ASAP7_75t_L g619 ( .A(n_306), .Y(n_619) );
AND2x4_ASAP7_75t_L g345 ( .A(n_307), .B(n_325), .Y(n_345) );
AND2x6_ASAP7_75t_L g347 ( .A(n_307), .B(n_314), .Y(n_347) );
INVx1_ASAP7_75t_L g393 ( .A(n_307), .Y(n_393) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_307), .B(n_314), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B1(n_315), .B2(n_316), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_310), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_455) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g513 ( .A(n_312), .Y(n_513) );
INVx2_ASAP7_75t_L g557 ( .A(n_312), .Y(n_557) );
INVx3_ASAP7_75t_L g676 ( .A(n_312), .Y(n_676) );
INVx6_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g421 ( .A(n_313), .Y(n_421) );
BUFx3_ASAP7_75t_L g493 ( .A(n_313), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_314), .B(n_319), .Y(n_334) );
AND2x2_ASAP7_75t_L g413 ( .A(n_314), .B(n_319), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g747 ( .A1(n_316), .A2(n_748), .B1(n_749), .B2(n_751), .C(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g458 ( .A(n_317), .Y(n_458) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g361 ( .A(n_320), .Y(n_361) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx4_ASAP7_75t_L g420 ( .A(n_323), .Y(n_420) );
INVx2_ASAP7_75t_SL g741 ( .A(n_323), .Y(n_741) );
INVx11_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx11_ASAP7_75t_L g450 ( .A(n_324), .Y(n_450) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g392 ( .A(n_326), .B(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g463 ( .A(n_328), .Y(n_463) );
BUFx3_ASAP7_75t_L g502 ( .A(n_328), .Y(n_502) );
BUFx2_ASAP7_75t_L g649 ( .A(n_328), .Y(n_649) );
BUFx3_ASAP7_75t_L g710 ( .A(n_328), .Y(n_710) );
BUFx2_ASAP7_75t_SL g750 ( .A(n_328), .Y(n_750) );
BUFx2_ASAP7_75t_SL g808 ( .A(n_328), .Y(n_808) );
AND2x2_ASAP7_75t_L g472 ( .A(n_329), .B(n_353), .Y(n_472) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x6_ASAP7_75t_L g339 ( .A(n_330), .B(n_340), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B1(n_335), .B2(n_336), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_333), .A2(n_820), .B1(n_821), .B2(n_822), .Y(n_819) );
BUFx2_ASAP7_75t_R g333 ( .A(n_334), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_337), .Y(n_336) );
BUFx4f_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g414 ( .A(n_338), .Y(n_414) );
BUFx2_ASAP7_75t_L g454 ( .A(n_338), .Y(n_454) );
BUFx2_ASAP7_75t_L g823 ( .A(n_338), .Y(n_823) );
INVx6_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g504 ( .A(n_339), .Y(n_504) );
INVx1_ASAP7_75t_SL g651 ( .A(n_339), .Y(n_651) );
INVx1_ASAP7_75t_L g489 ( .A(n_340), .Y(n_489) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx5_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g484 ( .A(n_344), .Y(n_484) );
INVx2_ASAP7_75t_L g704 ( .A(n_344), .Y(n_704) );
INVx2_ASAP7_75t_L g804 ( .A(n_344), .Y(n_804) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx4f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g517 ( .A(n_347), .Y(n_517) );
BUFx2_ASAP7_75t_L g640 ( .A(n_347), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_354), .B2(n_355), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_350), .A2(n_444), .B1(n_546), .B2(n_547), .Y(n_545) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_351), .A2(n_357), .B1(n_403), .B2(n_404), .Y(n_402) );
OAI22xp33_ASAP7_75t_SL g442 ( .A1(n_351), .A2(n_443), .B1(n_444), .B2(n_445), .Y(n_442) );
INVx4_ASAP7_75t_L g599 ( .A(n_351), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x4_ASAP7_75t_L g369 ( .A(n_352), .B(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g374 ( .A(n_352), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g488 ( .A(n_352), .B(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_355), .A2(n_598), .B1(n_833), .B2(n_834), .Y(n_832) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g444 ( .A(n_356), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g605 ( .A(n_357), .Y(n_605) );
OR2x6_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g481 ( .A(n_359), .B(n_361), .Y(n_481) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx4_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_364), .A2(n_477), .B(n_478), .Y(n_476) );
OAI21xp5_ASAP7_75t_SL g724 ( .A1(n_364), .A2(n_725), .B(n_726), .Y(n_724) );
INVx4_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx3_ASAP7_75t_L g401 ( .A(n_365), .Y(n_401) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_365), .Y(n_541) );
INVx2_ASAP7_75t_L g596 ( .A(n_365), .Y(n_596) );
INVx2_ASAP7_75t_L g798 ( .A(n_365), .Y(n_798) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx4_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g439 ( .A(n_368), .Y(n_439) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx4f_ASAP7_75t_SL g487 ( .A(n_369), .Y(n_487) );
BUFx2_ASAP7_75t_L g522 ( .A(n_369), .Y(n_522) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_369), .Y(n_627) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_369), .Y(n_689) );
INVx1_ASAP7_75t_L g375 ( .A(n_371), .Y(n_375) );
INVx2_ASAP7_75t_L g543 ( .A(n_372), .Y(n_543) );
BUFx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g771 ( .A(n_373), .Y(n_771) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx12f_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_374), .Y(n_479) );
INVx1_ASAP7_75t_L g526 ( .A(n_378), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_464), .B2(n_525), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_422), .B2(n_423), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND3x1_ASAP7_75t_L g387 ( .A(n_388), .B(n_405), .C(n_415), .Y(n_387) );
NOR3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_397), .C(n_402), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_394), .B2(n_395), .Y(n_389) );
BUFx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_392), .Y(n_431) );
INVx2_ASAP7_75t_L g533 ( .A(n_392), .Y(n_533) );
BUFx3_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_395), .A2(n_590), .B1(n_591), .B2(n_592), .Y(n_589) );
INVx2_ASAP7_75t_L g762 ( .A(n_395), .Y(n_762) );
BUFx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g536 ( .A(n_396), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx2_ASAP7_75t_L g441 ( .A(n_399), .Y(n_441) );
BUFx4f_ASAP7_75t_SL g523 ( .A(n_399), .Y(n_523) );
INVx3_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_410), .Y(n_405) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g668 ( .A(n_408), .Y(n_668) );
INVx1_ASAP7_75t_L g461 ( .A(n_409), .Y(n_461) );
INVx5_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx4_ASAP7_75t_L g453 ( .A(n_412), .Y(n_453) );
INVx3_ASAP7_75t_L g496 ( .A(n_412), .Y(n_496) );
BUFx3_ASAP7_75t_L g587 ( .A(n_412), .Y(n_587) );
INVx2_ASAP7_75t_L g615 ( .A(n_412), .Y(n_615) );
INVx8_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_419), .Y(n_415) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx3_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
BUFx3_ASAP7_75t_L g510 ( .A(n_418), .Y(n_510) );
BUFx3_ASAP7_75t_L g581 ( .A(n_418), .Y(n_581) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_446), .Y(n_426) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_435), .C(n_442), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g428 ( .A1(n_429), .A2(n_432), .B1(n_433), .B2(n_434), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI221xp5_ASAP7_75t_SL g759 ( .A1(n_431), .A2(n_760), .B1(n_761), .B2(n_763), .C(n_764), .Y(n_759) );
OAI21xp33_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_437), .B(n_438), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_436), .A2(n_625), .B(n_626), .Y(n_624) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_455), .C(n_459), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_SL g492 ( .A(n_450), .Y(n_492) );
INVx4_ASAP7_75t_L g512 ( .A(n_450), .Y(n_512) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_450), .Y(n_573) );
INVx5_ASAP7_75t_SL g693 ( .A(n_450), .Y(n_693) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g737 ( .A(n_453), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_458), .A2(n_575), .B1(n_828), .B2(n_829), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_462), .B2(n_463), .Y(n_459) );
OAI221xp5_ASAP7_75t_SL g582 ( .A1(n_463), .A2(n_553), .B1(n_583), .B2(n_584), .C(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g525 ( .A(n_464), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_498), .B2(n_524), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
XOR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_497), .Y(n_467) );
NAND3x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_475), .C(n_490), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
BUFx2_ASAP7_75t_L g812 ( .A(n_474), .Y(n_812) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_482), .Y(n_475) );
BUFx4f_ASAP7_75t_L g637 ( .A(n_479), .Y(n_637) );
INVx1_ASAP7_75t_SL g645 ( .A(n_480), .Y(n_645) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx3_ASAP7_75t_L g695 ( .A(n_481), .Y(n_695) );
BUFx2_ASAP7_75t_SL g732 ( .A(n_481), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .C(n_486), .Y(n_482) );
BUFx2_ASAP7_75t_L g831 ( .A(n_484), .Y(n_831) );
INVx1_ASAP7_75t_L g594 ( .A(n_487), .Y(n_594) );
INVx1_ASAP7_75t_L g520 ( .A(n_488), .Y(n_520) );
BUFx3_ASAP7_75t_L g623 ( .A(n_488), .Y(n_623) );
BUFx2_ASAP7_75t_L g765 ( .A(n_488), .Y(n_765) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_494), .Y(n_490) );
INVx1_ASAP7_75t_L g826 ( .A(n_492), .Y(n_826) );
INVx3_ASAP7_75t_L g575 ( .A(n_493), .Y(n_575) );
BUFx3_ASAP7_75t_L g507 ( .A(n_495), .Y(n_507) );
BUFx3_ASAP7_75t_L g551 ( .A(n_495), .Y(n_551) );
INVx3_ASAP7_75t_L g579 ( .A(n_495), .Y(n_579) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_495), .Y(n_654) );
INVx2_ASAP7_75t_L g524 ( .A(n_498), .Y(n_524) );
NAND4xp75_ASAP7_75t_L g499 ( .A(n_500), .B(n_505), .C(n_514), .D(n_521), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx4f_ASAP7_75t_SL g655 ( .A(n_510), .Y(n_655) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_515), .B(n_518), .Y(n_514) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_SL g729 ( .A(n_517), .Y(n_729) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g643 ( .A(n_520), .Y(n_643) );
INVx1_ASAP7_75t_L g538 ( .A(n_522), .Y(n_538) );
INVx1_ASAP7_75t_L g603 ( .A(n_523), .Y(n_603) );
INVx1_ASAP7_75t_L g562 ( .A(n_527), .Y(n_562) );
INVx1_ASAP7_75t_SL g560 ( .A(n_528), .Y(n_560) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_548), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_537), .C(n_545), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B1(n_534), .B2(n_535), .Y(n_530) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g591 ( .A(n_533), .Y(n_591) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g671 ( .A(n_536), .Y(n_671) );
OAI222xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_540), .B2(n_542), .C1(n_543), .C2(n_544), .Y(n_537) );
OAI222xp33_ASAP7_75t_L g766 ( .A1(n_540), .A2(n_767), .B1(n_768), .B2(n_769), .C1(n_770), .C2(n_772), .Y(n_766) );
INVx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g634 ( .A(n_541), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_555), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g778 ( .A(n_563), .Y(n_778) );
XNOR2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_719), .Y(n_563) );
OAI22xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_566), .B1(n_659), .B2(n_718), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_608), .B2(n_609), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g606 ( .A(n_570), .Y(n_606) );
AND2x2_ASAP7_75t_SL g570 ( .A(n_571), .B(n_588), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_582), .Y(n_571) );
OAI221xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_574), .B1(n_575), .B2(n_576), .C(n_577), .Y(n_572) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_593), .C(n_601), .Y(n_588) );
OAI222xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_596), .B2(n_597), .C1(n_598), .C2(n_600), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_596), .A2(n_700), .B(n_701), .Y(n_699) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AO22x1_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_628), .B1(n_629), .B2(n_658), .Y(n_609) );
INVx1_ASAP7_75t_SL g658 ( .A(n_610), .Y(n_658) );
NOR4xp75_ASAP7_75t_L g611 ( .A(n_612), .B(n_616), .C(n_620), .D(n_624), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_613), .B(n_614), .Y(n_612) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_615), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_617), .B(n_618), .Y(n_616) );
BUFx2_ASAP7_75t_L g756 ( .A(n_619), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_621), .B(n_622), .Y(n_620) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_627), .Y(n_836) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g657 ( .A(n_631), .Y(n_657) );
NAND3x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_646), .C(n_652), .Y(n_631) );
NOR2x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_638), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_635), .B(n_636), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .C(n_642), .Y(n_638) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_650), .Y(n_646) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g718 ( .A(n_659), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_680), .B2(n_681), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
XNOR2x2_ASAP7_75t_L g720 ( .A(n_663), .B(n_721), .Y(n_720) );
XOR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_679), .Y(n_663) );
NAND4xp75_ASAP7_75t_L g664 ( .A(n_665), .B(n_669), .C(n_674), .D(n_678), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
OA211x2_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B(n_672), .C(n_673), .Y(n_669) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
AO22x2_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_696), .B1(n_716), .B2(n_717), .Y(n_681) );
INVx1_ASAP7_75t_L g716 ( .A(n_682), .Y(n_716) );
NAND5xp2_ASAP7_75t_SL g683 ( .A(n_684), .B(n_685), .C(n_686), .D(n_690), .E(n_694), .Y(n_683) );
AND2x2_ASAP7_75t_SL g686 ( .A(n_687), .B(n_688), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_689), .Y(n_767) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx2_ASAP7_75t_L g717 ( .A(n_696), .Y(n_717) );
XOR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_715), .Y(n_696) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_698), .B(n_707), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .C(n_706), .Y(n_702) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
OAI22xp5_ASAP7_75t_SL g719 ( .A1(n_720), .A2(n_743), .B1(n_775), .B2(n_776), .Y(n_719) );
INVx1_ASAP7_75t_L g775 ( .A(n_720), .Y(n_775) );
XOR2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_742), .Y(n_721) );
NAND3x1_ASAP7_75t_L g722 ( .A(n_723), .B(n_733), .C(n_738), .Y(n_722) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .C(n_731), .Y(n_727) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx2_ASAP7_75t_L g776 ( .A(n_743), .Y(n_776) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g774 ( .A(n_745), .Y(n_774) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_746), .B(n_758), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_754), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
NOR2xp33_ASAP7_75t_SL g758 ( .A(n_759), .B(n_766), .Y(n_758) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVxp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
NOR2x1_ASAP7_75t_L g780 ( .A(n_781), .B(n_785), .Y(n_780) );
OR2x2_ASAP7_75t_SL g839 ( .A(n_781), .B(n_786), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_782), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_783), .B(n_815), .Y(n_842) );
CKINVDCx16_ASAP7_75t_R g815 ( .A(n_784), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_788), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
OAI222xp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_814), .B1(n_816), .B2(n_837), .C1(n_839), .C2(n_840), .Y(n_792) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_805), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_801), .Y(n_796) );
OAI21xp5_ASAP7_75t_SL g797 ( .A1(n_798), .A2(n_799), .B(n_800), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
NOR2x1_ASAP7_75t_L g805 ( .A(n_806), .B(n_810), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g838 ( .A(n_817), .Y(n_838) );
AND4x1_ASAP7_75t_L g817 ( .A(n_818), .B(n_824), .C(n_830), .D(n_835), .Y(n_817) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_841), .Y(n_840) );
endmodule