module fake_ibex_611_n_4999 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4999);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4999;

wire n_4557;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_962;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_3479;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_4569;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_2253;
wire n_4479;
wire n_3858;
wire n_4173;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_3060;
wire n_4124;
wire n_971;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_3293;
wire n_2550;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2625;
wire n_2444;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_4757;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4625;
wire n_4151;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_1471;
wire n_3441;
wire n_4559;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_1127;
wire n_947;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_2422;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_972;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_2223;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_977;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_1607;
wire n_2959;
wire n_2420;
wire n_2380;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1072;
wire n_2194;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_3096;
wire n_1278;
wire n_2059;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_950;
wire n_4282;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_985;
wire n_4611;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_4895;
wire n_3354;
wire n_4069;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_2574;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_1518;
wire n_4350;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_4686;
wire n_4682;
wire n_2914;
wire n_1833;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_4733;
wire n_987;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_1012;
wire n_960;
wire n_4412;
wire n_4266;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_3857;
wire n_2357;
wire n_4354;
wire n_2937;
wire n_3728;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_4539;
wire n_1205;
wire n_2969;
wire n_3550;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_2978;
wire n_3502;
wire n_3935;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_4926;
wire n_4688;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_969;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_3484;
wire n_2485;
wire n_4477;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_948;
wire n_3726;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4545;
wire n_2643;
wire n_4246;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_4491;
wire n_4672;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_4433;
wire n_3030;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4997;
wire n_4393;
wire n_3777;
wire n_4553;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_3633;
wire n_1731;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_2076;
wire n_974;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_959;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_965;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_2176;
wire n_2805;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_3787;
wire n_3445;
wire n_2080;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_4991;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_2142;
wire n_3703;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_954;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_998;
wire n_1729;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_4579;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_4636;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_2442;
wire n_1067;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_1662;
wire n_3443;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_1660;
wire n_4000;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_3712;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_976;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_3327;
wire n_1114;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_1885;
wire n_1989;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_1221;
wire n_3875;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_4565;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_956;
wire n_4597;
wire n_1812;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_4562;
wire n_1584;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_4196;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_2671;
wire n_3296;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_953;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_3036;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_3332;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_1442;
wire n_2168;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_3861;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_955;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_1640;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_4590;
wire n_4602;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2673;
wire n_2430;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_1743;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_4943;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_4159;
wire n_4372;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_3653;
wire n_4360;
wire n_4897;
wire n_963;
wire n_2139;
wire n_3693;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_3641;
wire n_4887;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_3722;
wire n_3802;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_4806;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_2859;
wire n_2564;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_2114;
wire n_1609;
wire n_3530;
wire n_1132;
wire n_4548;
wire n_1803;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_2660;
wire n_4604;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4126;
wire n_4103;
wire n_4710;
wire n_3282;
wire n_1003;
wire n_2708;
wire n_2748;
wire n_2224;
wire n_2233;
wire n_2499;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_1553;
wire n_3542;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_4504;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_2852;
wire n_2132;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_4747;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_2481;
wire n_4409;
wire n_1264;
wire n_2808;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_4152;
wire n_1352;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_4500;
wire n_1395;
wire n_1115;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_951;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_2414;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_3328;
wire n_2763;
wire n_994;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_961;
wire n_3735;
wire n_2127;
wire n_3228;
wire n_3028;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_2086;
wire n_4832;
wire n_3666;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2108;
wire n_2535;
wire n_2945;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_2894;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_975;
wire n_4900;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_2315;
wire n_3623;
wire n_2157;
wire n_3446;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_1105;
wire n_2898;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_4670;
wire n_4982;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_4053;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_1693;
wire n_2081;
wire n_2993;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_3989;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_967;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_3430;
wire n_1685;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_1398;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_4088;
wire n_2136;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4972;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_2262;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_983;
wire n_4224;
wire n_4868;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_4967;
wire n_1080;
wire n_2290;
wire n_957;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4668;
wire n_2383;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_2230;
wire n_3033;
wire n_2151;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_1606;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_979;
wire n_1999;
wire n_3810;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_2826;
wire n_2112;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_4671;
wire n_1326;
wire n_4981;
wire n_978;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_3618;
wire n_2727;
wire n_2719;
wire n_2213;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_3847;
wire n_2203;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_2646;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_4996;
wire n_4136;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1360;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_1452;
wire n_4953;
wire n_4570;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_2819;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_4407;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_3680;
wire n_3624;
wire n_4989;
wire n_2467;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1464;
wire n_1566;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_4929;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_1009;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_2525;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4958;
wire n_4297;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_964;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_3588;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1458;
wire n_1694;
wire n_2271;
wire n_2356;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_2642;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_4048;
wire n_4084;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_2849;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_4860;
wire n_4438;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_2665;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_993;
wire n_2581;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_3454;
wire n_4143;
wire n_4410;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_958;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_1433;
wire n_1907;
wire n_3994;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_4487;
wire n_1165;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_3042;
wire n_2561;
wire n_2491;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_3551;
wire n_4147;
wire n_3992;
wire n_4811;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_1419;
wire n_4738;
wire n_980;
wire n_1193;
wire n_3557;
wire n_2928;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_4086;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_966;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_1791;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_1164;
wire n_3749;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_4978;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_614),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_881),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_795),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_806),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_46),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_80),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_413),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_561),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_861),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_904),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_665),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_841),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_847),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_544),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_62),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_143),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_860),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_747),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_261),
.Y(n_965)
);

CKINVDCx16_ASAP7_75t_R g966 ( 
.A(n_94),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_642),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_731),
.Y(n_968)
);

BUFx10_ASAP7_75t_L g969 ( 
.A(n_883),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_923),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_694),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_903),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_941),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_311),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_482),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_306),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_195),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_125),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_778),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_136),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_944),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_302),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_711),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_629),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_27),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_139),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_627),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_933),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_27),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_776),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_117),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_629),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_798),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_552),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_783),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_765),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_397),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_831),
.Y(n_998)
);

INVxp67_ASAP7_75t_SL g999 ( 
.A(n_930),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_673),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_886),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_912),
.Y(n_1002)
);

INVx4_ASAP7_75t_R g1003 ( 
.A(n_230),
.Y(n_1003)
);

BUFx10_ASAP7_75t_L g1004 ( 
.A(n_879),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_935),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_748),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_795),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_614),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_353),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_914),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_465),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_360),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_99),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_47),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_842),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_842),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_851),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_524),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_884),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_410),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_151),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_834),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_42),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_426),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_579),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_79),
.Y(n_1026)
);

BUFx10_ASAP7_75t_L g1027 ( 
.A(n_461),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_292),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_762),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_826),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_124),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_744),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_843),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_89),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_404),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_372),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_201),
.Y(n_1037)
);

CKINVDCx14_ASAP7_75t_R g1038 ( 
.A(n_637),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_739),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_471),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_153),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_370),
.Y(n_1042)
);

BUFx10_ASAP7_75t_L g1043 ( 
.A(n_809),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_696),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_918),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_878),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_407),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_39),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_302),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_937),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_136),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_286),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_285),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_797),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_919),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_862),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_744),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_251),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_716),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_817),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_928),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_307),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_669),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_419),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_6),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_773),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_58),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_208),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_132),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_484),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_343),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_631),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_704),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_326),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_910),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_155),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_901),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_244),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_813),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_455),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_875),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_198),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_845),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_798),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_700),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_271),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_768),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_267),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_2),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_939),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_173),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_16),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_157),
.Y(n_1093)
);

INVx4_ASAP7_75t_R g1094 ( 
.A(n_903),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_657),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_907),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_718),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_14),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_822),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_147),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_454),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_381),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_610),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_881),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_834),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_410),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_829),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_342),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_243),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_206),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_934),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_492),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_733),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_104),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_902),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_439),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_169),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_246),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_235),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_882),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_874),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_852),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_802),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_394),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_877),
.Y(n_1125)
);

CKINVDCx16_ASAP7_75t_R g1126 ( 
.A(n_850),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_880),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_936),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_940),
.Y(n_1129)
);

BUFx10_ASAP7_75t_L g1130 ( 
.A(n_924),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_166),
.Y(n_1131)
);

BUFx10_ASAP7_75t_L g1132 ( 
.A(n_506),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_669),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_628),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_300),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_898),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_913),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_782),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_564),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_271),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_855),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_871),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_846),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_835),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_506),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_475),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_565),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_741),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_773),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_528),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_292),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_899),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_205),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_222),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_806),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_683),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_232),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_646),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_843),
.Y(n_1159)
);

BUFx5_ASAP7_75t_L g1160 ( 
.A(n_122),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_127),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_905),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_507),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_447),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_920),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_688),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_757),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_916),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_787),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_726),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_121),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_219),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_679),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_638),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_189),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_11),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_110),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_945),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_916),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_876),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_68),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_67),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_315),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_87),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_796),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_873),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_455),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_128),
.Y(n_1188)
);

BUFx10_ASAP7_75t_L g1189 ( 
.A(n_889),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_268),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_872),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_430),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_832),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_22),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_128),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_245),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_839),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_199),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_893),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_764),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_830),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_911),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_156),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_548),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_330),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_94),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_730),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_6),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_465),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_813),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_921),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_356),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_758),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_556),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_902),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_440),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_941),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_474),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_477),
.Y(n_1219)
);

CKINVDCx16_ASAP7_75t_R g1220 ( 
.A(n_705),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_501),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_942),
.Y(n_1222)
);

INVxp33_ASAP7_75t_R g1223 ( 
.A(n_100),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_871),
.Y(n_1224)
);

INVxp33_ASAP7_75t_SL g1225 ( 
.A(n_667),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_301),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_760),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_468),
.Y(n_1228)
);

BUFx10_ASAP7_75t_L g1229 ( 
.A(n_675),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_839),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_200),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_327),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_619),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_883),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_866),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_32),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_180),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_926),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_560),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_240),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_301),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_743),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_777),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_789),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_841),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_778),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_417),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_833),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_909),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_848),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_209),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_573),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_521),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_224),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_852),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_43),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_837),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_788),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_206),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_169),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_131),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_268),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_9),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_700),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_888),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_9),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_20),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_857),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_801),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_549),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_895),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_709),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_864),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_186),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_865),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_931),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_571),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_104),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_911),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_781),
.Y(n_1280)
);

BUFx10_ASAP7_75t_L g1281 ( 
.A(n_713),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_869),
.Y(n_1282)
);

CKINVDCx14_ASAP7_75t_R g1283 ( 
.A(n_362),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_402),
.Y(n_1284)
);

BUFx5_ASAP7_75t_L g1285 ( 
.A(n_559),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_929),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_890),
.Y(n_1287)
);

BUFx8_ASAP7_75t_SL g1288 ( 
.A(n_294),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_330),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_28),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_372),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_809),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_686),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_246),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_933),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_859),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_638),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_943),
.Y(n_1298)
);

BUFx8_ASAP7_75t_SL g1299 ( 
.A(n_747),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_811),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_858),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_14),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_892),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_908),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_894),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_514),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_407),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_853),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_401),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_849),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_723),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_523),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_80),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_358),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_923),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_763),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_296),
.Y(n_1317)
);

CKINVDCx14_ASAP7_75t_R g1318 ( 
.A(n_63),
.Y(n_1318)
);

BUFx5_ASAP7_75t_L g1319 ( 
.A(n_820),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_590),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_917),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_502),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_891),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_856),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_374),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_863),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_60),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_136),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_304),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_844),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_867),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_466),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_646),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_536),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_600),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_79),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_91),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_550),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_210),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_438),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_385),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_650),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_854),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_818),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_370),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_938),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_237),
.Y(n_1347)
);

BUFx8_ASAP7_75t_SL g1348 ( 
.A(n_368),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_184),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_69),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_312),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_439),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_801),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_363),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_545),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_836),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_909),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_128),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_885),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_887),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_43),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_706),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_334),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_563),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_742),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_372),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_896),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_200),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_550),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_467),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_253),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_507),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_828),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_814),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_51),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_55),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_525),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_371),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_925),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_224),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_732),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_932),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_394),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_312),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_125),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_106),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_91),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_808),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_935),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_23),
.Y(n_1390)
);

BUFx5_ASAP7_75t_L g1391 ( 
.A(n_838),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_651),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_39),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_906),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_217),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_223),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_33),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_50),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_922),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_870),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_725),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_391),
.Y(n_1402)
);

BUFx5_ASAP7_75t_L g1403 ( 
.A(n_271),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_690),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_927),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_900),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_922),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_257),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_868),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_442),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_514),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_807),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_915),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_115),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_210),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_792),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_840),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_796),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_262),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_185),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_707),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_125),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_585),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_946),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_768),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_837),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_368),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_759),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_94),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_508),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_819),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_442),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_146),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_566),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_724),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_351),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_897),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_85),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1283),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1023),
.Y(n_1440)
);

CKINVDCx16_ASAP7_75t_R g1441 ( 
.A(n_966),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1109),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1283),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1174),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1216),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1038),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1259),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1319),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1318),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1272),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_1009),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1151),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1247),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1288),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1072),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1386),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_992),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1348),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1371),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1319),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_989),
.Y(n_1461)
);

INVxp67_ASAP7_75t_SL g1462 ( 
.A(n_989),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1240),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1297),
.Y(n_1464)
);

INVxp33_ASAP7_75t_SL g1465 ( 
.A(n_1142),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_952),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1319),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1319),
.Y(n_1468)
);

INVxp33_ASAP7_75t_SL g1469 ( 
.A(n_1217),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_954),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_957),
.Y(n_1471)
);

INVxp33_ASAP7_75t_SL g1472 ( 
.A(n_1346),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_967),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_1073),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1073),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_975),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_976),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_980),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_990),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_982),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_1078),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_990),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_983),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_997),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1027),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1000),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1008),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1011),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1107),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1018),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1021),
.Y(n_1491)
);

INVxp33_ASAP7_75t_L g1492 ( 
.A(n_1099),
.Y(n_1492)
);

INVxp33_ASAP7_75t_L g1493 ( 
.A(n_1121),
.Y(n_1493)
);

INVxp67_ASAP7_75t_SL g1494 ( 
.A(n_1086),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1299),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1025),
.Y(n_1496)
);

INVxp33_ASAP7_75t_SL g1497 ( 
.A(n_947),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1133),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1026),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1028),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1031),
.Y(n_1501)
);

CKINVDCx14_ASAP7_75t_R g1502 ( 
.A(n_1027),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1035),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1041),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1086),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1051),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1067),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1202),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1074),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1080),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1088),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1103),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1108),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_990),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1225),
.B(n_0),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1117),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1150),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1154),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1175),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1176),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1177),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1181),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1184),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1188),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1194),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1204),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1212),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1226),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1062),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1231),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1233),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1319),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1239),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1220),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1252),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_951),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1254),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1260),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1118),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1263),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1266),
.Y(n_1541)
);

CKINVDCx16_ASAP7_75t_R g1542 ( 
.A(n_998),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1132),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1270),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1284),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1118),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1290),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1203),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1291),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1293),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1294),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1215),
.Y(n_1552)
);

CKINVDCx16_ASAP7_75t_R g1553 ( 
.A(n_1126),
.Y(n_1553)
);

INVxp33_ASAP7_75t_SL g1554 ( 
.A(n_961),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1322),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1508),
.B(n_1273),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1440),
.B(n_1424),
.Y(n_1557)
);

BUFx12f_ASAP7_75t_L g1558 ( 
.A(n_1454),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1442),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1448),
.A2(n_1467),
.B(n_1460),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1468),
.Y(n_1561)
);

XNOR2x2_ASAP7_75t_L g1562 ( 
.A(n_1515),
.B(n_953),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1457),
.B(n_1132),
.Y(n_1563)
);

NOR2x1_ASAP7_75t_L g1564 ( 
.A(n_1463),
.B(n_1201),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1455),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1444),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1532),
.A2(n_1059),
.B(n_960),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1461),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1459),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1479),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1462),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1445),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1447),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1502),
.B(n_1229),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1474),
.B(n_962),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1555),
.A2(n_1059),
.B(n_960),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1475),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1481),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1479),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1450),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1485),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1494),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1485),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1466),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1536),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1470),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1471),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1505),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1473),
.A2(n_1095),
.B(n_1091),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1479),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1482),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1464),
.B(n_1229),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1511),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1497),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1539),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1452),
.B(n_948),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_L g1597 ( 
.A(n_1482),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1482),
.Y(n_1598)
);

AND2x6_ASAP7_75t_L g1599 ( 
.A(n_1543),
.B(n_1203),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1476),
.Y(n_1600)
);

INVx5_ASAP7_75t_L g1601 ( 
.A(n_1514),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1546),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1548),
.B(n_965),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1477),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1478),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1480),
.Y(n_1606)
);

CKINVDCx16_ASAP7_75t_R g1607 ( 
.A(n_1441),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1483),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1498),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1514),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1439),
.B(n_971),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1484),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1486),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1487),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1492),
.B(n_1281),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1488),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1451),
.A2(n_977),
.B1(n_978),
.B2(n_974),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1490),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1554),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1491),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1552),
.B(n_1496),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1499),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1453),
.B(n_1255),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1500),
.B(n_984),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1501),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1458),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1503),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1504),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1506),
.A2(n_1095),
.B(n_1091),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1507),
.A2(n_1119),
.B(n_1100),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1469),
.A2(n_991),
.B1(n_994),
.B2(n_987),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1509),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1510),
.A2(n_1119),
.B(n_1100),
.Y(n_1633)
);

CKINVDCx16_ASAP7_75t_R g1634 ( 
.A(n_1542),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1534),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1449),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1514),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1493),
.B(n_1277),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1456),
.B(n_1311),
.Y(n_1639)
);

NOR2x1_ASAP7_75t_L g1640 ( 
.A(n_1512),
.B(n_1201),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1513),
.B(n_1012),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1516),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1517),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1518),
.B(n_1013),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1519),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1520),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1521),
.B(n_1014),
.Y(n_1647)
);

BUFx12f_ASAP7_75t_L g1648 ( 
.A(n_1495),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1522),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1523),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1524),
.B(n_1525),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1526),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1527),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1528),
.Y(n_1654)
);

OA21x2_ASAP7_75t_L g1655 ( 
.A1(n_1530),
.A2(n_1140),
.B(n_1124),
.Y(n_1655)
);

NOR2x1_ASAP7_75t_L g1656 ( 
.A(n_1531),
.B(n_1277),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1443),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1533),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1446),
.B(n_1416),
.Y(n_1659)
);

BUFx8_ASAP7_75t_L g1660 ( 
.A(n_1553),
.Y(n_1660)
);

AND2x6_ASAP7_75t_L g1661 ( 
.A(n_1535),
.B(n_985),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1537),
.Y(n_1662)
);

INVx6_ASAP7_75t_L g1663 ( 
.A(n_1472),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1538),
.B(n_1160),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1540),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1541),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1529),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1544),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1545),
.B(n_1160),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1547),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1549),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1550),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1551),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1439),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1489),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1448),
.A2(n_1173),
.B(n_1164),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1479),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1455),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1489),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_L g1680 ( 
.A(n_1439),
.B(n_1160),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1489),
.Y(n_1681)
);

OA21x2_ASAP7_75t_L g1682 ( 
.A1(n_1448),
.A2(n_1173),
.B(n_1164),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1455),
.B(n_1020),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1489),
.Y(n_1684)
);

AND2x6_ASAP7_75t_L g1685 ( 
.A(n_1485),
.B(n_985),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1485),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1448),
.A2(n_1221),
.B(n_1183),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1502),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1489),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1440),
.B(n_1344),
.Y(n_1690)
);

BUFx12f_ASAP7_75t_L g1691 ( 
.A(n_1454),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1455),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1489),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1455),
.B(n_1024),
.Y(n_1694)
);

INVx5_ASAP7_75t_L g1695 ( 
.A(n_1479),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1489),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1489),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1489),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1489),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1502),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1439),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_SL g1702 ( 
.A(n_1485),
.B(n_1431),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1489),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1489),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1479),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1455),
.Y(n_1706)
);

INVx4_ASAP7_75t_L g1707 ( 
.A(n_1439),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1489),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1485),
.Y(n_1709)
);

AND2x2_ASAP7_75t_SL g1710 ( 
.A(n_1441),
.B(n_958),
.Y(n_1710)
);

INVx5_ASAP7_75t_L g1711 ( 
.A(n_1479),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1508),
.B(n_958),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1508),
.B(n_959),
.Y(n_1713)
);

OA21x2_ASAP7_75t_L g1714 ( 
.A1(n_1448),
.A2(n_1221),
.B(n_1183),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1465),
.A2(n_1036),
.B1(n_1037),
.B2(n_1034),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1489),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1502),
.Y(n_1717)
);

OAI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1448),
.A2(n_1307),
.B(n_1278),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1455),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1489),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1455),
.B(n_1040),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1508),
.B(n_959),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1457),
.B(n_1285),
.Y(n_1723)
);

INVx4_ASAP7_75t_L g1724 ( 
.A(n_1439),
.Y(n_1724)
);

CKINVDCx8_ASAP7_75t_R g1725 ( 
.A(n_1441),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1502),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1489),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1455),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1489),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1457),
.B(n_1285),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1485),
.B(n_1285),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1455),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1489),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1455),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1455),
.B(n_1044),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1455),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1489),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1479),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1489),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1479),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1489),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1463),
.B(n_1327),
.Y(n_1742)
);

BUFx10_ASAP7_75t_L g1743 ( 
.A(n_1700),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1660),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1573),
.Y(n_1745)
);

CKINVDCx20_ASAP7_75t_R g1746 ( 
.A(n_1607),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1667),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1688),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1717),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1580),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1726),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1559),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1626),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1725),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1634),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1558),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1691),
.Y(n_1757)
);

CKINVDCx20_ASAP7_75t_R g1758 ( 
.A(n_1583),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1566),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1648),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1572),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1565),
.B(n_1047),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1635),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1594),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1619),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1581),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1563),
.B(n_969),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1663),
.Y(n_1768)
);

NOR2xp67_ASAP7_75t_L g1769 ( 
.A(n_1609),
.B(n_0),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1718),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1600),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1629),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1574),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1604),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1653),
.B(n_1285),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1686),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1642),
.Y(n_1777)
);

INVxp67_ASAP7_75t_L g1778 ( 
.A(n_1709),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1657),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1629),
.Y(n_1780)
);

CKINVDCx20_ASAP7_75t_R g1781 ( 
.A(n_1585),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1727),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_R g1783 ( 
.A(n_1702),
.B(n_1045),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1574),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1617),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1654),
.B(n_1285),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1615),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1638),
.Y(n_1788)
);

CKINVDCx20_ASAP7_75t_R g1789 ( 
.A(n_1636),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1615),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_SL g1791 ( 
.A(n_1659),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1563),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1631),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1592),
.B(n_999),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1646),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1715),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1710),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_R g1798 ( 
.A(n_1674),
.B(n_1081),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1701),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_1592),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1666),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1670),
.B(n_1403),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1638),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1707),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1724),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1671),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1576),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1651),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1599),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1599),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1599),
.Y(n_1811)
);

OA21x2_ASAP7_75t_L g1812 ( 
.A1(n_1560),
.A2(n_1329),
.B(n_1328),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_R g1813 ( 
.A(n_1680),
.B(n_1104),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1556),
.B(n_969),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1569),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1562),
.Y(n_1816)
);

HB1xp67_ASAP7_75t_L g1817 ( 
.A(n_1683),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1733),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_R g1819 ( 
.A(n_1685),
.B(n_1168),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1664),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1739),
.Y(n_1821)
);

CKINVDCx20_ASAP7_75t_R g1822 ( 
.A(n_1621),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1611),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1664),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1694),
.Y(n_1825)
);

INVx8_ASAP7_75t_L g1826 ( 
.A(n_1685),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1669),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1649),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1721),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1735),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_R g1831 ( 
.A(n_1685),
.B(n_1200),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1655),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_R g1833 ( 
.A(n_1684),
.B(n_1234),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1589),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_R g1835 ( 
.A(n_1698),
.B(n_1246),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_1575),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1630),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1633),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1649),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_1603),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1723),
.Y(n_1841)
);

CKINVDCx16_ASAP7_75t_R g1842 ( 
.A(n_1730),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1730),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1655),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1652),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_R g1846 ( 
.A(n_1708),
.B(n_1258),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1624),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1712),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1652),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1658),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1720),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1567),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1713),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1722),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1678),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1692),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1567),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1658),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1706),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1568),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1571),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1719),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1728),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1732),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1734),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1577),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1736),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1676),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1578),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1676),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1596),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1582),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1588),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1675),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1593),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1595),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1623),
.B(n_1131),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1641),
.B(n_1004),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1682),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1602),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1639),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1557),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1644),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1647),
.Y(n_1884)
);

BUFx10_ASAP7_75t_L g1885 ( 
.A(n_1690),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1656),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1731),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1605),
.B(n_1606),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1687),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1584),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1679),
.Y(n_1891)
);

CKINVDCx6p67_ASAP7_75t_R g1892 ( 
.A(n_1661),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1586),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1587),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1608),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_R g1896 ( 
.A(n_1613),
.B(n_1296),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1687),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1681),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1714),
.Y(n_1899)
);

NOR2xp67_ASAP7_75t_L g1900 ( 
.A(n_1689),
.B(n_1),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1742),
.A2(n_1298),
.B1(n_1357),
.B2(n_1300),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1693),
.Y(n_1902)
);

NAND2xp33_ASAP7_75t_R g1903 ( 
.A(n_1714),
.B(n_1048),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1696),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1661),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1697),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1699),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1703),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1704),
.Y(n_1909)
);

BUFx2_ASAP7_75t_L g1910 ( 
.A(n_1612),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1614),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1616),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1716),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1618),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1729),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1737),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1620),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1741),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1622),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1625),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1628),
.Y(n_1921)
);

NAND2xp33_ASAP7_75t_R g1922 ( 
.A(n_1627),
.B(n_1049),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1632),
.B(n_1052),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1643),
.Y(n_1924)
);

INVxp33_ASAP7_75t_L g1925 ( 
.A(n_1564),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1645),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1650),
.Y(n_1927)
);

INVx2_ASAP7_75t_SL g1928 ( 
.A(n_1640),
.Y(n_1928)
);

CKINVDCx20_ASAP7_75t_R g1929 ( 
.A(n_1662),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1665),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1668),
.Y(n_1931)
);

AND2x6_ASAP7_75t_L g1932 ( 
.A(n_1672),
.B(n_1362),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1673),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1561),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1661),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1601),
.B(n_1004),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_R g1937 ( 
.A(n_1601),
.B(n_1407),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1695),
.Y(n_1938)
);

BUFx6f_ASAP7_75t_L g1939 ( 
.A(n_1570),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1695),
.Y(n_1940)
);

NAND2xp33_ASAP7_75t_R g1941 ( 
.A(n_1711),
.B(n_1053),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1711),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1570),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1579),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1740),
.B(n_1043),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1579),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1590),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1590),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1591),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1591),
.Y(n_1950)
);

AND2x6_ASAP7_75t_L g1951 ( 
.A(n_1597),
.B(n_1362),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1598),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1598),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1610),
.Y(n_1954)
);

CKINVDCx20_ASAP7_75t_R g1955 ( 
.A(n_1610),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1637),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1740),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1677),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1677),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1705),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1705),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1738),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_1738),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1660),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1660),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1629),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1718),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1573),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1660),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1660),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1660),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1660),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1638),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1660),
.Y(n_1974)
);

CKINVDCx20_ASAP7_75t_R g1975 ( 
.A(n_1607),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1573),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1573),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1660),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1629),
.Y(n_1979)
);

CKINVDCx20_ASAP7_75t_R g1980 ( 
.A(n_1607),
.Y(n_1980)
);

CKINVDCx20_ASAP7_75t_R g1981 ( 
.A(n_1607),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1583),
.B(n_1043),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1718),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1573),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1573),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1573),
.Y(n_1986)
);

AND2x6_ASAP7_75t_L g1987 ( 
.A(n_1820),
.B(n_985),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1955),
.Y(n_1988)
);

INVx2_ASAP7_75t_SL g1989 ( 
.A(n_1743),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1911),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1860),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1772),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1861),
.Y(n_1993)
);

AO22x2_ASAP7_75t_L g1994 ( 
.A1(n_1816),
.A2(n_1223),
.B1(n_1195),
.B2(n_1198),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1866),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1832),
.Y(n_1996)
);

BUFx10_ASAP7_75t_L g1997 ( 
.A(n_1744),
.Y(n_1997)
);

CKINVDCx6p67_ASAP7_75t_R g1998 ( 
.A(n_1791),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1832),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1788),
.B(n_1058),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1817),
.B(n_1063),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1765),
.B(n_1163),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1844),
.Y(n_2003)
);

AND2x2_ASAP7_75t_SL g2004 ( 
.A(n_1842),
.B(n_1003),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1803),
.B(n_1064),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1875),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1743),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1758),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1876),
.Y(n_2009)
);

AND2x2_ASAP7_75t_SL g2010 ( 
.A(n_1783),
.B(n_1787),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1826),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1880),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1825),
.B(n_1065),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1872),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1873),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1808),
.A2(n_1403),
.B1(n_1069),
.B2(n_1071),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1847),
.B(n_1068),
.Y(n_2017)
);

INVx4_ASAP7_75t_L g2018 ( 
.A(n_1964),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1829),
.B(n_1830),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1883),
.B(n_1884),
.Y(n_2020)
);

INVx4_ASAP7_75t_SL g2021 ( 
.A(n_1932),
.Y(n_2021)
);

NAND2x1_ASAP7_75t_L g2022 ( 
.A(n_1932),
.B(n_1094),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1965),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1888),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1844),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1789),
.B(n_1017),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1933),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1745),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1822),
.A2(n_1082),
.B1(n_1085),
.B2(n_1076),
.Y(n_2029)
);

OR2x6_ASAP7_75t_L g2030 ( 
.A(n_1766),
.B(n_1055),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1969),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1970),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1826),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1971),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1750),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1919),
.B(n_1920),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_SL g2037 ( 
.A1(n_1896),
.A2(n_1189),
.B1(n_1213),
.B2(n_1130),
.Y(n_2037)
);

INVx6_ASAP7_75t_L g2038 ( 
.A(n_1782),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1968),
.Y(n_2039)
);

INVx3_ASAP7_75t_L g2040 ( 
.A(n_1972),
.Y(n_2040)
);

INVx2_ASAP7_75t_SL g2041 ( 
.A(n_1776),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1976),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1930),
.B(n_1089),
.Y(n_2043)
);

INVx8_ASAP7_75t_L g2044 ( 
.A(n_1791),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1855),
.A2(n_1093),
.B1(n_1101),
.B2(n_1092),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1966),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1977),
.Y(n_2047)
);

INVx4_ASAP7_75t_L g2048 ( 
.A(n_1974),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1767),
.B(n_1102),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1978),
.Y(n_2050)
);

INVxp67_ASAP7_75t_SL g2051 ( 
.A(n_1895),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1780),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1984),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1921),
.B(n_1106),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1985),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_1882),
.B(n_1110),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1881),
.B(n_1790),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1986),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1792),
.B(n_1112),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1877),
.B(n_1261),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_1768),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1778),
.B(n_1116),
.Y(n_2062)
);

INVx4_ASAP7_75t_L g2063 ( 
.A(n_1799),
.Y(n_2063)
);

INVx4_ASAP7_75t_SL g2064 ( 
.A(n_1932),
.Y(n_2064)
);

BUFx6f_ASAP7_75t_L g2065 ( 
.A(n_1826),
.Y(n_2065)
);

BUFx2_ASAP7_75t_L g2066 ( 
.A(n_1781),
.Y(n_2066)
);

INVx4_ASAP7_75t_L g2067 ( 
.A(n_1804),
.Y(n_2067)
);

BUFx6f_ASAP7_75t_L g2068 ( 
.A(n_1780),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1979),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1890),
.Y(n_2070)
);

INVx3_ASAP7_75t_L g2071 ( 
.A(n_1805),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1979),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1893),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1979),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1807),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1834),
.Y(n_2076)
);

CKINVDCx20_ASAP7_75t_R g2077 ( 
.A(n_1746),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_1794),
.A2(n_1403),
.B1(n_1139),
.B2(n_1145),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1894),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1856),
.A2(n_1146),
.B1(n_1147),
.B2(n_1134),
.Y(n_2080)
);

INVx4_ASAP7_75t_L g2081 ( 
.A(n_1764),
.Y(n_2081)
);

BUFx3_ASAP7_75t_L g2082 ( 
.A(n_1975),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1912),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1837),
.Y(n_2084)
);

BUFx3_ASAP7_75t_L g2085 ( 
.A(n_1980),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1931),
.B(n_1153),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1982),
.B(n_1156),
.Y(n_2087)
);

OAI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1800),
.A2(n_1158),
.B1(n_1161),
.B2(n_1157),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1905),
.Y(n_2089)
);

INVx1_ASAP7_75t_SL g2090 ( 
.A(n_1917),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1838),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1871),
.B(n_1929),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1926),
.B(n_1927),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1914),
.Y(n_2094)
);

INVx4_ASAP7_75t_L g2095 ( 
.A(n_1756),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_1981),
.B(n_1358),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_1763),
.B(n_1363),
.Y(n_2097)
);

BUFx3_ASAP7_75t_L g2098 ( 
.A(n_1757),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1924),
.Y(n_2099)
);

INVx8_ASAP7_75t_L g2100 ( 
.A(n_1932),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1923),
.B(n_1762),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1798),
.Y(n_2102)
);

AND2x6_ASAP7_75t_L g2103 ( 
.A(n_1824),
.B(n_1827),
.Y(n_2103)
);

BUFx10_ASAP7_75t_L g2104 ( 
.A(n_1760),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1833),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1859),
.B(n_1166),
.Y(n_2106)
);

INVx6_ASAP7_75t_L g2107 ( 
.A(n_1945),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1862),
.B(n_1171),
.Y(n_2108)
);

INVx1_ASAP7_75t_SL g2109 ( 
.A(n_1835),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_1878),
.B(n_963),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1863),
.B(n_1172),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1815),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_1814),
.B(n_1754),
.Y(n_2113)
);

INVx1_ASAP7_75t_SL g2114 ( 
.A(n_1846),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1864),
.B(n_1182),
.Y(n_2115)
);

INVx8_ASAP7_75t_L g2116 ( 
.A(n_1818),
.Y(n_2116)
);

NAND2xp33_ASAP7_75t_SL g2117 ( 
.A(n_1819),
.B(n_1187),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1865),
.B(n_1190),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1852),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1857),
.Y(n_2120)
);

BUFx6f_ASAP7_75t_L g2121 ( 
.A(n_1905),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_1905),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1867),
.B(n_1192),
.Y(n_2123)
);

BUFx4f_ASAP7_75t_L g2124 ( 
.A(n_1851),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1802),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1771),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_1821),
.Y(n_2127)
);

INVx4_ASAP7_75t_L g2128 ( 
.A(n_1940),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_1869),
.B(n_1196),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_1748),
.B(n_970),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1809),
.B(n_1205),
.Y(n_2131)
);

BUFx10_ASAP7_75t_L g2132 ( 
.A(n_1755),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1868),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1774),
.B(n_1206),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_1874),
.Y(n_2135)
);

INVx3_ASAP7_75t_L g2136 ( 
.A(n_1915),
.Y(n_2136)
);

AND2x6_ASAP7_75t_L g2137 ( 
.A(n_1870),
.B(n_985),
.Y(n_2137)
);

INVx3_ASAP7_75t_SL g2138 ( 
.A(n_1753),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1951),
.Y(n_2139)
);

BUFx2_ASAP7_75t_L g2140 ( 
.A(n_1937),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1777),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1795),
.B(n_1208),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1801),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1806),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1879),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1752),
.Y(n_2146)
);

INVx4_ASAP7_75t_L g2147 ( 
.A(n_1749),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1759),
.Y(n_2148)
);

INVx4_ASAP7_75t_L g2149 ( 
.A(n_1751),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1889),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1761),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1841),
.B(n_1214),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1843),
.B(n_1218),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1810),
.B(n_1219),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_1747),
.B(n_1779),
.Y(n_2155)
);

OR2x6_ASAP7_75t_L g2156 ( 
.A(n_1901),
.B(n_1055),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1934),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1775),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1786),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_1938),
.Y(n_2160)
);

INVx4_ASAP7_75t_L g2161 ( 
.A(n_1784),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1886),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1897),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1900),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1936),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1928),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_1951),
.Y(n_2167)
);

AND2x6_ASAP7_75t_L g2168 ( 
.A(n_1899),
.B(n_986),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1769),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1836),
.B(n_1232),
.Y(n_2170)
);

BUFx3_ASAP7_75t_L g2171 ( 
.A(n_1946),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1770),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1811),
.B(n_1236),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1891),
.Y(n_2174)
);

OAI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_1840),
.A2(n_1241),
.B1(n_1251),
.B2(n_1237),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_1831),
.B(n_1253),
.Y(n_2176)
);

NAND2x1p5_ASAP7_75t_L g2177 ( 
.A(n_1942),
.B(n_1337),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1898),
.Y(n_2178)
);

AO22x2_ASAP7_75t_L g2179 ( 
.A1(n_1903),
.A2(n_973),
.B1(n_979),
.B2(n_972),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_1887),
.B(n_1256),
.Y(n_2180)
);

BUFx6f_ASAP7_75t_L g2181 ( 
.A(n_1951),
.Y(n_2181)
);

INVxp67_ASAP7_75t_SL g2182 ( 
.A(n_1922),
.Y(n_2182)
);

NAND2xp33_ASAP7_75t_L g2183 ( 
.A(n_1935),
.B(n_1262),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1902),
.B(n_1264),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1904),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1967),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1941),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1906),
.Y(n_2188)
);

BUFx3_ASAP7_75t_L g2189 ( 
.A(n_1949),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1983),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1907),
.Y(n_2191)
);

BUFx3_ASAP7_75t_L g2192 ( 
.A(n_1950),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1908),
.B(n_1267),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1909),
.B(n_1274),
.Y(n_2194)
);

BUFx3_ASAP7_75t_L g2195 ( 
.A(n_1954),
.Y(n_2195)
);

INVx3_ASAP7_75t_L g2196 ( 
.A(n_1956),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_1885),
.B(n_1289),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1848),
.B(n_1302),
.Y(n_2198)
);

BUFx10_ASAP7_75t_L g2199 ( 
.A(n_1853),
.Y(n_2199)
);

BUFx2_ASAP7_75t_L g2200 ( 
.A(n_1854),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_1885),
.B(n_1306),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1913),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1916),
.B(n_1309),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_L g2204 ( 
.A(n_1797),
.B(n_1823),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1918),
.B(n_1312),
.Y(n_2205)
);

AND2x2_ASAP7_75t_SL g2206 ( 
.A(n_1813),
.B(n_1375),
.Y(n_2206)
);

INVx5_ASAP7_75t_L g2207 ( 
.A(n_1944),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_1785),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_1960),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1925),
.B(n_1314),
.Y(n_2210)
);

INVx4_ASAP7_75t_L g2211 ( 
.A(n_1963),
.Y(n_2211)
);

INVx4_ASAP7_75t_L g2212 ( 
.A(n_1892),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1828),
.Y(n_2213)
);

INVx3_ASAP7_75t_L g2214 ( 
.A(n_1839),
.Y(n_2214)
);

INVx1_ASAP7_75t_SL g2215 ( 
.A(n_1812),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1845),
.Y(n_2216)
);

BUFx6f_ASAP7_75t_L g2217 ( 
.A(n_1812),
.Y(n_2217)
);

BUFx6f_ASAP7_75t_L g2218 ( 
.A(n_1939),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1849),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1850),
.Y(n_2220)
);

BUFx3_ASAP7_75t_L g2221 ( 
.A(n_1858),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_1793),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1953),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1939),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1796),
.B(n_1317),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1947),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1939),
.B(n_1320),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_L g2228 ( 
.A1(n_1952),
.A2(n_1332),
.B1(n_1333),
.B2(n_1325),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1958),
.B(n_1334),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1958),
.B(n_1335),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_1958),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1959),
.Y(n_2232)
);

NOR2xp33_ASAP7_75t_L g2233 ( 
.A(n_1961),
.B(n_1336),
.Y(n_2233)
);

BUFx3_ASAP7_75t_L g2234 ( 
.A(n_1943),
.Y(n_2234)
);

AOI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_1948),
.A2(n_1339),
.B1(n_1341),
.B2(n_1338),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_L g2236 ( 
.A(n_1957),
.B(n_1342),
.Y(n_2236)
);

INVx2_ASAP7_75t_SL g2237 ( 
.A(n_1962),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1910),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1910),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1772),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_1743),
.Y(n_2241)
);

AND2x6_ASAP7_75t_L g2242 ( 
.A(n_1820),
.B(n_986),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1817),
.B(n_1349),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_1847),
.A2(n_1352),
.B1(n_1354),
.B2(n_1350),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_1973),
.B(n_1355),
.Y(n_2245)
);

BUFx2_ASAP7_75t_L g2246 ( 
.A(n_1758),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1772),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_1743),
.Y(n_2248)
);

BUFx3_ASAP7_75t_L g2249 ( 
.A(n_1955),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_1973),
.B(n_1366),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_1743),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1743),
.Y(n_2252)
);

INVx4_ASAP7_75t_SL g2253 ( 
.A(n_1932),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1817),
.B(n_1368),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1910),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1817),
.B(n_1370),
.Y(n_2256)
);

INVx5_ASAP7_75t_L g2257 ( 
.A(n_1743),
.Y(n_2257)
);

AND2x4_ASAP7_75t_L g2258 ( 
.A(n_1758),
.B(n_1056),
.Y(n_2258)
);

INVx4_ASAP7_75t_L g2259 ( 
.A(n_1743),
.Y(n_2259)
);

BUFx4f_ASAP7_75t_L g2260 ( 
.A(n_1773),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_1825),
.B(n_1372),
.Y(n_2261)
);

INVx5_ASAP7_75t_L g2262 ( 
.A(n_1743),
.Y(n_2262)
);

BUFx4f_ASAP7_75t_L g2263 ( 
.A(n_1773),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1910),
.Y(n_2264)
);

OAI22xp5_ASAP7_75t_L g2265 ( 
.A1(n_1847),
.A2(n_1438),
.B1(n_1380),
.B2(n_1383),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_1973),
.B(n_1377),
.Y(n_2266)
);

INVx2_ASAP7_75t_SL g2267 ( 
.A(n_1743),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_1825),
.B(n_1385),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1973),
.B(n_1387),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_1743),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1817),
.B(n_1433),
.Y(n_2271)
);

INVx4_ASAP7_75t_L g2272 ( 
.A(n_1743),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1772),
.Y(n_2273)
);

AND2x6_ASAP7_75t_L g2274 ( 
.A(n_1820),
.B(n_986),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_1973),
.B(n_1392),
.Y(n_2275)
);

INVx6_ASAP7_75t_L g2276 ( 
.A(n_1743),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_1743),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_1743),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_1758),
.B(n_1066),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1973),
.B(n_1393),
.Y(n_2280)
);

BUFx3_ASAP7_75t_L g2281 ( 
.A(n_1955),
.Y(n_2281)
);

BUFx6f_ASAP7_75t_L g2282 ( 
.A(n_1743),
.Y(n_2282)
);

AND2x6_ASAP7_75t_L g2283 ( 
.A(n_1820),
.B(n_986),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_1825),
.B(n_1396),
.Y(n_2284)
);

OR2x2_ASAP7_75t_L g2285 ( 
.A(n_1765),
.B(n_1434),
.Y(n_2285)
);

AND2x2_ASAP7_75t_SL g2286 ( 
.A(n_1842),
.B(n_1411),
.Y(n_2286)
);

OR2x2_ASAP7_75t_L g2287 ( 
.A(n_1765),
.B(n_1436),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_1825),
.B(n_1395),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1772),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_1825),
.B(n_1398),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_1825),
.B(n_1397),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_L g2292 ( 
.A(n_1825),
.B(n_1402),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_1825),
.B(n_1408),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2041),
.B(n_1410),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2014),
.Y(n_2295)
);

INVxp67_ASAP7_75t_L g2296 ( 
.A(n_2002),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2075),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2015),
.Y(n_2298)
);

INVxp67_ASAP7_75t_L g2299 ( 
.A(n_2066),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2076),
.Y(n_2300)
);

NAND2xp33_ASAP7_75t_L g2301 ( 
.A(n_2100),
.B(n_1429),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1991),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1993),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2084),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1995),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2017),
.B(n_1421),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2017),
.B(n_1422),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2006),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2091),
.Y(n_2309)
);

AND2x4_ASAP7_75t_SL g2310 ( 
.A(n_2007),
.B(n_1130),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_L g2311 ( 
.A(n_2019),
.B(n_1423),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2009),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2012),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2027),
.Y(n_2314)
);

NAND2x1p5_ASAP7_75t_L g2315 ( 
.A(n_2257),
.B(n_1042),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2119),
.Y(n_2316)
);

AND2x4_ASAP7_75t_L g2317 ( 
.A(n_2257),
.B(n_1075),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2129),
.B(n_1427),
.Y(n_2318)
);

NAND2x1p5_ASAP7_75t_L g2319 ( 
.A(n_2262),
.B(n_1042),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2120),
.Y(n_2320)
);

NOR2xp67_ASAP7_75t_L g2321 ( 
.A(n_2262),
.B(n_1),
.Y(n_2321)
);

AO22x2_ASAP7_75t_L g2322 ( 
.A1(n_2090),
.A2(n_1347),
.B1(n_1351),
.B2(n_1345),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2020),
.B(n_1430),
.Y(n_2323)
);

AND2x4_ASAP7_75t_L g2324 ( 
.A(n_2007),
.B(n_1083),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1990),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_2241),
.B(n_949),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2133),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2145),
.Y(n_2328)
);

INVx5_ASAP7_75t_L g2329 ( 
.A(n_2241),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2238),
.Y(n_2330)
);

AO22x2_ASAP7_75t_L g2331 ( 
.A1(n_2021),
.A2(n_1364),
.B1(n_1369),
.B2(n_1361),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2239),
.Y(n_2332)
);

AND2x6_ASAP7_75t_L g2333 ( 
.A(n_2252),
.B(n_1411),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2255),
.Y(n_2334)
);

NOR2xp67_ASAP7_75t_L g2335 ( 
.A(n_2259),
.B(n_2),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2150),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_2050),
.Y(n_2337)
);

NOR2xp67_ASAP7_75t_L g2338 ( 
.A(n_2272),
.B(n_2),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2245),
.B(n_1189),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_2252),
.B(n_1084),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2264),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2163),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2250),
.B(n_1376),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2172),
.Y(n_2344)
);

INVxp67_ASAP7_75t_L g2345 ( 
.A(n_2270),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2266),
.B(n_1378),
.Y(n_2346)
);

OR2x6_ASAP7_75t_L g2347 ( 
.A(n_2044),
.B(n_1079),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2206),
.A2(n_955),
.B1(n_956),
.B2(n_950),
.Y(n_2348)
);

NAND2x1p5_ASAP7_75t_L g2349 ( 
.A(n_2270),
.B(n_2278),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2269),
.B(n_1390),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_2278),
.Y(n_2351)
);

INVx8_ASAP7_75t_L g2352 ( 
.A(n_2282),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2275),
.B(n_964),
.Y(n_2353)
);

AOI22xp33_ASAP7_75t_L g2354 ( 
.A1(n_2049),
.A2(n_981),
.B1(n_988),
.B2(n_968),
.Y(n_2354)
);

AO21x1_ASAP7_75t_L g2355 ( 
.A1(n_2169),
.A2(n_1414),
.B(n_1404),
.Y(n_2355)
);

OAI221xp5_ASAP7_75t_L g2356 ( 
.A1(n_2060),
.A2(n_995),
.B1(n_1001),
.B2(n_996),
.C(n_993),
.Y(n_2356)
);

AOI22xp33_ASAP7_75t_L g2357 ( 
.A1(n_2049),
.A2(n_1002),
.B1(n_1006),
.B2(n_1005),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2028),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2035),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_2282),
.B(n_1115),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2186),
.Y(n_2361)
);

OR2x2_ASAP7_75t_L g2362 ( 
.A(n_2175),
.B(n_1010),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2190),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2039),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2042),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2047),
.Y(n_2366)
);

BUFx8_ASAP7_75t_L g2367 ( 
.A(n_2008),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2053),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2055),
.Y(n_2369)
);

OAI22xp33_ASAP7_75t_L g2370 ( 
.A1(n_2156),
.A2(n_1016),
.B1(n_1019),
.B2(n_1015),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2058),
.Y(n_2371)
);

INVx2_ASAP7_75t_SL g2372 ( 
.A(n_2276),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2070),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2073),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2079),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2280),
.B(n_1415),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2083),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2101),
.B(n_1419),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_2089),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2064),
.B(n_1123),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2094),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2099),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2112),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_2064),
.B(n_1125),
.Y(n_2384)
);

NAND2xp33_ASAP7_75t_L g2385 ( 
.A(n_2137),
.B(n_1391),
.Y(n_2385)
);

OAI22xp33_ASAP7_75t_L g2386 ( 
.A1(n_2156),
.A2(n_1029),
.B1(n_1030),
.B2(n_1022),
.Y(n_2386)
);

NAND3xp33_ASAP7_75t_L g2387 ( 
.A(n_2056),
.B(n_1070),
.C(n_1042),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_L g2388 ( 
.A(n_2089),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2157),
.Y(n_2389)
);

NOR2xp67_ASAP7_75t_L g2390 ( 
.A(n_2018),
.B(n_3),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2126),
.Y(n_2391)
);

AO22x2_ASAP7_75t_L g2392 ( 
.A1(n_2253),
.A2(n_1432),
.B1(n_1420),
.B2(n_1129),
.Y(n_2392)
);

CKINVDCx16_ASAP7_75t_R g2393 ( 
.A(n_2077),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2225),
.B(n_1032),
.Y(n_2394)
);

AND2x4_ASAP7_75t_L g2395 ( 
.A(n_2253),
.B(n_1127),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2141),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_1989),
.B(n_1141),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2143),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2144),
.Y(n_2399)
);

AND2x6_ASAP7_75t_SL g2400 ( 
.A(n_2155),
.B(n_1143),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2146),
.Y(n_2401)
);

AND2x6_ASAP7_75t_L g2402 ( 
.A(n_2139),
.B(n_1042),
.Y(n_2402)
);

AO22x1_ASAP7_75t_L g2403 ( 
.A1(n_2102),
.A2(n_1039),
.B1(n_1046),
.B2(n_1033),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2148),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2151),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2036),
.B(n_1050),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2248),
.B(n_1144),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2165),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2115),
.B(n_1054),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_1992),
.Y(n_2410)
);

INVx3_ASAP7_75t_L g2411 ( 
.A(n_2063),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_1996),
.Y(n_2412)
);

AOI22xp33_ASAP7_75t_L g2413 ( 
.A1(n_2059),
.A2(n_1060),
.B1(n_1061),
.B2(n_1057),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2177),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_1999),
.Y(n_2415)
);

BUFx8_ASAP7_75t_L g2416 ( 
.A(n_2246),
.Y(n_2416)
);

BUFx3_ASAP7_75t_L g2417 ( 
.A(n_1988),
.Y(n_2417)
);

AO22x2_ASAP7_75t_L g2418 ( 
.A1(n_2051),
.A2(n_1152),
.B1(n_1155),
.B2(n_1149),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2249),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2162),
.Y(n_2420)
);

NOR3xp33_ASAP7_75t_L g2421 ( 
.A(n_2093),
.B(n_1179),
.C(n_1170),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2118),
.B(n_2170),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2134),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2142),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2003),
.Y(n_2425)
);

INVxp67_ASAP7_75t_L g2426 ( 
.A(n_2097),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2067),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2000),
.B(n_1077),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_2281),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2227),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2267),
.B(n_2277),
.Y(n_2431)
);

NOR2xp33_ASAP7_75t_L g2432 ( 
.A(n_2092),
.B(n_1087),
.Y(n_2432)
);

AOI22xp33_ASAP7_75t_L g2433 ( 
.A1(n_2179),
.A2(n_1090),
.B1(n_1097),
.B2(n_1096),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2025),
.Y(n_2434)
);

NAND2x1p5_ASAP7_75t_L g2435 ( 
.A(n_2251),
.B(n_1070),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2285),
.B(n_1105),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2229),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2230),
.Y(n_2438)
);

AO22x2_ASAP7_75t_L g2439 ( 
.A1(n_2215),
.A2(n_1193),
.B1(n_1199),
.B2(n_1180),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_2010),
.B(n_2088),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2005),
.B(n_1111),
.Y(n_2441)
);

AO22x2_ASAP7_75t_L g2442 ( 
.A1(n_2182),
.A2(n_1235),
.B1(n_1242),
.B2(n_1210),
.Y(n_2442)
);

BUFx2_ASAP7_75t_L g2443 ( 
.A(n_1987),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2136),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_2287),
.B(n_1120),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2268),
.B(n_2288),
.Y(n_2446)
);

AO22x2_ASAP7_75t_L g2447 ( 
.A1(n_2109),
.A2(n_1245),
.B1(n_1248),
.B2(n_1244),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2213),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2216),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2291),
.B(n_1122),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2219),
.Y(n_2451)
);

HB1xp67_ASAP7_75t_L g2452 ( 
.A(n_2200),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2087),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2046),
.Y(n_2454)
);

AO22x2_ASAP7_75t_L g2455 ( 
.A1(n_2114),
.A2(n_1265),
.B1(n_1268),
.B2(n_1257),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2164),
.Y(n_2456)
);

A2O1A1Ixp33_ASAP7_75t_L g2457 ( 
.A1(n_2158),
.A2(n_1279),
.B(n_1282),
.C(n_1269),
.Y(n_2457)
);

INVx4_ASAP7_75t_L g2458 ( 
.A(n_2044),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2240),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2110),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_2068),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2292),
.B(n_1128),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2160),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2247),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2293),
.B(n_1148),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2236),
.Y(n_2466)
);

AO22x2_ASAP7_75t_L g2467 ( 
.A1(n_2026),
.A2(n_1305),
.B1(n_1308),
.B2(n_1286),
.Y(n_2467)
);

NOR2xp67_ASAP7_75t_L g2468 ( 
.A(n_2048),
.B(n_3),
.Y(n_2468)
);

NAND2x1p5_ASAP7_75t_L g2469 ( 
.A(n_2081),
.B(n_1098),
.Y(n_2469)
);

OR2x2_ASAP7_75t_SL g2470 ( 
.A(n_2222),
.B(n_1425),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2166),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2001),
.Y(n_2472)
);

AND2x2_ASAP7_75t_SL g2473 ( 
.A(n_2004),
.B(n_1098),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2243),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2254),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2256),
.Y(n_2476)
);

CKINVDCx11_ASAP7_75t_R g2477 ( 
.A(n_1997),
.Y(n_2477)
);

NAND2x1p5_ASAP7_75t_L g2478 ( 
.A(n_2124),
.B(n_1098),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2273),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2271),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2289),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2244),
.B(n_1162),
.Y(n_2482)
);

AO22x2_ASAP7_75t_L g2483 ( 
.A1(n_1994),
.A2(n_1321),
.B1(n_1330),
.B2(n_1315),
.Y(n_2483)
);

INVxp67_ASAP7_75t_L g2484 ( 
.A(n_2030),
.Y(n_2484)
);

NAND2x1_ASAP7_75t_L g2485 ( 
.A(n_1987),
.B(n_2242),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2220),
.Y(n_2486)
);

AO22x2_ASAP7_75t_L g2487 ( 
.A1(n_1994),
.A2(n_1356),
.B1(n_1360),
.B2(n_1331),
.Y(n_2487)
);

BUFx2_ASAP7_75t_L g2488 ( 
.A(n_1987),
.Y(n_2488)
);

A2O1A1Ixp33_ASAP7_75t_L g2489 ( 
.A1(n_2159),
.A2(n_1379),
.B(n_1388),
.C(n_1374),
.Y(n_2489)
);

AND2x4_ASAP7_75t_L g2490 ( 
.A(n_2071),
.B(n_1389),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2103),
.B(n_1405),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2226),
.Y(n_2492)
);

NAND2xp33_ASAP7_75t_L g2493 ( 
.A(n_2137),
.B(n_1391),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2103),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2265),
.B(n_1178),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2103),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_L g2497 ( 
.A(n_2068),
.Y(n_2497)
);

AND2x6_ASAP7_75t_L g2498 ( 
.A(n_2139),
.B(n_1098),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_2116),
.Y(n_2499)
);

OAI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2125),
.A2(n_1186),
.B1(n_1191),
.B2(n_1185),
.Y(n_2500)
);

HB1xp67_ASAP7_75t_L g2501 ( 
.A(n_2061),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2232),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2135),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2217),
.Y(n_2504)
);

INVxp67_ASAP7_75t_L g2505 ( 
.A(n_2096),
.Y(n_2505)
);

NOR3xp33_ASAP7_75t_L g2506 ( 
.A(n_2037),
.B(n_1426),
.C(n_1406),
.Y(n_2506)
);

BUFx6f_ASAP7_75t_L g2507 ( 
.A(n_2072),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2260),
.B(n_1207),
.Y(n_2508)
);

BUFx8_ASAP7_75t_L g2509 ( 
.A(n_2031),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2233),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2217),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2223),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2197),
.B(n_1211),
.Y(n_2513)
);

INVx4_ASAP7_75t_L g2514 ( 
.A(n_1998),
.Y(n_2514)
);

AOI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2029),
.A2(n_1227),
.B1(n_1230),
.B2(n_1224),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2235),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2107),
.Y(n_2517)
);

NAND2x1p5_ASAP7_75t_L g2518 ( 
.A(n_2171),
.B(n_1114),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2107),
.Y(n_2519)
);

NAND3xp33_ASAP7_75t_L g2520 ( 
.A(n_2201),
.B(n_2062),
.C(n_2123),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2212),
.B(n_1428),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2174),
.Y(n_2522)
);

NAND2xp33_ASAP7_75t_L g2523 ( 
.A(n_2137),
.B(n_1391),
.Y(n_2523)
);

AND2x4_ASAP7_75t_L g2524 ( 
.A(n_2127),
.B(n_1079),
.Y(n_2524)
);

INVx1_ASAP7_75t_SL g2525 ( 
.A(n_2189),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2121),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2078),
.B(n_1238),
.Y(n_2527)
);

AO22x2_ASAP7_75t_L g2528 ( 
.A1(n_2022),
.A2(n_1167),
.B1(n_1197),
.B2(n_1113),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2045),
.B(n_1243),
.Y(n_2529)
);

INVx2_ASAP7_75t_SL g2530 ( 
.A(n_2263),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2121),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2122),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2178),
.Y(n_2533)
);

AO22x2_ASAP7_75t_L g2534 ( 
.A1(n_2161),
.A2(n_1167),
.B1(n_1197),
.B2(n_1113),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2080),
.B(n_1249),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2185),
.Y(n_2536)
);

INVx2_ASAP7_75t_SL g2537 ( 
.A(n_2199),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2188),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2117),
.B(n_1394),
.Y(n_2539)
);

NAND2x1p5_ASAP7_75t_L g2540 ( 
.A(n_2192),
.B(n_1114),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_L g2541 ( 
.A(n_2013),
.B(n_1250),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2191),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2122),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_SL g2544 ( 
.A(n_2054),
.B(n_1418),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2195),
.B(n_1323),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2202),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_2211),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2152),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2153),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2147),
.Y(n_2550)
);

AO22x2_ASAP7_75t_L g2551 ( 
.A1(n_2258),
.A2(n_1399),
.B1(n_1437),
.B2(n_1323),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2231),
.Y(n_2552)
);

INVx3_ASAP7_75t_L g2553 ( 
.A(n_2149),
.Y(n_2553)
);

BUFx6f_ASAP7_75t_L g2554 ( 
.A(n_2072),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2221),
.Y(n_2555)
);

INVxp67_ASAP7_75t_L g2556 ( 
.A(n_2198),
.Y(n_2556)
);

NAND2xp33_ASAP7_75t_L g2557 ( 
.A(n_2168),
.B(n_1391),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2016),
.B(n_1271),
.Y(n_2558)
);

INVx6_ASAP7_75t_L g2559 ( 
.A(n_2104),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2106),
.Y(n_2560)
);

INVx2_ASAP7_75t_SL g2561 ( 
.A(n_2132),
.Y(n_2561)
);

AOI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2057),
.A2(n_1276),
.B1(n_1280),
.B2(n_1275),
.Y(n_2562)
);

NAND2x1p5_ASAP7_75t_L g2563 ( 
.A(n_2095),
.B(n_1114),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_2261),
.B(n_1287),
.Y(n_2564)
);

NAND2x1p5_ASAP7_75t_L g2565 ( 
.A(n_2196),
.B(n_1114),
.Y(n_2565)
);

NAND2x1p5_ASAP7_75t_L g2566 ( 
.A(n_2128),
.B(n_1135),
.Y(n_2566)
);

AND2x4_ASAP7_75t_L g2567 ( 
.A(n_2209),
.B(n_1399),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2108),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2111),
.Y(n_2569)
);

INVxp67_ASAP7_75t_L g2570 ( 
.A(n_2279),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2184),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2193),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2194),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2203),
.B(n_1292),
.Y(n_2574)
);

BUFx8_ASAP7_75t_L g2575 ( 
.A(n_2140),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2205),
.B(n_1295),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2043),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2086),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2242),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2214),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2242),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2274),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_2105),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2274),
.Y(n_2584)
);

HB1xp67_ASAP7_75t_L g2585 ( 
.A(n_2098),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2284),
.B(n_1301),
.Y(n_2586)
);

INVx1_ASAP7_75t_SL g2587 ( 
.A(n_2038),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2224),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2274),
.Y(n_2589)
);

AO22x2_ASAP7_75t_L g2590 ( 
.A1(n_2176),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2590)
);

CKINVDCx11_ASAP7_75t_R g2591 ( 
.A(n_2082),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2283),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_2085),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2234),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2290),
.B(n_1303),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2283),
.Y(n_2596)
);

BUFx4f_ASAP7_75t_L g2597 ( 
.A(n_2023),
.Y(n_2597)
);

AND2x4_ASAP7_75t_L g2598 ( 
.A(n_2131),
.B(n_4),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2283),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2228),
.B(n_1304),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2207),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2052),
.Y(n_2602)
);

INVxp67_ASAP7_75t_L g2603 ( 
.A(n_2130),
.Y(n_2603)
);

INVxp67_ASAP7_75t_L g2604 ( 
.A(n_2210),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2207),
.Y(n_2605)
);

AO22x2_ASAP7_75t_L g2606 ( 
.A1(n_2180),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2154),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2173),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2183),
.Y(n_2609)
);

OR2x2_ASAP7_75t_L g2610 ( 
.A(n_2204),
.B(n_1310),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2011),
.B(n_7),
.Y(n_2611)
);

AO22x2_ASAP7_75t_L g2612 ( 
.A1(n_2069),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2208),
.A2(n_1324),
.B1(n_1326),
.B2(n_1316),
.Y(n_2613)
);

AND2x4_ASAP7_75t_L g2614 ( 
.A(n_2011),
.B(n_7),
.Y(n_2614)
);

INVxp67_ASAP7_75t_L g2615 ( 
.A(n_2113),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2237),
.Y(n_2616)
);

AO22x2_ASAP7_75t_L g2617 ( 
.A1(n_2074),
.A2(n_2034),
.B1(n_2040),
.B2(n_2032),
.Y(n_2617)
);

NAND2x1p5_ASAP7_75t_L g2618 ( 
.A(n_2033),
.B(n_2065),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2187),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2033),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2065),
.Y(n_2621)
);

BUFx6f_ASAP7_75t_L g2622 ( 
.A(n_2167),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2168),
.Y(n_2623)
);

INVx5_ASAP7_75t_L g2624 ( 
.A(n_2167),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_2181),
.B(n_1400),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2181),
.B(n_1343),
.Y(n_2626)
);

AO22x2_ASAP7_75t_L g2627 ( 
.A1(n_2090),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_2627)
);

NAND2x1p5_ASAP7_75t_L g2628 ( 
.A(n_2257),
.B(n_1135),
.Y(n_2628)
);

AND2x4_ASAP7_75t_SL g2629 ( 
.A(n_2007),
.B(n_1135),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2014),
.Y(n_2630)
);

AO22x2_ASAP7_75t_L g2631 ( 
.A1(n_2090),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2257),
.B(n_12),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2024),
.A2(n_1359),
.B1(n_1365),
.B2(n_1353),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2014),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2014),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2014),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2075),
.Y(n_2637)
);

INVxp67_ASAP7_75t_L g2638 ( 
.A(n_2002),
.Y(n_2638)
);

OAI221xp5_ASAP7_75t_L g2639 ( 
.A1(n_2019),
.A2(n_1381),
.B1(n_1382),
.B2(n_1373),
.C(n_1367),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2014),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_2041),
.B(n_1435),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2075),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2075),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2014),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2075),
.Y(n_2645)
);

OAI221xp5_ASAP7_75t_L g2646 ( 
.A1(n_2019),
.A2(n_1412),
.B1(n_1413),
.B2(n_1409),
.C(n_1401),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2014),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2014),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2075),
.Y(n_2649)
);

INVxp67_ASAP7_75t_L g2650 ( 
.A(n_2002),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2257),
.B(n_12),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2017),
.B(n_1391),
.Y(n_2652)
);

OAI22xp33_ASAP7_75t_L g2653 ( 
.A1(n_2019),
.A2(n_1228),
.B1(n_1313),
.B2(n_1209),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2014),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2014),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2014),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2257),
.B(n_12),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2024),
.B(n_13),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2014),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2075),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2075),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2014),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2014),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2017),
.B(n_13),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2014),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2014),
.Y(n_2666)
);

INVxp67_ASAP7_75t_SL g2667 ( 
.A(n_2007),
.Y(n_2667)
);

CKINVDCx20_ASAP7_75t_R g2668 ( 
.A(n_2138),
.Y(n_2668)
);

INVxp67_ASAP7_75t_L g2669 ( 
.A(n_2002),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2014),
.Y(n_2670)
);

AND2x4_ASAP7_75t_L g2671 ( 
.A(n_2257),
.B(n_15),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2014),
.Y(n_2672)
);

NAND2xp33_ASAP7_75t_L g2673 ( 
.A(n_2100),
.B(n_1209),
.Y(n_2673)
);

AO22x2_ASAP7_75t_L g2674 ( 
.A1(n_2090),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_R g2675 ( 
.A(n_2050),
.B(n_15),
.Y(n_2675)
);

INVxp67_ASAP7_75t_L g2676 ( 
.A(n_2002),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2075),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2024),
.B(n_17),
.Y(n_2678)
);

OAI221xp5_ASAP7_75t_L g2679 ( 
.A1(n_2019),
.A2(n_1313),
.B1(n_1340),
.B2(n_1228),
.C(n_1209),
.Y(n_2679)
);

INVxp67_ASAP7_75t_L g2680 ( 
.A(n_2002),
.Y(n_2680)
);

OAI21xp33_ASAP7_75t_L g2681 ( 
.A1(n_2101),
.A2(n_1313),
.B(n_1228),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2014),
.Y(n_2682)
);

OAI22xp5_ASAP7_75t_L g2683 ( 
.A1(n_2024),
.A2(n_1340),
.B1(n_1384),
.B2(n_1313),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2024),
.B(n_18),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2014),
.Y(n_2685)
);

AO22x2_ASAP7_75t_L g2686 ( 
.A1(n_2090),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2014),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2075),
.Y(n_2688)
);

NAND2x1p5_ASAP7_75t_L g2689 ( 
.A(n_2257),
.B(n_1340),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2014),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2014),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2075),
.Y(n_2692)
);

INVxp67_ASAP7_75t_L g2693 ( 
.A(n_2002),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2014),
.Y(n_2694)
);

AND2x6_ASAP7_75t_L g2695 ( 
.A(n_2024),
.B(n_1340),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2014),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2257),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_2019),
.B(n_20),
.Y(n_2698)
);

INVxp67_ASAP7_75t_L g2699 ( 
.A(n_2002),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2014),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2014),
.Y(n_2701)
);

HB1xp67_ASAP7_75t_L g2702 ( 
.A(n_2007),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2024),
.B(n_21),
.Y(n_2703)
);

BUFx8_ASAP7_75t_L g2704 ( 
.A(n_2007),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2075),
.Y(n_2705)
);

NAND2x1p5_ASAP7_75t_L g2706 ( 
.A(n_2257),
.B(n_1384),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_2007),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_L g2708 ( 
.A(n_2019),
.B(n_22),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2075),
.Y(n_2709)
);

AND2x6_ASAP7_75t_L g2710 ( 
.A(n_2024),
.B(n_1384),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2014),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_L g2712 ( 
.A(n_2019),
.B(n_22),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2014),
.Y(n_2713)
);

OR2x2_ASAP7_75t_SL g2714 ( 
.A(n_2019),
.B(n_1417),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2075),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_2257),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2014),
.Y(n_2717)
);

BUFx6f_ASAP7_75t_L g2718 ( 
.A(n_2007),
.Y(n_2718)
);

AND2x4_ASAP7_75t_L g2719 ( 
.A(n_2257),
.B(n_23),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2014),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2014),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2014),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2017),
.B(n_23),
.Y(n_2723)
);

NOR2xp33_ASAP7_75t_L g2724 ( 
.A(n_2019),
.B(n_24),
.Y(n_2724)
);

AO22x2_ASAP7_75t_L g2725 ( 
.A1(n_2090),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2024),
.B(n_24),
.Y(n_2726)
);

BUFx8_ASAP7_75t_L g2727 ( 
.A(n_2007),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2014),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2257),
.B(n_25),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_2050),
.Y(n_2730)
);

AO22x2_ASAP7_75t_L g2731 ( 
.A1(n_2090),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2075),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2014),
.Y(n_2733)
);

INVxp67_ASAP7_75t_L g2734 ( 
.A(n_2002),
.Y(n_2734)
);

AO22x2_ASAP7_75t_L g2735 ( 
.A1(n_2090),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2735)
);

AO22x2_ASAP7_75t_L g2736 ( 
.A1(n_2090),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2736)
);

OR2x6_ASAP7_75t_L g2737 ( 
.A(n_2044),
.B(n_1007),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2075),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2024),
.B(n_29),
.Y(n_2739)
);

INVx3_ASAP7_75t_L g2740 ( 
.A(n_2007),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2075),
.Y(n_2741)
);

INVxp67_ASAP7_75t_L g2742 ( 
.A(n_2002),
.Y(n_2742)
);

AO22x2_ASAP7_75t_L g2743 ( 
.A1(n_2090),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2075),
.Y(n_2744)
);

NAND2x1p5_ASAP7_75t_L g2745 ( 
.A(n_2257),
.B(n_1007),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2024),
.B(n_31),
.Y(n_2746)
);

INVxp67_ASAP7_75t_L g2747 ( 
.A(n_2002),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2019),
.B(n_32),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2024),
.B(n_33),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2041),
.B(n_1136),
.Y(n_2750)
);

BUFx6f_ASAP7_75t_L g2751 ( 
.A(n_2218),
.Y(n_2751)
);

NAND2x1p5_ASAP7_75t_L g2752 ( 
.A(n_2257),
.B(n_1136),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2075),
.Y(n_2753)
);

NAND3x1_ASAP7_75t_L g2754 ( 
.A(n_2019),
.B(n_33),
.C(n_34),
.Y(n_2754)
);

BUFx6f_ASAP7_75t_L g2755 ( 
.A(n_2007),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2017),
.B(n_34),
.Y(n_2756)
);

BUFx3_ASAP7_75t_L g2757 ( 
.A(n_2007),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2014),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2024),
.B(n_35),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2014),
.Y(n_2760)
);

AND2x6_ASAP7_75t_L g2761 ( 
.A(n_2024),
.B(n_1137),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2075),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2024),
.B(n_35),
.Y(n_2763)
);

NAND2xp33_ASAP7_75t_L g2764 ( 
.A(n_2100),
.B(n_1137),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2014),
.Y(n_2765)
);

AND2x4_ASAP7_75t_L g2766 ( 
.A(n_2257),
.B(n_35),
.Y(n_2766)
);

NAND2x1p5_ASAP7_75t_L g2767 ( 
.A(n_2257),
.B(n_1138),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2024),
.B(n_36),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2014),
.Y(n_2769)
);

NAND2x1p5_ASAP7_75t_L g2770 ( 
.A(n_2257),
.B(n_1159),
.Y(n_2770)
);

OAI22xp33_ASAP7_75t_L g2771 ( 
.A1(n_2019),
.A2(n_1165),
.B1(n_1169),
.B2(n_1159),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2024),
.B(n_36),
.Y(n_2772)
);

NOR2xp33_ASAP7_75t_L g2773 ( 
.A(n_2019),
.B(n_36),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2075),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2075),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2075),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2014),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2014),
.Y(n_2778)
);

NOR3xp33_ASAP7_75t_L g2779 ( 
.A(n_2019),
.B(n_39),
.C(n_38),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2014),
.Y(n_2780)
);

A2O1A1Ixp33_ASAP7_75t_L g2781 ( 
.A1(n_2101),
.A2(n_1169),
.B(n_1222),
.C(n_1165),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2014),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2014),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2014),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2075),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2014),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2014),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2024),
.B(n_37),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2014),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2017),
.B(n_37),
.Y(n_2790)
);

NAND2xp33_ASAP7_75t_L g2791 ( 
.A(n_2100),
.B(n_1169),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2024),
.B(n_37),
.Y(n_2792)
);

AOI22xp33_ASAP7_75t_L g2793 ( 
.A1(n_2286),
.A2(n_1417),
.B1(n_1222),
.B2(n_41),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2014),
.Y(n_2794)
);

NAND2x1p5_ASAP7_75t_L g2795 ( 
.A(n_2257),
.B(n_1222),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2014),
.Y(n_2796)
);

OAI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2024),
.A2(n_1417),
.B1(n_41),
.B2(n_38),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2024),
.B(n_40),
.Y(n_2798)
);

AND2x4_ASAP7_75t_L g2799 ( 
.A(n_2257),
.B(n_40),
.Y(n_2799)
);

AOI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2019),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_2800)
);

INVxp67_ASAP7_75t_L g2801 ( 
.A(n_2002),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2014),
.Y(n_2802)
);

OAI221xp5_ASAP7_75t_L g2803 ( 
.A1(n_2019),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.C(n_46),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2075),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2257),
.B(n_44),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2017),
.B(n_45),
.Y(n_2806)
);

AOI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2019),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2807)
);

AND2x4_ASAP7_75t_L g2808 ( 
.A(n_2257),
.B(n_47),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2322),
.B(n_48),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2446),
.B(n_49),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_L g2811 ( 
.A(n_2461),
.Y(n_2811)
);

AOI21x1_ASAP7_75t_L g2812 ( 
.A1(n_2439),
.A2(n_49),
.B(n_50),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_SL g2813 ( 
.A(n_2473),
.B(n_717),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2472),
.B(n_51),
.Y(n_2814)
);

AOI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2673),
.A2(n_52),
.B(n_53),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2322),
.B(n_52),
.Y(n_2816)
);

INVx1_ASAP7_75t_SL g2817 ( 
.A(n_2352),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_SL g2818 ( 
.A(n_2329),
.B(n_717),
.Y(n_2818)
);

BUFx3_ASAP7_75t_L g2819 ( 
.A(n_2704),
.Y(n_2819)
);

AOI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2764),
.A2(n_2791),
.B(n_2681),
.Y(n_2820)
);

BUFx12f_ASAP7_75t_L g2821 ( 
.A(n_2477),
.Y(n_2821)
);

INVx4_ASAP7_75t_L g2822 ( 
.A(n_2352),
.Y(n_2822)
);

INVx3_ASAP7_75t_L g2823 ( 
.A(n_2718),
.Y(n_2823)
);

NOR2xp67_ASAP7_75t_L g2824 ( 
.A(n_2329),
.B(n_53),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2378),
.A2(n_54),
.B(n_55),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2474),
.B(n_54),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2475),
.B(n_54),
.Y(n_2827)
);

BUFx12f_ASAP7_75t_L g2828 ( 
.A(n_2704),
.Y(n_2828)
);

NAND3xp33_ASAP7_75t_L g2829 ( 
.A(n_2520),
.B(n_56),
.C(n_57),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2504),
.A2(n_56),
.B(n_57),
.Y(n_2830)
);

AOI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2296),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2831)
);

AOI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2511),
.A2(n_58),
.B(n_59),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2476),
.B(n_60),
.Y(n_2833)
);

NAND3xp33_ASAP7_75t_L g2834 ( 
.A(n_2781),
.B(n_61),
.C(n_62),
.Y(n_2834)
);

AOI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_2385),
.A2(n_2523),
.B(n_2493),
.Y(n_2835)
);

OAI21xp33_ASAP7_75t_L g2836 ( 
.A1(n_2439),
.A2(n_61),
.B(n_62),
.Y(n_2836)
);

AND2x4_ASAP7_75t_L g2837 ( 
.A(n_2329),
.B(n_61),
.Y(n_2837)
);

AOI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2557),
.A2(n_63),
.B(n_64),
.Y(n_2838)
);

OAI21xp33_ASAP7_75t_L g2839 ( 
.A1(n_2421),
.A2(n_63),
.B(n_64),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2295),
.Y(n_2840)
);

A2O1A1Ixp33_ASAP7_75t_L g2841 ( 
.A1(n_2423),
.A2(n_2424),
.B(n_2708),
.C(n_2698),
.Y(n_2841)
);

AOI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2510),
.A2(n_65),
.B(n_66),
.Y(n_2842)
);

AOI22xp5_ASAP7_75t_L g2843 ( 
.A1(n_2801),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2480),
.B(n_67),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2344),
.A2(n_68),
.B(n_69),
.Y(n_2845)
);

AND2x4_ASAP7_75t_L g2846 ( 
.A(n_2755),
.B(n_70),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2453),
.B(n_71),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2298),
.Y(n_2848)
);

AOI22x1_ASAP7_75t_L g2849 ( 
.A1(n_2528),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_2849)
);

A2O1A1Ixp33_ASAP7_75t_L g2850 ( 
.A1(n_2712),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_2850)
);

NOR3xp33_ASAP7_75t_L g2851 ( 
.A(n_2440),
.B(n_74),
.C(n_75),
.Y(n_2851)
);

INVxp67_ASAP7_75t_L g2852 ( 
.A(n_2727),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2361),
.A2(n_75),
.B(n_76),
.Y(n_2853)
);

O2A1O1Ixp33_ASAP7_75t_L g2854 ( 
.A1(n_2457),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_2854)
);

A2O1A1Ixp33_ASAP7_75t_L g2855 ( 
.A1(n_2724),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_2855)
);

AOI21xp5_ASAP7_75t_L g2856 ( 
.A1(n_2363),
.A2(n_78),
.B(n_79),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2630),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2634),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2548),
.B(n_78),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2635),
.Y(n_2860)
);

AOI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2602),
.A2(n_80),
.B(n_81),
.Y(n_2861)
);

AOI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2638),
.A2(n_2650),
.B1(n_2676),
.B2(n_2669),
.Y(n_2862)
);

O2A1O1Ixp5_ASAP7_75t_L g2863 ( 
.A1(n_2355),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2549),
.B(n_82),
.Y(n_2864)
);

OR2x6_ASAP7_75t_L g2865 ( 
.A(n_2737),
.B(n_83),
.Y(n_2865)
);

BUFx4f_ASAP7_75t_L g2866 ( 
.A(n_2737),
.Y(n_2866)
);

AOI21xp5_ASAP7_75t_L g2867 ( 
.A1(n_2466),
.A2(n_84),
.B(n_85),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2636),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2516),
.B(n_84),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2316),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2750),
.A2(n_86),
.B(n_87),
.Y(n_2871)
);

OR2x2_ASAP7_75t_L g2872 ( 
.A(n_2680),
.B(n_87),
.Y(n_2872)
);

AOI21xp5_ASAP7_75t_L g2873 ( 
.A1(n_2320),
.A2(n_88),
.B(n_89),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_2755),
.B(n_718),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2327),
.A2(n_88),
.B(n_89),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2478),
.B(n_719),
.Y(n_2876)
);

AOI21xp5_ASAP7_75t_L g2877 ( 
.A1(n_2328),
.A2(n_2342),
.B(n_2336),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2297),
.A2(n_2304),
.B(n_2300),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2804),
.A2(n_90),
.B(n_91),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2571),
.B(n_2572),
.Y(n_2880)
);

HB1xp67_ASAP7_75t_L g2881 ( 
.A(n_2501),
.Y(n_2881)
);

AOI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2693),
.A2(n_95),
.B1(n_92),
.B2(n_93),
.Y(n_2882)
);

AOI21xp5_ASAP7_75t_L g2883 ( 
.A1(n_2309),
.A2(n_93),
.B(n_95),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2573),
.B(n_96),
.Y(n_2884)
);

BUFx12f_ASAP7_75t_L g2885 ( 
.A(n_2591),
.Y(n_2885)
);

O2A1O1Ixp33_ASAP7_75t_L g2886 ( 
.A1(n_2489),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2366),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2664),
.B(n_100),
.Y(n_2888)
);

INVx3_ASAP7_75t_L g2889 ( 
.A(n_2565),
.Y(n_2889)
);

AOI21xp5_ASAP7_75t_L g2890 ( 
.A1(n_2637),
.A2(n_101),
.B(n_102),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2640),
.Y(n_2891)
);

NOR2x1_ASAP7_75t_L g2892 ( 
.A(n_2668),
.B(n_103),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_SL g2893 ( 
.A(n_2458),
.B(n_103),
.Y(n_2893)
);

AOI21x1_ASAP7_75t_L g2894 ( 
.A1(n_2623),
.A2(n_103),
.B(n_104),
.Y(n_2894)
);

AOI21x1_ASAP7_75t_L g2895 ( 
.A1(n_2579),
.A2(n_105),
.B(n_106),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2714),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2374),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2723),
.B(n_107),
.Y(n_2898)
);

AOI21xp5_ASAP7_75t_L g2899 ( 
.A1(n_2642),
.A2(n_107),
.B(n_108),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2756),
.B(n_108),
.Y(n_2900)
);

INVx4_ASAP7_75t_L g2901 ( 
.A(n_2559),
.Y(n_2901)
);

BUFx2_ASAP7_75t_L g2902 ( 
.A(n_2333),
.Y(n_2902)
);

AOI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2643),
.A2(n_109),
.B(n_110),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2375),
.Y(n_2904)
);

INVx2_ASAP7_75t_SL g2905 ( 
.A(n_2559),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2645),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2644),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2649),
.A2(n_109),
.B(n_110),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2422),
.B(n_109),
.Y(n_2909)
);

AOI21xp5_ASAP7_75t_L g2910 ( 
.A1(n_2660),
.A2(n_111),
.B(n_112),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2647),
.Y(n_2911)
);

AOI21x1_ASAP7_75t_L g2912 ( 
.A1(n_2581),
.A2(n_111),
.B(n_112),
.Y(n_2912)
);

O2A1O1Ixp33_ASAP7_75t_L g2913 ( 
.A1(n_2779),
.A2(n_114),
.B(n_111),
.C(n_113),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2648),
.Y(n_2914)
);

INVx1_ASAP7_75t_SL g2915 ( 
.A(n_2707),
.Y(n_2915)
);

INVx3_ASAP7_75t_L g2916 ( 
.A(n_2435),
.Y(n_2916)
);

BUFx12f_ASAP7_75t_L g2917 ( 
.A(n_2509),
.Y(n_2917)
);

NOR2x1_ASAP7_75t_L g2918 ( 
.A(n_2499),
.B(n_115),
.Y(n_2918)
);

AOI22xp5_ASAP7_75t_L g2919 ( 
.A1(n_2699),
.A2(n_2742),
.B1(n_2747),
.B2(n_2734),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2661),
.A2(n_116),
.B(n_117),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2677),
.A2(n_116),
.B(n_118),
.Y(n_2921)
);

OR2x2_ASAP7_75t_L g2922 ( 
.A(n_2426),
.B(n_116),
.Y(n_2922)
);

NAND3xp33_ASAP7_75t_L g2923 ( 
.A(n_2387),
.B(n_118),
.C(n_119),
.Y(n_2923)
);

BUFx12f_ASAP7_75t_L g2924 ( 
.A(n_2509),
.Y(n_2924)
);

O2A1O1Ixp33_ASAP7_75t_L g2925 ( 
.A1(n_2604),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_2925)
);

AOI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2688),
.A2(n_119),
.B(n_120),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2790),
.B(n_120),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2443),
.B(n_720),
.Y(n_2928)
);

BUFx12f_ASAP7_75t_L g2929 ( 
.A(n_2367),
.Y(n_2929)
);

O2A1O1Ixp33_ASAP7_75t_L g2930 ( 
.A1(n_2318),
.A2(n_126),
.B(n_123),
.C(n_124),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2556),
.B(n_2505),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2692),
.A2(n_2709),
.B(n_2705),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2806),
.B(n_123),
.Y(n_2933)
);

OAI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2658),
.A2(n_123),
.B(n_124),
.Y(n_2934)
);

O2A1O1Ixp33_ASAP7_75t_L g2935 ( 
.A1(n_2748),
.A2(n_129),
.B(n_126),
.C(n_127),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2715),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2654),
.B(n_129),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2732),
.A2(n_130),
.B(n_131),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2738),
.A2(n_132),
.B(n_133),
.Y(n_2939)
);

HB1xp67_ASAP7_75t_L g2940 ( 
.A(n_2757),
.Y(n_2940)
);

OAI21xp33_ASAP7_75t_SL g2941 ( 
.A1(n_2678),
.A2(n_132),
.B(n_133),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2655),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2656),
.B(n_134),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2659),
.B(n_134),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2662),
.B(n_135),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2663),
.B(n_137),
.Y(n_2946)
);

BUFx3_ASAP7_75t_L g2947 ( 
.A(n_2349),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2665),
.B(n_2666),
.Y(n_2948)
);

AOI21x1_ASAP7_75t_L g2949 ( 
.A1(n_2582),
.A2(n_137),
.B(n_138),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2741),
.A2(n_138),
.B(n_139),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_2744),
.A2(n_2762),
.B(n_2753),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2670),
.B(n_140),
.Y(n_2952)
);

BUFx3_ASAP7_75t_L g2953 ( 
.A(n_2707),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2672),
.Y(n_2954)
);

O2A1O1Ixp5_ASAP7_75t_L g2955 ( 
.A1(n_2485),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_2603),
.B(n_2570),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2353),
.B(n_141),
.Y(n_2957)
);

A2O1A1Ixp33_ASAP7_75t_L g2958 ( 
.A1(n_2773),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2428),
.B(n_143),
.Y(n_2959)
);

NOR2x1_ASAP7_75t_L g2960 ( 
.A(n_2514),
.B(n_144),
.Y(n_2960)
);

A2O1A1Ixp33_ASAP7_75t_L g2961 ( 
.A1(n_2430),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2961)
);

O2A1O1Ixp5_ASAP7_75t_L g2962 ( 
.A1(n_2485),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_2962)
);

NOR2xp33_ASAP7_75t_L g2963 ( 
.A(n_2299),
.B(n_148),
.Y(n_2963)
);

NOR3xp33_ASAP7_75t_L g2964 ( 
.A(n_2803),
.B(n_149),
.C(n_150),
.Y(n_2964)
);

AND2x4_ASAP7_75t_L g2965 ( 
.A(n_2414),
.B(n_150),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2682),
.B(n_2685),
.Y(n_2966)
);

AND2x2_ASAP7_75t_L g2967 ( 
.A(n_2441),
.B(n_151),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_SL g2968 ( 
.A(n_2337),
.B(n_152),
.Y(n_2968)
);

OAI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2684),
.A2(n_152),
.B(n_153),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2687),
.B(n_154),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_2393),
.Y(n_2971)
);

NAND2x1p5_ASAP7_75t_L g2972 ( 
.A(n_2597),
.B(n_154),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2443),
.B(n_721),
.Y(n_2973)
);

O2A1O1Ixp5_ASAP7_75t_L g2974 ( 
.A1(n_2653),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2690),
.B(n_2691),
.Y(n_2975)
);

O2A1O1Ixp5_ASAP7_75t_L g2976 ( 
.A1(n_2771),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_2379),
.Y(n_2977)
);

OAI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2793),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2461),
.Y(n_2979)
);

AOI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2774),
.A2(n_160),
.B(n_161),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2615),
.B(n_2484),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2775),
.Y(n_2982)
);

OAI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2331),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2776),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2785),
.A2(n_164),
.B(n_165),
.Y(n_2985)
);

HB1xp67_ASAP7_75t_L g2986 ( 
.A(n_2452),
.Y(n_2986)
);

AOI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2703),
.A2(n_164),
.B(n_165),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2694),
.B(n_2802),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2696),
.B(n_165),
.Y(n_2989)
);

OAI21xp33_ASAP7_75t_L g2990 ( 
.A1(n_2311),
.A2(n_166),
.B(n_167),
.Y(n_2990)
);

NAND2x1_ASAP7_75t_L g2991 ( 
.A(n_2695),
.B(n_166),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2700),
.B(n_167),
.Y(n_2992)
);

A2O1A1Ixp33_ASAP7_75t_L g2993 ( 
.A1(n_2437),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_2993)
);

A2O1A1Ixp33_ASAP7_75t_L g2994 ( 
.A1(n_2438),
.A2(n_171),
.B(n_168),
.C(n_170),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2398),
.Y(n_2995)
);

OAI21xp33_ASAP7_75t_L g2996 ( 
.A1(n_2323),
.A2(n_170),
.B(n_171),
.Y(n_2996)
);

NAND3xp33_ASAP7_75t_L g2997 ( 
.A(n_2679),
.B(n_170),
.C(n_172),
.Y(n_2997)
);

INVx1_ASAP7_75t_SL g2998 ( 
.A(n_2525),
.Y(n_2998)
);

AOI21xp5_ASAP7_75t_L g2999 ( 
.A1(n_2726),
.A2(n_172),
.B(n_173),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2701),
.Y(n_3000)
);

AOI21x1_ASAP7_75t_L g3001 ( 
.A1(n_2584),
.A2(n_174),
.B(n_175),
.Y(n_3001)
);

BUFx2_ASAP7_75t_L g3002 ( 
.A(n_2333),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2362),
.B(n_175),
.Y(n_3003)
);

AOI21xp5_ASAP7_75t_L g3004 ( 
.A1(n_2739),
.A2(n_176),
.B(n_177),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2461),
.Y(n_3005)
);

A2O1A1Ixp33_ASAP7_75t_L g3006 ( 
.A1(n_2746),
.A2(n_178),
.B(n_176),
.C(n_177),
.Y(n_3006)
);

NOR2xp33_ASAP7_75t_L g3007 ( 
.A(n_2610),
.B(n_176),
.Y(n_3007)
);

NOR2xp67_ASAP7_75t_L g3008 ( 
.A(n_2697),
.B(n_177),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2711),
.Y(n_3009)
);

AND2x6_ASAP7_75t_SL g3010 ( 
.A(n_2347),
.B(n_178),
.Y(n_3010)
);

OA22x2_ASAP7_75t_L g3011 ( 
.A1(n_2347),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_3011)
);

AOI21xp5_ASAP7_75t_L g3012 ( 
.A1(n_2749),
.A2(n_179),
.B(n_181),
.Y(n_3012)
);

INVx3_ASAP7_75t_L g3013 ( 
.A(n_2379),
.Y(n_3013)
);

O2A1O1Ixp5_ASAP7_75t_L g3014 ( 
.A1(n_2596),
.A2(n_2589),
.B(n_2599),
.C(n_2592),
.Y(n_3014)
);

A2O1A1Ixp33_ASAP7_75t_L g3015 ( 
.A1(n_2759),
.A2(n_2768),
.B(n_2772),
.C(n_2763),
.Y(n_3015)
);

OAI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2788),
.A2(n_181),
.B(n_182),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2713),
.B(n_182),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2399),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2717),
.B(n_2789),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2720),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2792),
.A2(n_183),
.B(n_184),
.Y(n_3021)
);

AOI21xp5_ASAP7_75t_L g3022 ( 
.A1(n_2798),
.A2(n_185),
.B(n_186),
.Y(n_3022)
);

AOI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2410),
.A2(n_187),
.B(n_188),
.Y(n_3023)
);

AO21x1_ASAP7_75t_L g3024 ( 
.A1(n_2797),
.A2(n_722),
.B(n_721),
.Y(n_3024)
);

AOI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2412),
.A2(n_2425),
.B(n_2415),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2721),
.B(n_188),
.Y(n_3026)
);

BUFx2_ASAP7_75t_SL g3027 ( 
.A(n_2716),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_SL g3028 ( 
.A(n_2488),
.B(n_722),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2722),
.B(n_2728),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_L g3030 ( 
.A(n_2356),
.B(n_2306),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_SL g3031 ( 
.A(n_2488),
.B(n_723),
.Y(n_3031)
);

AOI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2434),
.A2(n_189),
.B(n_190),
.Y(n_3032)
);

AOI21xp5_ASAP7_75t_L g3033 ( 
.A1(n_2454),
.A2(n_2464),
.B(n_2459),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2447),
.B(n_190),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2401),
.Y(n_3035)
);

NOR2xp33_ASAP7_75t_SL g3036 ( 
.A(n_2730),
.B(n_191),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2733),
.B(n_191),
.Y(n_3037)
);

O2A1O1Ixp33_ASAP7_75t_L g3038 ( 
.A1(n_2307),
.A2(n_194),
.B(n_192),
.C(n_193),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2518),
.B(n_727),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2758),
.B(n_2794),
.Y(n_3040)
);

AOI21x1_ASAP7_75t_L g3041 ( 
.A1(n_2494),
.A2(n_193),
.B(n_194),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2436),
.A2(n_2445),
.B1(n_2462),
.B2(n_2394),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2302),
.Y(n_3043)
);

INVxp67_ASAP7_75t_SL g3044 ( 
.A(n_2751),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2760),
.B(n_2780),
.Y(n_3045)
);

AOI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2479),
.A2(n_195),
.B(n_196),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2481),
.A2(n_196),
.B(n_197),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2765),
.B(n_2796),
.Y(n_3048)
);

AOI22x1_ASAP7_75t_L g3049 ( 
.A1(n_2315),
.A2(n_2319),
.B1(n_2689),
.B2(n_2628),
.Y(n_3049)
);

AO32x2_ASAP7_75t_L g3050 ( 
.A1(n_2683),
.A2(n_202),
.A3(n_199),
.B1(n_201),
.B2(n_203),
.Y(n_3050)
);

OAI21xp33_ASAP7_75t_L g3051 ( 
.A1(n_2339),
.A2(n_202),
.B(n_203),
.Y(n_3051)
);

AND2x4_ASAP7_75t_L g3052 ( 
.A(n_2667),
.B(n_204),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2769),
.B(n_204),
.Y(n_3053)
);

HB1xp67_ASAP7_75t_L g3054 ( 
.A(n_2702),
.Y(n_3054)
);

NOR2xp33_ASAP7_75t_L g3055 ( 
.A(n_2639),
.B(n_204),
.Y(n_3055)
);

OAI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_2343),
.A2(n_205),
.B(n_206),
.Y(n_3056)
);

AOI21x1_ASAP7_75t_L g3057 ( 
.A1(n_2496),
.A2(n_205),
.B(n_207),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_SL g3058 ( 
.A(n_2540),
.B(n_727),
.Y(n_3058)
);

OAI22xp5_ASAP7_75t_L g3059 ( 
.A1(n_2433),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_3059)
);

AOI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2497),
.A2(n_207),
.B(n_208),
.Y(n_3060)
);

A2O1A1Ixp33_ASAP7_75t_L g3061 ( 
.A1(n_2652),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2777),
.Y(n_3062)
);

OAI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2346),
.A2(n_212),
.B(n_213),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2778),
.B(n_212),
.Y(n_3064)
);

OR2x2_ASAP7_75t_L g3065 ( 
.A(n_2470),
.B(n_213),
.Y(n_3065)
);

AOI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2507),
.A2(n_214),
.B(n_215),
.Y(n_3066)
);

AOI21x1_ASAP7_75t_L g3067 ( 
.A1(n_2612),
.A2(n_214),
.B(n_215),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2303),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2782),
.Y(n_3069)
);

A2O1A1Ixp33_ASAP7_75t_L g3070 ( 
.A1(n_2800),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_3070)
);

AND2x4_ASAP7_75t_L g3071 ( 
.A(n_2351),
.B(n_216),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_2646),
.B(n_217),
.Y(n_3072)
);

AOI21xp5_ASAP7_75t_L g3073 ( 
.A1(n_2507),
.A2(n_218),
.B(n_219),
.Y(n_3073)
);

BUFx12f_ASAP7_75t_L g3074 ( 
.A(n_2416),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2783),
.Y(n_3075)
);

INVx4_ASAP7_75t_L g3076 ( 
.A(n_2740),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2784),
.B(n_2786),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2554),
.A2(n_2588),
.B(n_2376),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2787),
.B(n_2305),
.Y(n_3079)
);

AOI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2350),
.A2(n_220),
.B(n_221),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_2294),
.B(n_220),
.Y(n_3081)
);

OAI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_2392),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2308),
.B(n_225),
.Y(n_3083)
);

OAI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_2392),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_3084)
);

AOI21x1_ASAP7_75t_L g3085 ( 
.A1(n_2612),
.A2(n_229),
.B(n_230),
.Y(n_3085)
);

O2A1O1Ixp33_ASAP7_75t_L g3086 ( 
.A1(n_2409),
.A2(n_232),
.B(n_229),
.C(n_231),
.Y(n_3086)
);

A2O1A1Ixp33_ASAP7_75t_L g3087 ( 
.A1(n_2807),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_2535),
.B(n_2432),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2312),
.B(n_233),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2313),
.B(n_234),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2325),
.B(n_235),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2330),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_SL g3093 ( 
.A(n_2397),
.B(n_728),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2332),
.B(n_236),
.Y(n_3094)
);

O2A1O1Ixp5_ASAP7_75t_L g3095 ( 
.A1(n_2625),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2751),
.Y(n_3096)
);

AO21x1_ASAP7_75t_L g3097 ( 
.A1(n_2491),
.A2(n_729),
.B(n_728),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2397),
.B(n_731),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2609),
.A2(n_2449),
.B(n_2448),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2451),
.A2(n_239),
.B(n_240),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2334),
.B(n_241),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2460),
.B(n_241),
.Y(n_3102)
);

AOI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2486),
.A2(n_241),
.B(n_242),
.Y(n_3103)
);

BUFx4f_ASAP7_75t_L g3104 ( 
.A(n_2695),
.Y(n_3104)
);

BUFx6f_ASAP7_75t_L g3105 ( 
.A(n_2751),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2314),
.A2(n_245),
.B(n_247),
.Y(n_3106)
);

OR2x6_ASAP7_75t_L g3107 ( 
.A(n_2530),
.B(n_247),
.Y(n_3107)
);

INVx3_ASAP7_75t_L g3108 ( 
.A(n_2388),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2341),
.B(n_248),
.Y(n_3109)
);

AO21x1_ASAP7_75t_L g3110 ( 
.A1(n_2491),
.A2(n_733),
.B(n_732),
.Y(n_3110)
);

O2A1O1Ixp5_ASAP7_75t_L g3111 ( 
.A1(n_2539),
.A2(n_2567),
.B(n_2384),
.C(n_2395),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2492),
.A2(n_249),
.B(n_250),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_2407),
.B(n_734),
.Y(n_3113)
);

AND2x2_ASAP7_75t_SL g3114 ( 
.A(n_2301),
.B(n_249),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2358),
.Y(n_3115)
);

OAI21xp5_ASAP7_75t_L g3116 ( 
.A1(n_2574),
.A2(n_2576),
.B(n_2558),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2502),
.A2(n_252),
.B(n_253),
.Y(n_3117)
);

BUFx6f_ASAP7_75t_L g3118 ( 
.A(n_2388),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2359),
.A2(n_2365),
.B(n_2364),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_SL g3120 ( 
.A(n_2407),
.B(n_734),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2370),
.B(n_254),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2386),
.B(n_254),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_SL g3123 ( 
.A1(n_2706),
.A2(n_255),
.B(n_256),
.Y(n_3123)
);

OAI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2527),
.A2(n_255),
.B(n_256),
.Y(n_3124)
);

A2O1A1Ixp33_ASAP7_75t_L g3125 ( 
.A1(n_2368),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2369),
.Y(n_3126)
);

BUFx4f_ASAP7_75t_L g3127 ( 
.A(n_2695),
.Y(n_3127)
);

AND2x6_ASAP7_75t_L g3128 ( 
.A(n_2531),
.B(n_257),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2408),
.B(n_2371),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2373),
.B(n_258),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2377),
.B(n_258),
.Y(n_3131)
);

AOI21xp5_ASAP7_75t_L g3132 ( 
.A1(n_2381),
.A2(n_258),
.B(n_259),
.Y(n_3132)
);

BUFx6f_ASAP7_75t_L g3133 ( 
.A(n_2531),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2382),
.Y(n_3134)
);

INVxp67_ASAP7_75t_SL g3135 ( 
.A(n_2629),
.Y(n_3135)
);

OAI321xp33_ASAP7_75t_L g3136 ( 
.A1(n_2348),
.A2(n_261),
.A3(n_263),
.B1(n_259),
.B2(n_260),
.C(n_262),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_2335),
.B(n_735),
.Y(n_3137)
);

OAI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2383),
.A2(n_262),
.B(n_263),
.Y(n_3138)
);

AOI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_2389),
.A2(n_264),
.B(n_265),
.Y(n_3139)
);

INVx2_ASAP7_75t_SL g3140 ( 
.A(n_2431),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2338),
.B(n_736),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2391),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_2396),
.A2(n_266),
.B(n_267),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2404),
.Y(n_3144)
);

OAI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2405),
.A2(n_266),
.B(n_267),
.Y(n_3145)
);

OAI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_2551),
.A2(n_272),
.B1(n_269),
.B2(n_270),
.Y(n_3146)
);

INVxp67_ASAP7_75t_L g3147 ( 
.A(n_2534),
.Y(n_3147)
);

OAI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_2551),
.A2(n_272),
.B1(n_269),
.B2(n_270),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_2455),
.B(n_269),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2420),
.Y(n_3150)
);

AOI21xp5_ASAP7_75t_L g3151 ( 
.A1(n_2544),
.A2(n_270),
.B(n_272),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2419),
.B(n_273),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_2675),
.B(n_736),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2522),
.B(n_274),
.Y(n_3154)
);

AOI21xp5_ASAP7_75t_L g3155 ( 
.A1(n_2580),
.A2(n_274),
.B(n_275),
.Y(n_3155)
);

A2O1A1Ixp33_ASAP7_75t_L g3156 ( 
.A1(n_2390),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2533),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2512),
.Y(n_3158)
);

OR2x6_ASAP7_75t_L g3159 ( 
.A(n_2632),
.B(n_276),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2536),
.B(n_276),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2471),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2538),
.B(n_277),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2542),
.B(n_278),
.Y(n_3163)
);

NOR2xp33_ASAP7_75t_L g3164 ( 
.A(n_2429),
.B(n_278),
.Y(n_3164)
);

AOI21xp33_ASAP7_75t_L g3165 ( 
.A1(n_2406),
.A2(n_279),
.B(n_280),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2546),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2513),
.B(n_2560),
.Y(n_3167)
);

BUFx2_ASAP7_75t_L g3168 ( 
.A(n_2416),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_2526),
.A2(n_2543),
.B(n_2532),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2568),
.B(n_2569),
.Y(n_3170)
);

AOI21xp5_ASAP7_75t_L g3171 ( 
.A1(n_2616),
.A2(n_2456),
.B(n_2552),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2577),
.B(n_279),
.Y(n_3172)
);

BUFx2_ASAP7_75t_SL g3173 ( 
.A(n_2537),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2578),
.B(n_280),
.Y(n_3174)
);

BUFx4f_ASAP7_75t_L g3175 ( 
.A(n_2710),
.Y(n_3175)
);

AOI21x1_ASAP7_75t_L g3176 ( 
.A1(n_2617),
.A2(n_281),
.B(n_282),
.Y(n_3176)
);

OAI22xp5_ASAP7_75t_L g3177 ( 
.A1(n_2418),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_3177)
);

O2A1O1Ixp33_ASAP7_75t_L g3178 ( 
.A1(n_2506),
.A2(n_283),
.B(n_281),
.C(n_282),
.Y(n_3178)
);

OAI21xp33_ASAP7_75t_L g3179 ( 
.A1(n_2418),
.A2(n_283),
.B(n_284),
.Y(n_3179)
);

BUFx8_ASAP7_75t_L g3180 ( 
.A(n_2429),
.Y(n_3180)
);

AOI21xp5_ASAP7_75t_L g3181 ( 
.A1(n_2444),
.A2(n_2608),
.B(n_2607),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2450),
.B(n_285),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_2632),
.B(n_2651),
.Y(n_3183)
);

OAI22xp5_ASAP7_75t_L g3184 ( 
.A1(n_2483),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_3184)
);

NAND3xp33_ASAP7_75t_L g3185 ( 
.A(n_2468),
.B(n_287),
.C(n_288),
.Y(n_3185)
);

BUFx2_ASAP7_75t_L g3186 ( 
.A(n_2575),
.Y(n_3186)
);

AOI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_2503),
.A2(n_2463),
.B(n_2594),
.Y(n_3187)
);

AND2x2_ASAP7_75t_SL g3188 ( 
.A(n_2651),
.B(n_289),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2555),
.A2(n_290),
.B(n_291),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2606),
.Y(n_3190)
);

AOI22xp5_ASAP7_75t_L g3191 ( 
.A1(n_2465),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_3191)
);

AOI21xp5_ASAP7_75t_L g3192 ( 
.A1(n_2641),
.A2(n_293),
.B(n_294),
.Y(n_3192)
);

HB1xp67_ASAP7_75t_L g3193 ( 
.A(n_2345),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2606),
.Y(n_3194)
);

OAI21x1_ASAP7_75t_L g3195 ( 
.A1(n_2745),
.A2(n_295),
.B(n_296),
.Y(n_3195)
);

AOI21xp5_ASAP7_75t_L g3196 ( 
.A1(n_2626),
.A2(n_297),
.B(n_298),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2529),
.B(n_297),
.Y(n_3197)
);

INVx4_ASAP7_75t_L g3198 ( 
.A(n_2624),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_2575),
.Y(n_3199)
);

A2O1A1Ixp33_ASAP7_75t_L g3200 ( 
.A1(n_2598),
.A2(n_299),
.B(n_297),
.C(n_298),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2590),
.Y(n_3201)
);

AOI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_2600),
.A2(n_298),
.B(n_299),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2354),
.B(n_299),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2357),
.B(n_300),
.Y(n_3204)
);

INVxp67_ASAP7_75t_L g3205 ( 
.A(n_2324),
.Y(n_3205)
);

O2A1O1Ixp33_ASAP7_75t_L g3206 ( 
.A1(n_2482),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2431),
.B(n_303),
.Y(n_3207)
);

AOI21xp5_ASAP7_75t_L g3208 ( 
.A1(n_2495),
.A2(n_303),
.B(n_304),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2710),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2500),
.B(n_305),
.Y(n_3210)
);

INVx4_ASAP7_75t_L g3211 ( 
.A(n_2624),
.Y(n_3211)
);

NOR2xp67_ASAP7_75t_SL g3212 ( 
.A(n_2550),
.B(n_2553),
.Y(n_3212)
);

OAI21x1_ASAP7_75t_L g3213 ( 
.A1(n_2752),
.A2(n_306),
.B(n_307),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2633),
.B(n_307),
.Y(n_3214)
);

A2O1A1Ixp33_ASAP7_75t_L g3215 ( 
.A1(n_2321),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_3215)
);

AOI221xp5_ASAP7_75t_L g3216 ( 
.A1(n_2487),
.A2(n_2467),
.B1(n_2442),
.B2(n_2567),
.C(n_2490),
.Y(n_3216)
);

A2O1A1Ixp33_ASAP7_75t_L g3217 ( 
.A1(n_2611),
.A2(n_315),
.B(n_313),
.C(n_314),
.Y(n_3217)
);

AOI22x1_ASAP7_75t_L g3218 ( 
.A1(n_2469),
.A2(n_317),
.B1(n_314),
.B2(n_316),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2541),
.B(n_2564),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_2590),
.A2(n_316),
.B(n_317),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2627),
.Y(n_3221)
);

A2O1A1Ixp33_ASAP7_75t_L g3222 ( 
.A1(n_2611),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_3222)
);

A2O1A1Ixp33_ASAP7_75t_L g3223 ( 
.A1(n_2614),
.A2(n_2490),
.B(n_2384),
.C(n_2395),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_SL g3224 ( 
.A(n_2657),
.B(n_2671),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2413),
.B(n_319),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2442),
.B(n_320),
.Y(n_3226)
);

AO32x1_ASAP7_75t_L g3227 ( 
.A1(n_2627),
.A2(n_322),
.A3(n_320),
.B1(n_321),
.B2(n_323),
.Y(n_3227)
);

OAI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_2487),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2563),
.A2(n_321),
.B(n_322),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2631),
.Y(n_3230)
);

AOI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_2586),
.A2(n_323),
.B(n_324),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2631),
.Y(n_3232)
);

BUFx6f_ASAP7_75t_L g3233 ( 
.A(n_2622),
.Y(n_3233)
);

AO21x1_ASAP7_75t_L g3234 ( 
.A1(n_2767),
.A2(n_738),
.B(n_737),
.Y(n_3234)
);

OAI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_2595),
.A2(n_2754),
.B(n_2710),
.Y(n_3235)
);

AOI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_2566),
.A2(n_325),
.B(n_327),
.Y(n_3236)
);

NOR2x1_ASAP7_75t_L g3237 ( 
.A(n_2411),
.B(n_328),
.Y(n_3237)
);

NOR3xp33_ASAP7_75t_L g3238 ( 
.A(n_2403),
.B(n_328),
.C(n_329),
.Y(n_3238)
);

BUFx2_ASAP7_75t_L g3239 ( 
.A(n_2585),
.Y(n_3239)
);

AOI21xp5_ASAP7_75t_L g3240 ( 
.A1(n_2620),
.A2(n_328),
.B(n_329),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_2517),
.B(n_329),
.Y(n_3241)
);

NOR2xp33_ASAP7_75t_L g3242 ( 
.A(n_3088),
.B(n_2400),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2948),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2820),
.A2(n_2686),
.B(n_2674),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2887),
.Y(n_3245)
);

OAI22xp5_ASAP7_75t_L g3246 ( 
.A1(n_2866),
.A2(n_2674),
.B1(n_2725),
.B2(n_2686),
.Y(n_3246)
);

AND2x2_ASAP7_75t_L g3247 ( 
.A(n_2809),
.B(n_2725),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2966),
.Y(n_3248)
);

OAI21x1_ASAP7_75t_L g3249 ( 
.A1(n_3014),
.A2(n_2835),
.B(n_3078),
.Y(n_3249)
);

INVx3_ASAP7_75t_L g3250 ( 
.A(n_2828),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2880),
.B(n_2467),
.Y(n_3251)
);

AOI21x1_ASAP7_75t_L g3252 ( 
.A1(n_3201),
.A2(n_2735),
.B(n_2731),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3030),
.B(n_2519),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2810),
.B(n_2524),
.Y(n_3254)
);

AOI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_3015),
.A2(n_2736),
.B(n_2735),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2840),
.B(n_2848),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_3104),
.A2(n_2743),
.B(n_2736),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2857),
.B(n_2524),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2858),
.B(n_2545),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_3219),
.B(n_2593),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_2860),
.B(n_2545),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2868),
.B(n_2583),
.Y(n_3262)
);

NOR2xp33_ASAP7_75t_L g3263 ( 
.A(n_3042),
.B(n_2417),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2897),
.Y(n_3264)
);

INVx5_ASAP7_75t_L g3265 ( 
.A(n_2865),
.Y(n_3265)
);

INVx6_ASAP7_75t_L g3266 ( 
.A(n_2822),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2891),
.B(n_2340),
.Y(n_3267)
);

INVx4_ASAP7_75t_L g3268 ( 
.A(n_2819),
.Y(n_3268)
);

INVxp67_ASAP7_75t_L g3269 ( 
.A(n_2881),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2907),
.B(n_2340),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_L g3271 ( 
.A(n_3183),
.B(n_3224),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3104),
.A2(n_2743),
.B(n_2731),
.Y(n_3272)
);

BUFx6f_ASAP7_75t_L g3273 ( 
.A(n_3118),
.Y(n_3273)
);

O2A1O1Ixp33_ASAP7_75t_L g3274 ( 
.A1(n_3116),
.A2(n_2326),
.B(n_2729),
.C(n_2719),
.Y(n_3274)
);

NOR3xp33_ASAP7_75t_SL g3275 ( 
.A(n_2971),
.B(n_2619),
.C(n_2508),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_2865),
.A2(n_2795),
.B1(n_2770),
.B2(n_2766),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_2917),
.Y(n_3277)
);

HB1xp67_ASAP7_75t_L g3278 ( 
.A(n_2986),
.Y(n_3278)
);

AND2x2_ASAP7_75t_L g3279 ( 
.A(n_2816),
.B(n_2766),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_3127),
.A2(n_3175),
.B(n_3099),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_3127),
.A2(n_2622),
.B(n_2380),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_3175),
.A2(n_2380),
.B(n_2624),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2904),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2911),
.B(n_2360),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2975),
.Y(n_3285)
);

BUFx6f_ASAP7_75t_L g3286 ( 
.A(n_3118),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2995),
.Y(n_3287)
);

CKINVDCx14_ASAP7_75t_R g3288 ( 
.A(n_2924),
.Y(n_3288)
);

OAI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_3159),
.A2(n_2799),
.B1(n_2808),
.B2(n_2805),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2914),
.B(n_2360),
.Y(n_3290)
);

O2A1O1Ixp5_ASAP7_75t_L g3291 ( 
.A1(n_3235),
.A2(n_2605),
.B(n_2601),
.C(n_2317),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_2877),
.A2(n_2761),
.B(n_2621),
.Y(n_3292)
);

HB1xp67_ASAP7_75t_L g3293 ( 
.A(n_3239),
.Y(n_3293)
);

OAI22xp5_ASAP7_75t_L g3294 ( 
.A1(n_3159),
.A2(n_2805),
.B1(n_2808),
.B2(n_2799),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_2878),
.A2(n_2761),
.B(n_2317),
.Y(n_3295)
);

A2O1A1Ixp33_ASAP7_75t_L g3296 ( 
.A1(n_2836),
.A2(n_2521),
.B(n_2310),
.C(n_2427),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2942),
.B(n_2587),
.Y(n_3297)
);

INVx3_ASAP7_75t_L g3298 ( 
.A(n_2929),
.Y(n_3298)
);

AOI21x1_ASAP7_75t_L g3299 ( 
.A1(n_3190),
.A2(n_2521),
.B(n_2761),
.Y(n_3299)
);

AOI22xp33_ASAP7_75t_L g3300 ( 
.A1(n_3216),
.A2(n_2561),
.B1(n_2547),
.B2(n_2402),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_SL g3301 ( 
.A(n_3114),
.B(n_2372),
.Y(n_3301)
);

BUFx3_ASAP7_75t_L g3302 ( 
.A(n_3074),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2988),
.Y(n_3303)
);

NAND2x1p5_ASAP7_75t_L g3304 ( 
.A(n_2901),
.B(n_2618),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3019),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_3018),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_SL g3307 ( 
.A(n_2896),
.B(n_2613),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3029),
.Y(n_3308)
);

OAI22xp5_ASAP7_75t_L g3309 ( 
.A1(n_3188),
.A2(n_2515),
.B1(n_2562),
.B2(n_2498),
.Y(n_3309)
);

AOI221xp5_ASAP7_75t_L g3310 ( 
.A1(n_3146),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_3310)
);

INVx8_ASAP7_75t_L g3311 ( 
.A(n_2821),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3147),
.A2(n_2498),
.B1(n_2402),
.B2(n_333),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_2932),
.A2(n_2498),
.B(n_2402),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3040),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_2902),
.B(n_331),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3045),
.Y(n_3316)
);

A2O1A1Ixp33_ASAP7_75t_L g3317 ( 
.A1(n_3179),
.A2(n_333),
.B(n_331),
.C(n_332),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_3034),
.B(n_332),
.Y(n_3318)
);

O2A1O1Ixp33_ASAP7_75t_L g3319 ( 
.A1(n_2913),
.A2(n_337),
.B(n_335),
.C(n_336),
.Y(n_3319)
);

INVx6_ASAP7_75t_L g3320 ( 
.A(n_3180),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3035),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3043),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_2951),
.A2(n_336),
.B(n_337),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3068),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3126),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3144),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3150),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3048),
.Y(n_3328)
);

AOI21xp5_ASAP7_75t_L g3329 ( 
.A1(n_3169),
.A2(n_3033),
.B(n_3025),
.Y(n_3329)
);

OAI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_2997),
.A2(n_338),
.B(n_339),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_SL g3331 ( 
.A(n_3002),
.B(n_338),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3077),
.Y(n_3332)
);

BUFx3_ASAP7_75t_L g3333 ( 
.A(n_3186),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_2893),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3119),
.A2(n_340),
.B(n_341),
.Y(n_3335)
);

BUFx2_ASAP7_75t_L g3336 ( 
.A(n_2947),
.Y(n_3336)
);

INVx1_ASAP7_75t_SL g3337 ( 
.A(n_2817),
.Y(n_3337)
);

BUFx6f_ASAP7_75t_L g3338 ( 
.A(n_3118),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_SL g3339 ( 
.A(n_2852),
.B(n_342),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_2870),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_2954),
.B(n_343),
.Y(n_3341)
);

BUFx8_ASAP7_75t_L g3342 ( 
.A(n_2885),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_2889),
.B(n_3049),
.Y(n_3343)
);

BUFx6f_ASAP7_75t_L g3344 ( 
.A(n_3133),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_SL g3345 ( 
.A(n_2889),
.B(n_344),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_3223),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_3346)
);

AND2x6_ASAP7_75t_L g3347 ( 
.A(n_3194),
.B(n_345),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3000),
.B(n_346),
.Y(n_3348)
);

INVxp67_ASAP7_75t_SL g3349 ( 
.A(n_3205),
.Y(n_3349)
);

AOI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_2991),
.A2(n_3044),
.B(n_3171),
.Y(n_3350)
);

AOI21xp5_ASAP7_75t_L g3351 ( 
.A1(n_3187),
.A2(n_346),
.B(n_347),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3009),
.B(n_347),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_2906),
.Y(n_3353)
);

AO32x1_ASAP7_75t_L g3354 ( 
.A1(n_3221),
.A2(n_350),
.A3(n_348),
.B1(n_349),
.B2(n_351),
.Y(n_3354)
);

OAI22x1_ASAP7_75t_L g3355 ( 
.A1(n_2972),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3020),
.B(n_348),
.Y(n_3356)
);

O2A1O1Ixp33_ASAP7_75t_L g3357 ( 
.A1(n_2850),
.A2(n_351),
.B(n_349),
.C(n_350),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3062),
.B(n_352),
.Y(n_3358)
);

O2A1O1Ixp5_ASAP7_75t_L g3359 ( 
.A1(n_2813),
.A2(n_354),
.B(n_352),
.C(n_353),
.Y(n_3359)
);

AOI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_3039),
.A2(n_353),
.B(n_354),
.Y(n_3360)
);

A2O1A1Ixp33_ASAP7_75t_L g3361 ( 
.A1(n_2839),
.A2(n_357),
.B(n_355),
.C(n_356),
.Y(n_3361)
);

AOI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_3058),
.A2(n_355),
.B(n_356),
.Y(n_3362)
);

A2O1A1Ixp33_ASAP7_75t_L g3363 ( 
.A1(n_2990),
.A2(n_358),
.B(n_355),
.C(n_357),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3069),
.B(n_359),
.Y(n_3364)
);

AOI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_3209),
.A2(n_359),
.B(n_360),
.Y(n_3365)
);

O2A1O1Ixp5_ASAP7_75t_L g3366 ( 
.A1(n_3124),
.A2(n_361),
.B(n_359),
.C(n_360),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_SL g3367 ( 
.A(n_3111),
.B(n_361),
.Y(n_3367)
);

NOR3xp33_ASAP7_75t_L g3368 ( 
.A(n_3153),
.B(n_362),
.C(n_363),
.Y(n_3368)
);

BUFx6f_ASAP7_75t_L g3369 ( 
.A(n_3133),
.Y(n_3369)
);

O2A1O1Ixp33_ASAP7_75t_L g3370 ( 
.A1(n_2855),
.A2(n_366),
.B(n_364),
.C(n_365),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3075),
.B(n_364),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3079),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3115),
.B(n_366),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3149),
.B(n_367),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3134),
.B(n_368),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_2998),
.B(n_369),
.Y(n_3376)
);

AOI21x1_ASAP7_75t_L g3377 ( 
.A1(n_2812),
.A2(n_739),
.B(n_738),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_2909),
.B(n_371),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3092),
.Y(n_3379)
);

OAI21xp33_ASAP7_75t_L g3380 ( 
.A1(n_2968),
.A2(n_373),
.B(n_375),
.Y(n_3380)
);

INVx2_ASAP7_75t_L g3381 ( 
.A(n_2936),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3142),
.B(n_373),
.Y(n_3382)
);

INVx3_ASAP7_75t_L g3383 ( 
.A(n_3076),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3129),
.B(n_375),
.Y(n_3384)
);

O2A1O1Ixp33_ASAP7_75t_L g3385 ( 
.A1(n_2958),
.A2(n_378),
.B(n_376),
.C(n_377),
.Y(n_3385)
);

OAI21x1_ASAP7_75t_L g3386 ( 
.A1(n_2894),
.A2(n_379),
.B(n_377),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3157),
.Y(n_3387)
);

HB1xp67_ASAP7_75t_L g3388 ( 
.A(n_3054),
.Y(n_3388)
);

AOI21xp5_ASAP7_75t_L g3389 ( 
.A1(n_3181),
.A2(n_376),
.B(n_377),
.Y(n_3389)
);

BUFx2_ASAP7_75t_L g3390 ( 
.A(n_3133),
.Y(n_3390)
);

NOR2xp33_ASAP7_75t_L g3391 ( 
.A(n_2931),
.B(n_379),
.Y(n_3391)
);

NOR2xp33_ASAP7_75t_L g3392 ( 
.A(n_2862),
.B(n_379),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3166),
.Y(n_3393)
);

OAI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_2974),
.A2(n_380),
.B(n_382),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_2919),
.B(n_382),
.Y(n_3395)
);

NAND2x1p5_ASAP7_75t_L g3396 ( 
.A(n_3199),
.B(n_383),
.Y(n_3396)
);

A2O1A1Ixp33_ASAP7_75t_L g3397 ( 
.A1(n_2996),
.A2(n_385),
.B(n_383),
.C(n_384),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3003),
.B(n_383),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3007),
.B(n_384),
.Y(n_3399)
);

AO32x2_ASAP7_75t_L g3400 ( 
.A1(n_3184),
.A2(n_3228),
.A3(n_3177),
.B1(n_3148),
.B2(n_3082),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_2982),
.Y(n_3401)
);

AND2x4_ASAP7_75t_L g3402 ( 
.A(n_2823),
.B(n_2916),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_2869),
.A2(n_385),
.B(n_386),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_3167),
.B(n_386),
.Y(n_3404)
);

AOI21xp5_ASAP7_75t_L g3405 ( 
.A1(n_2934),
.A2(n_386),
.B(n_387),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3161),
.Y(n_3406)
);

AOI22xp33_ASAP7_75t_L g3407 ( 
.A1(n_2964),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_3407)
);

O2A1O1Ixp33_ASAP7_75t_L g3408 ( 
.A1(n_2935),
.A2(n_389),
.B(n_387),
.C(n_388),
.Y(n_3408)
);

BUFx2_ASAP7_75t_L g3409 ( 
.A(n_3128),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_2981),
.B(n_388),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_SL g3411 ( 
.A(n_3008),
.B(n_390),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_SL g3412 ( 
.A(n_2824),
.B(n_3052),
.Y(n_3412)
);

AO21x1_ASAP7_75t_L g3413 ( 
.A1(n_3220),
.A2(n_3232),
.B(n_3230),
.Y(n_3413)
);

OAI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_3095),
.A2(n_390),
.B(n_391),
.Y(n_3414)
);

O2A1O1Ixp33_ASAP7_75t_L g3415 ( 
.A1(n_3093),
.A2(n_395),
.B(n_392),
.C(n_393),
.Y(n_3415)
);

CKINVDCx5p33_ASAP7_75t_R g3416 ( 
.A(n_3168),
.Y(n_3416)
);

INVxp67_ASAP7_75t_SL g3417 ( 
.A(n_2811),
.Y(n_3417)
);

AOI21xp5_ASAP7_75t_L g3418 ( 
.A1(n_2969),
.A2(n_396),
.B(n_397),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_2984),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3158),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3055),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_3421)
);

O2A1O1Ixp33_ASAP7_75t_L g3422 ( 
.A1(n_3098),
.A2(n_401),
.B(n_399),
.C(n_400),
.Y(n_3422)
);

AOI21xp5_ASAP7_75t_L g3423 ( 
.A1(n_3016),
.A2(n_3170),
.B(n_2834),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_2959),
.B(n_399),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_SL g3425 ( 
.A(n_3036),
.B(n_400),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_2967),
.B(n_401),
.Y(n_3426)
);

O2A1O1Ixp33_ASAP7_75t_L g3427 ( 
.A1(n_3113),
.A2(n_3120),
.B(n_3165),
.C(n_3226),
.Y(n_3427)
);

AOI21xp5_ASAP7_75t_L g3428 ( 
.A1(n_2928),
.A2(n_402),
.B(n_403),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_3233),
.B(n_402),
.Y(n_3429)
);

AND2x4_ASAP7_75t_L g3430 ( 
.A(n_2823),
.B(n_403),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_2973),
.A2(n_403),
.B(n_404),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_2937),
.Y(n_3432)
);

BUFx12f_ASAP7_75t_L g3433 ( 
.A(n_3010),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_3028),
.A2(n_404),
.B(n_405),
.Y(n_3434)
);

A2O1A1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_2941),
.A2(n_408),
.B(n_405),
.C(n_406),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3197),
.B(n_406),
.Y(n_3436)
);

AOI21x1_ASAP7_75t_L g3437 ( 
.A1(n_3067),
.A2(n_741),
.B(n_740),
.Y(n_3437)
);

OR2x2_ASAP7_75t_L g3438 ( 
.A(n_2915),
.B(n_406),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3218),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_2957),
.B(n_2859),
.Y(n_3440)
);

NOR2xp33_ASAP7_75t_R g3441 ( 
.A(n_3128),
.B(n_2905),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_2864),
.B(n_408),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3195),
.Y(n_3443)
);

CKINVDCx5p33_ASAP7_75t_R g3444 ( 
.A(n_3173),
.Y(n_3444)
);

OAI21xp33_ASAP7_75t_SL g3445 ( 
.A1(n_3213),
.A2(n_409),
.B(n_410),
.Y(n_3445)
);

INVx3_ASAP7_75t_L g3446 ( 
.A(n_2953),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_L g3447 ( 
.A(n_2956),
.B(n_409),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_2965),
.B(n_411),
.Y(n_3448)
);

AOI21xp5_ASAP7_75t_L g3449 ( 
.A1(n_3031),
.A2(n_411),
.B(n_412),
.Y(n_3449)
);

CKINVDCx16_ASAP7_75t_R g3450 ( 
.A(n_3107),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_3140),
.B(n_3065),
.Y(n_3451)
);

A2O1A1Ixp33_ASAP7_75t_L g3452 ( 
.A1(n_2854),
.A2(n_415),
.B(n_413),
.C(n_414),
.Y(n_3452)
);

O2A1O1Ixp33_ASAP7_75t_L g3453 ( 
.A1(n_3156),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_3453)
);

OR2x6_ASAP7_75t_SL g3454 ( 
.A(n_2983),
.B(n_416),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_2943),
.Y(n_3455)
);

OAI22xp5_ASAP7_75t_L g3456 ( 
.A1(n_3200),
.A2(n_418),
.B1(n_416),
.B2(n_417),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_2944),
.Y(n_3457)
);

OAI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_2976),
.A2(n_417),
.B(n_418),
.Y(n_3458)
);

AOI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_3072),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_3459)
);

OAI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_3191),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_2811),
.Y(n_3461)
);

A2O1A1Ixp33_ASAP7_75t_L g3462 ( 
.A1(n_2886),
.A2(n_3056),
.B(n_3063),
.C(n_3038),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_2884),
.B(n_2814),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_2979),
.Y(n_3464)
);

NOR2xp33_ASAP7_75t_L g3465 ( 
.A(n_3182),
.B(n_422),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2945),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_2965),
.B(n_422),
.Y(n_3467)
);

O2A1O1Ixp33_ASAP7_75t_L g3468 ( 
.A1(n_3070),
.A2(n_425),
.B(n_423),
.C(n_424),
.Y(n_3468)
);

CKINVDCx5p33_ASAP7_75t_R g3469 ( 
.A(n_3027),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_2946),
.Y(n_3470)
);

A2O1A1Ixp33_ASAP7_75t_SL g3471 ( 
.A1(n_3238),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_3471)
);

OAI21xp33_ASAP7_75t_SL g3472 ( 
.A1(n_3138),
.A2(n_427),
.B(n_428),
.Y(n_3472)
);

O2A1O1Ixp33_ASAP7_75t_L g3473 ( 
.A1(n_3087),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_SL g3474 ( 
.A(n_3233),
.B(n_429),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_2979),
.Y(n_3475)
);

INVx3_ASAP7_75t_L g3476 ( 
.A(n_3198),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_2826),
.B(n_430),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3005),
.Y(n_3478)
);

O2A1O1Ixp33_ASAP7_75t_L g3479 ( 
.A1(n_3178),
.A2(n_433),
.B(n_431),
.C(n_432),
.Y(n_3479)
);

AOI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_2876),
.A2(n_431),
.B(n_432),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3005),
.B(n_431),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_2827),
.B(n_432),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_2952),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_2833),
.B(n_2844),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_SL g3485 ( 
.A(n_3128),
.B(n_433),
.Y(n_3485)
);

OR2x6_ASAP7_75t_L g3486 ( 
.A(n_3123),
.B(n_433),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3137),
.A2(n_434),
.B(n_435),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3203),
.B(n_434),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_R g3489 ( 
.A(n_3085),
.B(n_434),
.Y(n_3489)
);

OAI21xp33_ASAP7_75t_L g3490 ( 
.A1(n_3051),
.A2(n_435),
.B(n_436),
.Y(n_3490)
);

OAI22xp5_ASAP7_75t_L g3491 ( 
.A1(n_3217),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3204),
.B(n_436),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3141),
.A2(n_437),
.B(n_438),
.Y(n_3493)
);

BUFx2_ASAP7_75t_L g3494 ( 
.A(n_3135),
.Y(n_3494)
);

INVx2_ASAP7_75t_L g3495 ( 
.A(n_3096),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3121),
.B(n_437),
.Y(n_3496)
);

BUFx8_ASAP7_75t_L g3497 ( 
.A(n_2837),
.Y(n_3497)
);

NOR3xp33_ASAP7_75t_SL g3498 ( 
.A(n_3084),
.B(n_439),
.C(n_440),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3105),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3122),
.B(n_440),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3105),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_SL g3502 ( 
.A(n_3105),
.B(n_2849),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3011),
.B(n_441),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_SL g3504 ( 
.A(n_3237),
.B(n_443),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3225),
.B(n_444),
.Y(n_3505)
);

AND2x4_ASAP7_75t_L g3506 ( 
.A(n_2940),
.B(n_445),
.Y(n_3506)
);

OAI22x1_ASAP7_75t_L g3507 ( 
.A1(n_2892),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_2895),
.Y(n_3508)
);

BUFx2_ASAP7_75t_L g3509 ( 
.A(n_3198),
.Y(n_3509)
);

AOI22xp5_ASAP7_75t_L g3510 ( 
.A1(n_2851),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_3510)
);

BUFx6f_ASAP7_75t_L g3511 ( 
.A(n_3211),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_2970),
.Y(n_3512)
);

BUFx6f_ASAP7_75t_L g3513 ( 
.A(n_3211),
.Y(n_3513)
);

AOI22xp5_ASAP7_75t_L g3514 ( 
.A1(n_3081),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_3514)
);

OA21x2_ASAP7_75t_L g3515 ( 
.A1(n_2955),
.A2(n_2962),
.B(n_3145),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_2838),
.A2(n_2829),
.B(n_2987),
.Y(n_3516)
);

INVx2_ASAP7_75t_SL g3517 ( 
.A(n_2837),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_2872),
.B(n_449),
.Y(n_3518)
);

AND2x4_ASAP7_75t_L g3519 ( 
.A(n_2977),
.B(n_450),
.Y(n_3519)
);

AOI21xp5_ASAP7_75t_L g3520 ( 
.A1(n_2999),
.A2(n_450),
.B(n_451),
.Y(n_3520)
);

AO22x1_ASAP7_75t_L g3521 ( 
.A1(n_2960),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_2922),
.B(n_452),
.Y(n_3522)
);

OR2x2_ASAP7_75t_L g3523 ( 
.A(n_2888),
.B(n_452),
.Y(n_3523)
);

OR2x6_ASAP7_75t_L g3524 ( 
.A(n_3229),
.B(n_453),
.Y(n_3524)
);

NOR2xp67_ASAP7_75t_L g3525 ( 
.A(n_3193),
.B(n_2963),
.Y(n_3525)
);

O2A1O1Ixp5_ASAP7_75t_L g3526 ( 
.A1(n_3024),
.A2(n_456),
.B(n_454),
.C(n_455),
.Y(n_3526)
);

AOI22xp5_ASAP7_75t_L g3527 ( 
.A1(n_3164),
.A2(n_458),
.B1(n_456),
.B2(n_457),
.Y(n_3527)
);

AOI22xp5_ASAP7_75t_L g3528 ( 
.A1(n_3152),
.A2(n_3059),
.B1(n_3102),
.B2(n_2978),
.Y(n_3528)
);

INVx3_ASAP7_75t_L g3529 ( 
.A(n_3071),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_2989),
.Y(n_3530)
);

A2O1A1Ixp33_ASAP7_75t_L g3531 ( 
.A1(n_2930),
.A2(n_460),
.B(n_458),
.C(n_459),
.Y(n_3531)
);

INVx3_ASAP7_75t_L g3532 ( 
.A(n_3071),
.Y(n_3532)
);

AND2x4_ASAP7_75t_L g3533 ( 
.A(n_3013),
.B(n_459),
.Y(n_3533)
);

OR2x2_ASAP7_75t_L g3534 ( 
.A(n_2898),
.B(n_459),
.Y(n_3534)
);

BUFx6f_ASAP7_75t_L g3535 ( 
.A(n_3013),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_2912),
.Y(n_3536)
);

OAI21xp5_ASAP7_75t_L g3537 ( 
.A1(n_3004),
.A2(n_461),
.B(n_462),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_2992),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_2847),
.B(n_462),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_SL g3540 ( 
.A(n_2846),
.B(n_462),
.Y(n_3540)
);

BUFx6f_ASAP7_75t_L g3541 ( 
.A(n_3108),
.Y(n_3541)
);

A2O1A1Ixp33_ASAP7_75t_L g3542 ( 
.A1(n_3206),
.A2(n_465),
.B(n_463),
.C(n_464),
.Y(n_3542)
);

O2A1O1Ixp33_ASAP7_75t_L g3543 ( 
.A1(n_3210),
.A2(n_466),
.B(n_463),
.C(n_464),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3017),
.Y(n_3544)
);

NOR2xp67_ASAP7_75t_L g3545 ( 
.A(n_3108),
.B(n_463),
.Y(n_3545)
);

OA21x2_ASAP7_75t_L g3546 ( 
.A1(n_2863),
.A2(n_464),
.B(n_466),
.Y(n_3546)
);

AOI22xp33_ASAP7_75t_L g3547 ( 
.A1(n_3185),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_3547)
);

A2O1A1Ixp33_ASAP7_75t_SL g3548 ( 
.A1(n_3136),
.A2(n_469),
.B(n_467),
.C(n_468),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_2918),
.B(n_469),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_SL g3550 ( 
.A(n_3234),
.B(n_470),
.Y(n_3550)
);

O2A1O1Ixp5_ASAP7_75t_L g3551 ( 
.A1(n_2818),
.A2(n_2874),
.B(n_3110),
.C(n_3097),
.Y(n_3551)
);

NOR2xp33_ASAP7_75t_L g3552 ( 
.A(n_3207),
.B(n_470),
.Y(n_3552)
);

O2A1O1Ixp33_ASAP7_75t_L g3553 ( 
.A1(n_3214),
.A2(n_472),
.B(n_470),
.C(n_471),
.Y(n_3553)
);

OAI22xp5_ASAP7_75t_L g3554 ( 
.A1(n_3222),
.A2(n_474),
.B1(n_472),
.B2(n_473),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3012),
.A2(n_472),
.B(n_473),
.Y(n_3555)
);

A2O1A1Ixp33_ASAP7_75t_L g3556 ( 
.A1(n_3236),
.A2(n_475),
.B(n_473),
.C(n_474),
.Y(n_3556)
);

O2A1O1Ixp33_ASAP7_75t_L g3557 ( 
.A1(n_2925),
.A2(n_478),
.B(n_476),
.C(n_477),
.Y(n_3557)
);

AOI21xp5_ASAP7_75t_L g3558 ( 
.A1(n_3021),
.A2(n_476),
.B(n_478),
.Y(n_3558)
);

AOI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3022),
.A2(n_479),
.B(n_480),
.Y(n_3559)
);

A2O1A1Ixp33_ASAP7_75t_L g3560 ( 
.A1(n_3086),
.A2(n_482),
.B(n_480),
.C(n_481),
.Y(n_3560)
);

BUFx5_ASAP7_75t_L g3561 ( 
.A(n_3212),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_2949),
.Y(n_3562)
);

O2A1O1Ixp33_ASAP7_75t_L g3563 ( 
.A1(n_3215),
.A2(n_483),
.B(n_481),
.C(n_482),
.Y(n_3563)
);

HB1xp67_ASAP7_75t_L g3564 ( 
.A(n_2900),
.Y(n_3564)
);

A2O1A1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_2825),
.A2(n_484),
.B(n_481),
.C(n_483),
.Y(n_3565)
);

BUFx12f_ASAP7_75t_L g3566 ( 
.A(n_3227),
.Y(n_3566)
);

O2A1O1Ixp33_ASAP7_75t_L g3567 ( 
.A1(n_3006),
.A2(n_487),
.B(n_485),
.C(n_486),
.Y(n_3567)
);

BUFx3_ASAP7_75t_L g3568 ( 
.A(n_3241),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3001),
.Y(n_3569)
);

BUFx3_ASAP7_75t_L g3570 ( 
.A(n_3154),
.Y(n_3570)
);

AOI21xp33_ASAP7_75t_L g3571 ( 
.A1(n_2927),
.A2(n_487),
.B(n_488),
.Y(n_3571)
);

OAI22xp5_ASAP7_75t_L g3572 ( 
.A1(n_2933),
.A2(n_491),
.B1(n_489),
.B2(n_490),
.Y(n_3572)
);

OAI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_2831),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_3573)
);

AOI22xp5_ASAP7_75t_L g3574 ( 
.A1(n_2843),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3026),
.B(n_494),
.Y(n_3575)
);

INVxp67_ASAP7_75t_L g3576 ( 
.A(n_3160),
.Y(n_3576)
);

AND2x4_ASAP7_75t_L g3577 ( 
.A(n_3192),
.B(n_495),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_3176),
.B(n_495),
.Y(n_3578)
);

AND2x6_ASAP7_75t_L g3579 ( 
.A(n_3083),
.B(n_496),
.Y(n_3579)
);

OR2x2_ASAP7_75t_L g3580 ( 
.A(n_3037),
.B(n_496),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_SL g3581 ( 
.A(n_2882),
.B(n_2923),
.Y(n_3581)
);

AO32x1_ASAP7_75t_L g3582 ( 
.A1(n_3227),
.A2(n_498),
.A3(n_496),
.B1(n_497),
.B2(n_499),
.Y(n_3582)
);

OR2x2_ASAP7_75t_L g3583 ( 
.A(n_3053),
.B(n_498),
.Y(n_3583)
);

A2O1A1Ixp33_ASAP7_75t_L g3584 ( 
.A1(n_3208),
.A2(n_500),
.B(n_498),
.C(n_499),
.Y(n_3584)
);

O2A1O1Ixp5_ASAP7_75t_SL g3585 ( 
.A1(n_3172),
.A2(n_3174),
.B(n_3163),
.C(n_3162),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_SL g3586 ( 
.A(n_3061),
.B(n_499),
.Y(n_3586)
);

A2O1A1Ixp33_ASAP7_75t_L g3587 ( 
.A1(n_3202),
.A2(n_502),
.B(n_500),
.C(n_501),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_3089),
.A2(n_501),
.B(n_502),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_R g3589 ( 
.A(n_3041),
.B(n_503),
.Y(n_3589)
);

CKINVDCx20_ASAP7_75t_R g3590 ( 
.A(n_3091),
.Y(n_3590)
);

BUFx4f_ASAP7_75t_L g3591 ( 
.A(n_3125),
.Y(n_3591)
);

AO21x2_ASAP7_75t_L g3592 ( 
.A1(n_3057),
.A2(n_503),
.B(n_504),
.Y(n_3592)
);

OAI22xp5_ASAP7_75t_L g3593 ( 
.A1(n_2961),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3064),
.B(n_504),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_3090),
.A2(n_3131),
.B(n_3130),
.Y(n_3595)
);

A2O1A1Ixp33_ASAP7_75t_L g3596 ( 
.A1(n_3080),
.A2(n_507),
.B(n_505),
.C(n_506),
.Y(n_3596)
);

INVx3_ASAP7_75t_L g3597 ( 
.A(n_3094),
.Y(n_3597)
);

NAND3xp33_ASAP7_75t_SL g3598 ( 
.A(n_3231),
.B(n_2842),
.C(n_2867),
.Y(n_3598)
);

AOI22xp33_ASAP7_75t_L g3599 ( 
.A1(n_3151),
.A2(n_509),
.B1(n_505),
.B2(n_508),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_SL g3600 ( 
.A(n_2993),
.B(n_509),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3101),
.Y(n_3601)
);

AND2x4_ASAP7_75t_L g3602 ( 
.A(n_3109),
.B(n_510),
.Y(n_3602)
);

OAI22x1_ASAP7_75t_L g3603 ( 
.A1(n_3050),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_3603)
);

AOI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3196),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_2994),
.B(n_512),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3100),
.B(n_513),
.Y(n_3606)
);

AND2x2_ASAP7_75t_SL g3607 ( 
.A(n_3050),
.B(n_514),
.Y(n_3607)
);

AND2x2_ASAP7_75t_SL g3608 ( 
.A(n_3050),
.B(n_515),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_2871),
.A2(n_2832),
.B(n_2830),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_2861),
.A2(n_515),
.B(n_516),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3112),
.Y(n_3611)
);

BUFx3_ASAP7_75t_L g3612 ( 
.A(n_3060),
.Y(n_3612)
);

HB1xp67_ASAP7_75t_L g3613 ( 
.A(n_3189),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3132),
.B(n_516),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_L g3615 ( 
.A1(n_3240),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_3615)
);

NOR3xp33_ASAP7_75t_L g3616 ( 
.A(n_3139),
.B(n_3143),
.C(n_3106),
.Y(n_3616)
);

INVxp67_ASAP7_75t_L g3617 ( 
.A(n_3117),
.Y(n_3617)
);

NOR2xp33_ASAP7_75t_L g3618 ( 
.A(n_3155),
.B(n_3066),
.Y(n_3618)
);

A2O1A1Ixp33_ASAP7_75t_L g3619 ( 
.A1(n_3103),
.A2(n_522),
.B(n_520),
.C(n_521),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_3073),
.B(n_522),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_2845),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_2853),
.A2(n_2873),
.B(n_2856),
.Y(n_3622)
);

INVx4_ASAP7_75t_L g3623 ( 
.A(n_3023),
.Y(n_3623)
);

NAND2xp33_ASAP7_75t_SL g3624 ( 
.A(n_2875),
.B(n_526),
.Y(n_3624)
);

INVx2_ASAP7_75t_L g3625 ( 
.A(n_2879),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3032),
.B(n_526),
.Y(n_3626)
);

NOR2xp33_ASAP7_75t_R g3627 ( 
.A(n_2883),
.B(n_526),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_L g3628 ( 
.A(n_3046),
.B(n_527),
.Y(n_3628)
);

O2A1O1Ixp33_ASAP7_75t_L g3629 ( 
.A1(n_3047),
.A2(n_2910),
.B(n_2920),
.C(n_2908),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_2890),
.B(n_529),
.Y(n_3630)
);

A2O1A1Ixp33_ASAP7_75t_L g3631 ( 
.A1(n_2985),
.A2(n_531),
.B(n_529),
.C(n_530),
.Y(n_3631)
);

BUFx12f_ASAP7_75t_L g3632 ( 
.A(n_2899),
.Y(n_3632)
);

OAI21x1_ASAP7_75t_L g3633 ( 
.A1(n_2903),
.A2(n_531),
.B(n_530),
.Y(n_3633)
);

A2O1A1Ixp33_ASAP7_75t_L g3634 ( 
.A1(n_2921),
.A2(n_531),
.B(n_529),
.C(n_530),
.Y(n_3634)
);

AOI22xp33_ASAP7_75t_L g3635 ( 
.A1(n_2926),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.Y(n_3635)
);

NOR2xp33_ASAP7_75t_R g3636 ( 
.A(n_2938),
.B(n_532),
.Y(n_3636)
);

BUFx6f_ASAP7_75t_L g3637 ( 
.A(n_2939),
.Y(n_3637)
);

HB1xp67_ASAP7_75t_L g3638 ( 
.A(n_2950),
.Y(n_3638)
);

AOI22xp5_ASAP7_75t_L g3639 ( 
.A1(n_2980),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_3639)
);

BUFx2_ASAP7_75t_L g3640 ( 
.A(n_3180),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_2880),
.B(n_535),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_2880),
.B(n_535),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_2887),
.Y(n_3643)
);

A2O1A1Ixp33_ASAP7_75t_L g3644 ( 
.A1(n_2815),
.A2(n_539),
.B(n_537),
.C(n_538),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_2948),
.Y(n_3645)
);

OR2x6_ASAP7_75t_L g3646 ( 
.A(n_2828),
.B(n_539),
.Y(n_3646)
);

AOI21xp5_ASAP7_75t_L g3647 ( 
.A1(n_2820),
.A2(n_540),
.B(n_541),
.Y(n_3647)
);

AOI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_2820),
.A2(n_540),
.B(n_541),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_3118),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_SL g3650 ( 
.A(n_2866),
.B(n_542),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_2887),
.Y(n_3651)
);

OR2x6_ASAP7_75t_L g3652 ( 
.A(n_2828),
.B(n_542),
.Y(n_3652)
);

OAI21x1_ASAP7_75t_L g3653 ( 
.A1(n_3014),
.A2(n_545),
.B(n_544),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_SL g3654 ( 
.A(n_2866),
.B(n_543),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_SL g3655 ( 
.A(n_2866),
.B(n_543),
.Y(n_3655)
);

O2A1O1Ixp33_ASAP7_75t_L g3656 ( 
.A1(n_2841),
.A2(n_546),
.B(n_544),
.C(n_545),
.Y(n_3656)
);

BUFx6f_ASAP7_75t_L g3657 ( 
.A(n_3118),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_SL g3658 ( 
.A(n_2828),
.B(n_546),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_2809),
.B(n_546),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3379),
.Y(n_3660)
);

INVx3_ASAP7_75t_L g3661 ( 
.A(n_3266),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3243),
.B(n_547),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3387),
.Y(n_3663)
);

BUFx2_ASAP7_75t_SL g3664 ( 
.A(n_3265),
.Y(n_3664)
);

BUFx2_ASAP7_75t_SL g3665 ( 
.A(n_3265),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3420),
.Y(n_3666)
);

NOR2xp33_ASAP7_75t_L g3667 ( 
.A(n_3242),
.B(n_547),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3245),
.Y(n_3668)
);

INVx3_ASAP7_75t_L g3669 ( 
.A(n_3268),
.Y(n_3669)
);

INVx8_ASAP7_75t_L g3670 ( 
.A(n_3311),
.Y(n_3670)
);

INVx2_ASAP7_75t_SL g3671 ( 
.A(n_3320),
.Y(n_3671)
);

BUFx6f_ASAP7_75t_L g3672 ( 
.A(n_3511),
.Y(n_3672)
);

CKINVDCx11_ASAP7_75t_R g3673 ( 
.A(n_3311),
.Y(n_3673)
);

BUFx3_ASAP7_75t_L g3674 ( 
.A(n_3469),
.Y(n_3674)
);

INVx1_ASAP7_75t_SL g3675 ( 
.A(n_3444),
.Y(n_3675)
);

INVx3_ASAP7_75t_SL g3676 ( 
.A(n_3320),
.Y(n_3676)
);

BUFx6f_ASAP7_75t_L g3677 ( 
.A(n_3511),
.Y(n_3677)
);

BUFx12f_ASAP7_75t_L g3678 ( 
.A(n_3342),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3264),
.Y(n_3679)
);

BUFx6f_ASAP7_75t_L g3680 ( 
.A(n_3511),
.Y(n_3680)
);

INVx5_ASAP7_75t_L g3681 ( 
.A(n_3646),
.Y(n_3681)
);

CKINVDCx20_ASAP7_75t_R g3682 ( 
.A(n_3288),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3256),
.Y(n_3683)
);

AND2x4_ASAP7_75t_L g3684 ( 
.A(n_3640),
.B(n_549),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3441),
.Y(n_3685)
);

INVx4_ASAP7_75t_L g3686 ( 
.A(n_3302),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3283),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3247),
.B(n_548),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3287),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3306),
.Y(n_3690)
);

BUFx3_ASAP7_75t_L g3691 ( 
.A(n_3333),
.Y(n_3691)
);

BUFx12f_ASAP7_75t_L g3692 ( 
.A(n_3652),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3393),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3321),
.Y(n_3694)
);

BUFx6f_ASAP7_75t_L g3695 ( 
.A(n_3513),
.Y(n_3695)
);

INVx4_ASAP7_75t_L g3696 ( 
.A(n_3250),
.Y(n_3696)
);

BUFx2_ASAP7_75t_R g3697 ( 
.A(n_3416),
.Y(n_3697)
);

BUFx3_ASAP7_75t_L g3698 ( 
.A(n_3336),
.Y(n_3698)
);

BUFx3_ASAP7_75t_L g3699 ( 
.A(n_3277),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3643),
.Y(n_3700)
);

BUFx3_ASAP7_75t_L g3701 ( 
.A(n_3298),
.Y(n_3701)
);

INVx3_ASAP7_75t_L g3702 ( 
.A(n_3513),
.Y(n_3702)
);

BUFx6f_ASAP7_75t_L g3703 ( 
.A(n_3513),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3651),
.Y(n_3704)
);

INVx1_ASAP7_75t_SL g3705 ( 
.A(n_3337),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3406),
.Y(n_3706)
);

INVx5_ASAP7_75t_L g3707 ( 
.A(n_3450),
.Y(n_3707)
);

INVxp67_ASAP7_75t_SL g3708 ( 
.A(n_3278),
.Y(n_3708)
);

CKINVDCx20_ASAP7_75t_R g3709 ( 
.A(n_3497),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3322),
.Y(n_3710)
);

INVx6_ASAP7_75t_L g3711 ( 
.A(n_3433),
.Y(n_3711)
);

INVx1_ASAP7_75t_SL g3712 ( 
.A(n_3509),
.Y(n_3712)
);

INVx3_ASAP7_75t_L g3713 ( 
.A(n_3383),
.Y(n_3713)
);

INVx1_ASAP7_75t_SL g3714 ( 
.A(n_3293),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3324),
.B(n_551),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3325),
.Y(n_3716)
);

BUFx2_ASAP7_75t_L g3717 ( 
.A(n_3409),
.Y(n_3717)
);

BUFx12f_ASAP7_75t_L g3718 ( 
.A(n_3396),
.Y(n_3718)
);

INVx1_ASAP7_75t_SL g3719 ( 
.A(n_3446),
.Y(n_3719)
);

INVx6_ASAP7_75t_SL g3720 ( 
.A(n_3486),
.Y(n_3720)
);

INVx3_ASAP7_75t_SL g3721 ( 
.A(n_3506),
.Y(n_3721)
);

INVx1_ASAP7_75t_SL g3722 ( 
.A(n_3494),
.Y(n_3722)
);

NAND2x1p5_ASAP7_75t_L g3723 ( 
.A(n_3476),
.B(n_3430),
.Y(n_3723)
);

INVx1_ASAP7_75t_SL g3724 ( 
.A(n_3388),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3326),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3327),
.Y(n_3726)
);

BUFx3_ASAP7_75t_L g3727 ( 
.A(n_3304),
.Y(n_3727)
);

BUFx2_ASAP7_75t_L g3728 ( 
.A(n_3417),
.Y(n_3728)
);

CKINVDCx11_ASAP7_75t_R g3729 ( 
.A(n_3454),
.Y(n_3729)
);

NAND2x1p5_ASAP7_75t_L g3730 ( 
.A(n_3430),
.B(n_551),
.Y(n_3730)
);

INVx1_ASAP7_75t_SL g3731 ( 
.A(n_3448),
.Y(n_3731)
);

NAND2x1p5_ASAP7_75t_L g3732 ( 
.A(n_3519),
.B(n_553),
.Y(n_3732)
);

INVx4_ASAP7_75t_L g3733 ( 
.A(n_3529),
.Y(n_3733)
);

AND2x2_ASAP7_75t_SL g3734 ( 
.A(n_3485),
.B(n_554),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_SL g3735 ( 
.A(n_3246),
.B(n_554),
.Y(n_3735)
);

BUFx2_ASAP7_75t_L g3736 ( 
.A(n_3390),
.Y(n_3736)
);

NAND2x1p5_ASAP7_75t_L g3737 ( 
.A(n_3519),
.B(n_554),
.Y(n_3737)
);

BUFx4_ASAP7_75t_SL g3738 ( 
.A(n_3590),
.Y(n_3738)
);

BUFx2_ASAP7_75t_L g3739 ( 
.A(n_3273),
.Y(n_3739)
);

INVx5_ASAP7_75t_L g3740 ( 
.A(n_3286),
.Y(n_3740)
);

INVx3_ASAP7_75t_L g3741 ( 
.A(n_3402),
.Y(n_3741)
);

BUFx3_ASAP7_75t_L g3742 ( 
.A(n_3402),
.Y(n_3742)
);

INVx2_ASAP7_75t_SL g3743 ( 
.A(n_3561),
.Y(n_3743)
);

AOI22xp33_ASAP7_75t_L g3744 ( 
.A1(n_3591),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_3744)
);

AND2x2_ASAP7_75t_L g3745 ( 
.A(n_3340),
.B(n_555),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_3353),
.Y(n_3746)
);

INVx4_ASAP7_75t_L g3747 ( 
.A(n_3532),
.Y(n_3747)
);

BUFx3_ASAP7_75t_L g3748 ( 
.A(n_3517),
.Y(n_3748)
);

INVx2_ASAP7_75t_SL g3749 ( 
.A(n_3561),
.Y(n_3749)
);

INVxp67_ASAP7_75t_SL g3750 ( 
.A(n_3269),
.Y(n_3750)
);

INVx3_ASAP7_75t_L g3751 ( 
.A(n_3561),
.Y(n_3751)
);

BUFx2_ASAP7_75t_SL g3752 ( 
.A(n_3276),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3248),
.Y(n_3753)
);

BUFx2_ASAP7_75t_L g3754 ( 
.A(n_3286),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3285),
.Y(n_3755)
);

INVx1_ASAP7_75t_SL g3756 ( 
.A(n_3467),
.Y(n_3756)
);

BUFx5_ASAP7_75t_L g3757 ( 
.A(n_3632),
.Y(n_3757)
);

BUFx4f_ASAP7_75t_SL g3758 ( 
.A(n_3301),
.Y(n_3758)
);

BUFx6f_ASAP7_75t_L g3759 ( 
.A(n_3286),
.Y(n_3759)
);

CKINVDCx20_ASAP7_75t_R g3760 ( 
.A(n_3275),
.Y(n_3760)
);

BUFx3_ASAP7_75t_L g3761 ( 
.A(n_3533),
.Y(n_3761)
);

INVx2_ASAP7_75t_L g3762 ( 
.A(n_3381),
.Y(n_3762)
);

INVx3_ASAP7_75t_L g3763 ( 
.A(n_3535),
.Y(n_3763)
);

BUFx3_ASAP7_75t_L g3764 ( 
.A(n_3338),
.Y(n_3764)
);

CKINVDCx20_ASAP7_75t_R g3765 ( 
.A(n_3289),
.Y(n_3765)
);

INVx3_ASAP7_75t_L g3766 ( 
.A(n_3535),
.Y(n_3766)
);

INVx3_ASAP7_75t_L g3767 ( 
.A(n_3535),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3303),
.B(n_557),
.Y(n_3768)
);

BUFx3_ASAP7_75t_L g3769 ( 
.A(n_3338),
.Y(n_3769)
);

BUFx2_ASAP7_75t_L g3770 ( 
.A(n_3338),
.Y(n_3770)
);

BUFx2_ASAP7_75t_L g3771 ( 
.A(n_3344),
.Y(n_3771)
);

CKINVDCx11_ASAP7_75t_R g3772 ( 
.A(n_3294),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3401),
.Y(n_3773)
);

BUFx3_ASAP7_75t_L g3774 ( 
.A(n_3344),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3305),
.B(n_558),
.Y(n_3775)
);

BUFx3_ASAP7_75t_L g3776 ( 
.A(n_3344),
.Y(n_3776)
);

BUFx2_ASAP7_75t_L g3777 ( 
.A(n_3369),
.Y(n_3777)
);

INVx5_ASAP7_75t_L g3778 ( 
.A(n_3369),
.Y(n_3778)
);

AOI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_3313),
.A2(n_3502),
.B(n_3295),
.Y(n_3779)
);

BUFx12f_ASAP7_75t_L g3780 ( 
.A(n_3438),
.Y(n_3780)
);

BUFx3_ASAP7_75t_L g3781 ( 
.A(n_3369),
.Y(n_3781)
);

BUFx6f_ASAP7_75t_SL g3782 ( 
.A(n_3347),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3308),
.Y(n_3783)
);

OR2x2_ASAP7_75t_L g3784 ( 
.A(n_3251),
.B(n_558),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3314),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3316),
.Y(n_3786)
);

INVx4_ASAP7_75t_L g3787 ( 
.A(n_3649),
.Y(n_3787)
);

AOI22xp33_ASAP7_75t_SL g3788 ( 
.A1(n_3309),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3328),
.Y(n_3789)
);

INVxp67_ASAP7_75t_SL g3790 ( 
.A(n_3267),
.Y(n_3790)
);

CKINVDCx11_ASAP7_75t_R g3791 ( 
.A(n_3524),
.Y(n_3791)
);

INVx4_ASAP7_75t_L g3792 ( 
.A(n_3649),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3419),
.B(n_559),
.Y(n_3793)
);

INVx1_ASAP7_75t_SL g3794 ( 
.A(n_3378),
.Y(n_3794)
);

CKINVDCx20_ASAP7_75t_R g3795 ( 
.A(n_3424),
.Y(n_3795)
);

INVx5_ASAP7_75t_SL g3796 ( 
.A(n_3524),
.Y(n_3796)
);

INVx4_ASAP7_75t_L g3797 ( 
.A(n_3657),
.Y(n_3797)
);

AND2x4_ASAP7_75t_L g3798 ( 
.A(n_3279),
.B(n_562),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3332),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_3263),
.B(n_3260),
.Y(n_3800)
);

NAND2x1p5_ASAP7_75t_L g3801 ( 
.A(n_3282),
.B(n_561),
.Y(n_3801)
);

INVx1_ASAP7_75t_SL g3802 ( 
.A(n_3426),
.Y(n_3802)
);

BUFx3_ASAP7_75t_L g3803 ( 
.A(n_3657),
.Y(n_3803)
);

INVx5_ASAP7_75t_L g3804 ( 
.A(n_3541),
.Y(n_3804)
);

HB1xp67_ASAP7_75t_L g3805 ( 
.A(n_3372),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3318),
.B(n_562),
.Y(n_3806)
);

INVx4_ASAP7_75t_L g3807 ( 
.A(n_3579),
.Y(n_3807)
);

BUFx6f_ASAP7_75t_L g3808 ( 
.A(n_3461),
.Y(n_3808)
);

BUFx2_ASAP7_75t_SL g3809 ( 
.A(n_3545),
.Y(n_3809)
);

OAI22xp33_ASAP7_75t_SL g3810 ( 
.A1(n_3339),
.A2(n_3658),
.B1(n_3412),
.B2(n_3272),
.Y(n_3810)
);

NAND2x1p5_ASAP7_75t_L g3811 ( 
.A(n_3425),
.B(n_563),
.Y(n_3811)
);

BUFx8_ASAP7_75t_L g3812 ( 
.A(n_3503),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3645),
.B(n_564),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3564),
.B(n_565),
.Y(n_3814)
);

BUFx3_ASAP7_75t_L g3815 ( 
.A(n_3297),
.Y(n_3815)
);

BUFx2_ASAP7_75t_R g3816 ( 
.A(n_3650),
.Y(n_3816)
);

INVx4_ASAP7_75t_L g3817 ( 
.A(n_3579),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3262),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3432),
.B(n_565),
.Y(n_3819)
);

INVx3_ASAP7_75t_L g3820 ( 
.A(n_3570),
.Y(n_3820)
);

INVx4_ASAP7_75t_L g3821 ( 
.A(n_3579),
.Y(n_3821)
);

OR2x6_ASAP7_75t_L g3822 ( 
.A(n_3257),
.B(n_566),
.Y(n_3822)
);

NAND2x1p5_ASAP7_75t_L g3823 ( 
.A(n_3654),
.B(n_566),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3270),
.Y(n_3824)
);

BUFx6f_ASAP7_75t_L g3825 ( 
.A(n_3464),
.Y(n_3825)
);

INVx4_ASAP7_75t_L g3826 ( 
.A(n_3579),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3284),
.Y(n_3827)
);

BUFx3_ASAP7_75t_L g3828 ( 
.A(n_3568),
.Y(n_3828)
);

INVx3_ASAP7_75t_L g3829 ( 
.A(n_3602),
.Y(n_3829)
);

CKINVDCx8_ASAP7_75t_R g3830 ( 
.A(n_3347),
.Y(n_3830)
);

BUFx3_ASAP7_75t_L g3831 ( 
.A(n_3258),
.Y(n_3831)
);

BUFx6f_ASAP7_75t_L g3832 ( 
.A(n_3475),
.Y(n_3832)
);

INVx1_ASAP7_75t_SL g3833 ( 
.A(n_3259),
.Y(n_3833)
);

BUFx6f_ASAP7_75t_SL g3834 ( 
.A(n_3347),
.Y(n_3834)
);

NAND2x1p5_ASAP7_75t_L g3835 ( 
.A(n_3655),
.B(n_567),
.Y(n_3835)
);

BUFx2_ASAP7_75t_L g3836 ( 
.A(n_3443),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3290),
.Y(n_3837)
);

OAI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3300),
.A2(n_3498),
.B1(n_3254),
.B2(n_3334),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3455),
.B(n_3457),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3261),
.Y(n_3840)
);

BUFx8_ASAP7_75t_SL g3841 ( 
.A(n_3374),
.Y(n_3841)
);

AND2x2_ASAP7_75t_L g3842 ( 
.A(n_3659),
.B(n_567),
.Y(n_3842)
);

INVx4_ASAP7_75t_L g3843 ( 
.A(n_3549),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3341),
.Y(n_3844)
);

INVx5_ASAP7_75t_L g3845 ( 
.A(n_3597),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3437),
.Y(n_3846)
);

INVx6_ASAP7_75t_L g3847 ( 
.A(n_3577),
.Y(n_3847)
);

HB1xp67_ASAP7_75t_L g3848 ( 
.A(n_3349),
.Y(n_3848)
);

BUFx3_ASAP7_75t_L g3849 ( 
.A(n_3478),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3377),
.Y(n_3850)
);

INVx3_ASAP7_75t_L g3851 ( 
.A(n_3602),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3466),
.B(n_568),
.Y(n_3852)
);

INVx3_ASAP7_75t_L g3853 ( 
.A(n_3299),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3348),
.Y(n_3854)
);

BUFx8_ASAP7_75t_SL g3855 ( 
.A(n_3253),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3607),
.B(n_568),
.Y(n_3856)
);

BUFx3_ASAP7_75t_L g3857 ( 
.A(n_3495),
.Y(n_3857)
);

INVx3_ASAP7_75t_L g3858 ( 
.A(n_3523),
.Y(n_3858)
);

INVx2_ASAP7_75t_SL g3859 ( 
.A(n_3355),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3470),
.B(n_569),
.Y(n_3860)
);

CKINVDCx16_ASAP7_75t_R g3861 ( 
.A(n_3489),
.Y(n_3861)
);

AOI22xp5_ASAP7_75t_L g3862 ( 
.A1(n_3307),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_3862)
);

NAND2x1p5_ASAP7_75t_L g3863 ( 
.A(n_3411),
.B(n_572),
.Y(n_3863)
);

INVx1_ASAP7_75t_SL g3864 ( 
.A(n_3534),
.Y(n_3864)
);

INVx3_ASAP7_75t_L g3865 ( 
.A(n_3252),
.Y(n_3865)
);

CKINVDCx14_ASAP7_75t_R g3866 ( 
.A(n_3376),
.Y(n_3866)
);

INVx3_ASAP7_75t_SL g3867 ( 
.A(n_3343),
.Y(n_3867)
);

INVx3_ASAP7_75t_L g3868 ( 
.A(n_3499),
.Y(n_3868)
);

CKINVDCx20_ASAP7_75t_R g3869 ( 
.A(n_3451),
.Y(n_3869)
);

BUFx3_ASAP7_75t_L g3870 ( 
.A(n_3501),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3352),
.Y(n_3871)
);

BUFx3_ASAP7_75t_L g3872 ( 
.A(n_3391),
.Y(n_3872)
);

BUFx2_ASAP7_75t_L g3873 ( 
.A(n_3566),
.Y(n_3873)
);

BUFx12f_ASAP7_75t_L g3874 ( 
.A(n_3623),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3386),
.Y(n_3875)
);

BUFx2_ASAP7_75t_SL g3876 ( 
.A(n_3525),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3483),
.B(n_572),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3356),
.Y(n_3878)
);

INVx5_ASAP7_75t_L g3879 ( 
.A(n_3630),
.Y(n_3879)
);

BUFx6f_ASAP7_75t_L g3880 ( 
.A(n_3612),
.Y(n_3880)
);

INVx3_ASAP7_75t_L g3881 ( 
.A(n_3580),
.Y(n_3881)
);

BUFx3_ASAP7_75t_L g3882 ( 
.A(n_3447),
.Y(n_3882)
);

INVx3_ASAP7_75t_L g3883 ( 
.A(n_3583),
.Y(n_3883)
);

INVx1_ASAP7_75t_SL g3884 ( 
.A(n_3281),
.Y(n_3884)
);

OAI22xp5_ASAP7_75t_L g3885 ( 
.A1(n_3528),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.Y(n_3885)
);

INVx4_ASAP7_75t_L g3886 ( 
.A(n_3592),
.Y(n_3886)
);

BUFx12f_ASAP7_75t_L g3887 ( 
.A(n_3637),
.Y(n_3887)
);

AOI22xp33_ASAP7_75t_L g3888 ( 
.A1(n_3616),
.A2(n_575),
.B1(n_573),
.B2(n_574),
.Y(n_3888)
);

BUFx2_ASAP7_75t_L g3889 ( 
.A(n_3413),
.Y(n_3889)
);

INVxp67_ASAP7_75t_SL g3890 ( 
.A(n_3255),
.Y(n_3890)
);

INVx1_ASAP7_75t_SL g3891 ( 
.A(n_3540),
.Y(n_3891)
);

HB1xp67_ASAP7_75t_L g3892 ( 
.A(n_3440),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3512),
.Y(n_3893)
);

BUFx6f_ASAP7_75t_L g3894 ( 
.A(n_3637),
.Y(n_3894)
);

INVx2_ASAP7_75t_SL g3895 ( 
.A(n_3345),
.Y(n_3895)
);

BUFx3_ASAP7_75t_L g3896 ( 
.A(n_3410),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_L g3897 ( 
.A(n_3392),
.B(n_575),
.Y(n_3897)
);

BUFx3_ASAP7_75t_L g3898 ( 
.A(n_3522),
.Y(n_3898)
);

BUFx2_ASAP7_75t_R g3899 ( 
.A(n_3496),
.Y(n_3899)
);

BUFx12f_ASAP7_75t_L g3900 ( 
.A(n_3608),
.Y(n_3900)
);

INVx3_ASAP7_75t_L g3901 ( 
.A(n_3633),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3530),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3358),
.Y(n_3903)
);

BUFx3_ASAP7_75t_L g3904 ( 
.A(n_3641),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3538),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3364),
.Y(n_3906)
);

NAND2x1_ASAP7_75t_L g3907 ( 
.A(n_3508),
.B(n_576),
.Y(n_3907)
);

BUFx4_ASAP7_75t_SL g3908 ( 
.A(n_3544),
.Y(n_3908)
);

INVx1_ASAP7_75t_SL g3909 ( 
.A(n_3627),
.Y(n_3909)
);

INVx2_ASAP7_75t_SL g3910 ( 
.A(n_3507),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3601),
.Y(n_3911)
);

BUFx6f_ASAP7_75t_L g3912 ( 
.A(n_3429),
.Y(n_3912)
);

AND2x4_ASAP7_75t_L g3913 ( 
.A(n_3504),
.B(n_577),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3400),
.B(n_576),
.Y(n_3914)
);

AOI22xp5_ASAP7_75t_L g3915 ( 
.A1(n_3395),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.Y(n_3915)
);

BUFx6f_ASAP7_75t_L g3916 ( 
.A(n_3474),
.Y(n_3916)
);

BUFx3_ASAP7_75t_L g3917 ( 
.A(n_3642),
.Y(n_3917)
);

INVxp67_ASAP7_75t_SL g3918 ( 
.A(n_3244),
.Y(n_3918)
);

BUFx4f_ASAP7_75t_L g3919 ( 
.A(n_3546),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3371),
.Y(n_3920)
);

INVx2_ASAP7_75t_L g3921 ( 
.A(n_3546),
.Y(n_3921)
);

INVx2_ASAP7_75t_SL g3922 ( 
.A(n_3636),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3400),
.B(n_578),
.Y(n_3923)
);

BUFx2_ASAP7_75t_L g3924 ( 
.A(n_3638),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3373),
.Y(n_3925)
);

BUFx6f_ASAP7_75t_L g3926 ( 
.A(n_3271),
.Y(n_3926)
);

INVx4_ASAP7_75t_L g3927 ( 
.A(n_3515),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3400),
.B(n_3603),
.Y(n_3928)
);

AND2x4_ASAP7_75t_L g3929 ( 
.A(n_3296),
.B(n_580),
.Y(n_3929)
);

BUFx3_ASAP7_75t_L g3930 ( 
.A(n_3404),
.Y(n_3930)
);

BUFx3_ASAP7_75t_L g3931 ( 
.A(n_3518),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3375),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3653),
.Y(n_3933)
);

BUFx2_ASAP7_75t_L g3934 ( 
.A(n_3613),
.Y(n_3934)
);

BUFx3_ASAP7_75t_L g3935 ( 
.A(n_3384),
.Y(n_3935)
);

AOI22xp5_ASAP7_75t_L g3936 ( 
.A1(n_3380),
.A2(n_581),
.B1(n_578),
.B2(n_580),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3382),
.Y(n_3937)
);

INVx3_ASAP7_75t_L g3938 ( 
.A(n_3515),
.Y(n_3938)
);

INVxp67_ASAP7_75t_SL g3939 ( 
.A(n_3274),
.Y(n_3939)
);

BUFx2_ASAP7_75t_L g3940 ( 
.A(n_3445),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3576),
.B(n_581),
.Y(n_3941)
);

OR2x2_ASAP7_75t_L g3942 ( 
.A(n_3463),
.B(n_581),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3484),
.B(n_582),
.Y(n_3943)
);

INVx2_ASAP7_75t_SL g3944 ( 
.A(n_3481),
.Y(n_3944)
);

INVx4_ASAP7_75t_L g3945 ( 
.A(n_3439),
.Y(n_3945)
);

AND2x4_ASAP7_75t_L g3946 ( 
.A(n_3315),
.B(n_583),
.Y(n_3946)
);

INVx6_ASAP7_75t_L g3947 ( 
.A(n_3291),
.Y(n_3947)
);

INVx3_ASAP7_75t_L g3948 ( 
.A(n_3398),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_3611),
.B(n_582),
.Y(n_3949)
);

HB1xp67_ASAP7_75t_L g3950 ( 
.A(n_3617),
.Y(n_3950)
);

BUFx4f_ASAP7_75t_L g3951 ( 
.A(n_3521),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_3500),
.Y(n_3952)
);

BUFx2_ASAP7_75t_L g3953 ( 
.A(n_3472),
.Y(n_3953)
);

INVx1_ASAP7_75t_SL g3954 ( 
.A(n_3331),
.Y(n_3954)
);

BUFx3_ASAP7_75t_L g3955 ( 
.A(n_3465),
.Y(n_3955)
);

INVx8_ASAP7_75t_L g3956 ( 
.A(n_3368),
.Y(n_3956)
);

OR2x6_ASAP7_75t_L g3957 ( 
.A(n_3280),
.B(n_3312),
.Y(n_3957)
);

BUFx6f_ASAP7_75t_L g3958 ( 
.A(n_3626),
.Y(n_3958)
);

INVx4_ASAP7_75t_L g3959 ( 
.A(n_3625),
.Y(n_3959)
);

INVx2_ASAP7_75t_SL g3960 ( 
.A(n_3436),
.Y(n_3960)
);

NOR2xp33_ASAP7_75t_L g3961 ( 
.A(n_3552),
.B(n_582),
.Y(n_3961)
);

BUFx10_ASAP7_75t_L g3962 ( 
.A(n_3620),
.Y(n_3962)
);

HB1xp67_ASAP7_75t_L g3963 ( 
.A(n_3367),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3354),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3354),
.Y(n_3965)
);

BUFx2_ASAP7_75t_L g3966 ( 
.A(n_3249),
.Y(n_3966)
);

OR2x2_ASAP7_75t_L g3967 ( 
.A(n_3539),
.B(n_583),
.Y(n_3967)
);

AND2x2_ASAP7_75t_L g3968 ( 
.A(n_3536),
.B(n_584),
.Y(n_3968)
);

BUFx12f_ASAP7_75t_L g3969 ( 
.A(n_3589),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3595),
.B(n_584),
.Y(n_3970)
);

INVx5_ASAP7_75t_L g3971 ( 
.A(n_3562),
.Y(n_3971)
);

BUFx3_ASAP7_75t_L g3972 ( 
.A(n_3399),
.Y(n_3972)
);

INVx2_ASAP7_75t_SL g3973 ( 
.A(n_3572),
.Y(n_3973)
);

AND2x4_ASAP7_75t_L g3974 ( 
.A(n_3537),
.B(n_585),
.Y(n_3974)
);

INVxp67_ASAP7_75t_SL g3975 ( 
.A(n_3427),
.Y(n_3975)
);

INVxp67_ASAP7_75t_L g3976 ( 
.A(n_3442),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3578),
.Y(n_3977)
);

INVx4_ASAP7_75t_L g3978 ( 
.A(n_3569),
.Y(n_3978)
);

CKINVDCx5p33_ASAP7_75t_R g3979 ( 
.A(n_3514),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3575),
.Y(n_3980)
);

BUFx6f_ASAP7_75t_L g3981 ( 
.A(n_3505),
.Y(n_3981)
);

HB1xp67_ASAP7_75t_L g3982 ( 
.A(n_3621),
.Y(n_3982)
);

INVx1_ASAP7_75t_SL g3983 ( 
.A(n_3477),
.Y(n_3983)
);

BUFx6f_ASAP7_75t_L g3984 ( 
.A(n_3488),
.Y(n_3984)
);

BUFx5_ASAP7_75t_L g3985 ( 
.A(n_3624),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3421),
.B(n_586),
.Y(n_3986)
);

INVx2_ASAP7_75t_L g3987 ( 
.A(n_3526),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3582),
.Y(n_3988)
);

AOI22xp5_ASAP7_75t_L g3989 ( 
.A1(n_3573),
.A2(n_588),
.B1(n_586),
.B2(n_587),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_3366),
.Y(n_3990)
);

BUFx12f_ASAP7_75t_L g3991 ( 
.A(n_3527),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_L g3992 ( 
.A1(n_3581),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_3992)
);

BUFx3_ASAP7_75t_L g3993 ( 
.A(n_3482),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3594),
.Y(n_3994)
);

INVx3_ASAP7_75t_L g3995 ( 
.A(n_3606),
.Y(n_3995)
);

BUFx3_ASAP7_75t_L g3996 ( 
.A(n_3492),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3550),
.Y(n_3997)
);

CKINVDCx16_ASAP7_75t_R g3998 ( 
.A(n_3346),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3614),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3459),
.B(n_587),
.Y(n_4000)
);

CKINVDCx14_ASAP7_75t_R g4001 ( 
.A(n_3460),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3605),
.Y(n_4002)
);

NOR2xp33_ASAP7_75t_L g4003 ( 
.A(n_3571),
.B(n_588),
.Y(n_4003)
);

BUFx12f_ASAP7_75t_L g4004 ( 
.A(n_3548),
.Y(n_4004)
);

BUFx6f_ASAP7_75t_L g4005 ( 
.A(n_3618),
.Y(n_4005)
);

BUFx2_ASAP7_75t_L g4006 ( 
.A(n_3394),
.Y(n_4006)
);

INVx6_ASAP7_75t_L g4007 ( 
.A(n_3471),
.Y(n_4007)
);

BUFx2_ASAP7_75t_L g4008 ( 
.A(n_3458),
.Y(n_4008)
);

BUFx2_ASAP7_75t_L g4009 ( 
.A(n_3330),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3490),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3543),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3553),
.Y(n_4012)
);

OAI21x1_ASAP7_75t_L g4013 ( 
.A1(n_3938),
.A2(n_3779),
.B(n_3846),
.Y(n_4013)
);

AOI21xp33_ASAP7_75t_SL g4014 ( 
.A1(n_3670),
.A2(n_3456),
.B(n_3491),
.Y(n_4014)
);

OA21x2_ASAP7_75t_L g4015 ( 
.A1(n_3873),
.A2(n_3551),
.B(n_3329),
.Y(n_4015)
);

OAI21x1_ASAP7_75t_L g4016 ( 
.A1(n_3850),
.A2(n_3350),
.B(n_3292),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3794),
.B(n_589),
.Y(n_4017)
);

INVx2_ASAP7_75t_L g4018 ( 
.A(n_3668),
.Y(n_4018)
);

OAI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_4001),
.A2(n_3317),
.B1(n_3510),
.B2(n_3435),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3805),
.Y(n_4020)
);

INVx1_ASAP7_75t_SL g4021 ( 
.A(n_3908),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3679),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3660),
.Y(n_4023)
);

OAI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_3734),
.A2(n_3585),
.B(n_3361),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3892),
.B(n_3462),
.Y(n_4025)
);

OAI21x1_ASAP7_75t_L g4026 ( 
.A1(n_3865),
.A2(n_3622),
.B(n_3516),
.Y(n_4026)
);

AOI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3900),
.A2(n_3598),
.B1(n_3310),
.B2(n_3586),
.Y(n_4027)
);

OAI21x1_ASAP7_75t_L g4028 ( 
.A1(n_3853),
.A2(n_3901),
.B(n_3907),
.Y(n_4028)
);

AND2x4_ASAP7_75t_L g4029 ( 
.A(n_3685),
.B(n_3556),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3683),
.B(n_3423),
.Y(n_4030)
);

AOI22xp33_ASAP7_75t_L g4031 ( 
.A1(n_3991),
.A2(n_3628),
.B1(n_3600),
.B2(n_3554),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3663),
.Y(n_4032)
);

INVx4_ASAP7_75t_L g4033 ( 
.A(n_3673),
.Y(n_4033)
);

OAI21xp5_ASAP7_75t_L g4034 ( 
.A1(n_3951),
.A2(n_3397),
.B(n_3363),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3753),
.Y(n_4035)
);

OAI21x1_ASAP7_75t_L g4036 ( 
.A1(n_3907),
.A2(n_3609),
.B(n_3629),
.Y(n_4036)
);

NOR2xp67_ASAP7_75t_L g4037 ( 
.A(n_3681),
.B(n_3405),
.Y(n_4037)
);

AOI22xp5_ASAP7_75t_L g4038 ( 
.A1(n_3998),
.A2(n_3407),
.B1(n_3574),
.B2(n_3593),
.Y(n_4038)
);

OAI21x1_ASAP7_75t_L g4039 ( 
.A1(n_3921),
.A2(n_3933),
.B(n_3875),
.Y(n_4039)
);

NAND2x1p5_ASAP7_75t_L g4040 ( 
.A(n_3681),
.B(n_3604),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3687),
.Y(n_4041)
);

OAI21x1_ASAP7_75t_L g4042 ( 
.A1(n_3751),
.A2(n_3648),
.B(n_3647),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_4005),
.B(n_3414),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_3802),
.B(n_590),
.Y(n_4044)
);

BUFx2_ASAP7_75t_L g4045 ( 
.A(n_3685),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3755),
.Y(n_4046)
);

BUFx3_ASAP7_75t_L g4047 ( 
.A(n_3669),
.Y(n_4047)
);

CKINVDCx16_ASAP7_75t_R g4048 ( 
.A(n_3709),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3689),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3783),
.Y(n_4050)
);

OAI21x1_ASAP7_75t_SL g4051 ( 
.A1(n_3807),
.A2(n_3418),
.B(n_3656),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3785),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3818),
.B(n_3403),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3786),
.Y(n_4054)
);

NAND2x1p5_ASAP7_75t_L g4055 ( 
.A(n_3686),
.B(n_3639),
.Y(n_4055)
);

INVx2_ASAP7_75t_L g4056 ( 
.A(n_3690),
.Y(n_4056)
);

OR2x6_ASAP7_75t_L g4057 ( 
.A(n_3664),
.B(n_3665),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3789),
.Y(n_4058)
);

BUFx2_ASAP7_75t_L g4059 ( 
.A(n_3720),
.Y(n_4059)
);

AND2x4_ASAP7_75t_L g4060 ( 
.A(n_3817),
.B(n_3365),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3824),
.B(n_3588),
.Y(n_4061)
);

AND2x4_ASAP7_75t_L g4062 ( 
.A(n_3821),
.B(n_3644),
.Y(n_4062)
);

OA21x2_ASAP7_75t_L g4063 ( 
.A1(n_3873),
.A2(n_3359),
.B(n_3389),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3694),
.Y(n_4064)
);

OA21x2_ASAP7_75t_L g4065 ( 
.A1(n_3918),
.A2(n_3351),
.B(n_3323),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3827),
.B(n_3408),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3837),
.B(n_3335),
.Y(n_4067)
);

INVx2_ASAP7_75t_L g4068 ( 
.A(n_3700),
.Y(n_4068)
);

OAI21x1_ASAP7_75t_L g4069 ( 
.A1(n_3988),
.A2(n_3610),
.B(n_3362),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_3704),
.Y(n_4070)
);

BUFx2_ASAP7_75t_L g4071 ( 
.A(n_3672),
.Y(n_4071)
);

CKINVDCx20_ASAP7_75t_R g4072 ( 
.A(n_3682),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3799),
.B(n_3542),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_3746),
.Y(n_4074)
);

OAI21x1_ASAP7_75t_L g4075 ( 
.A1(n_3990),
.A2(n_3360),
.B(n_3480),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3693),
.Y(n_4076)
);

OR2x2_ASAP7_75t_L g4077 ( 
.A(n_3724),
.B(n_590),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3706),
.Y(n_4078)
);

OA21x2_ASAP7_75t_L g4079 ( 
.A1(n_3889),
.A2(n_3493),
.B(n_3487),
.Y(n_4079)
);

INVx8_ASAP7_75t_L g4080 ( 
.A(n_3678),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3893),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3902),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_3840),
.B(n_3531),
.Y(n_4083)
);

AND2x4_ASAP7_75t_L g4084 ( 
.A(n_3826),
.B(n_3596),
.Y(n_4084)
);

AOI221xp5_ASAP7_75t_L g4085 ( 
.A1(n_3897),
.A2(n_3319),
.B1(n_3557),
.B2(n_3479),
.C(n_3422),
.Y(n_4085)
);

OAI21x1_ASAP7_75t_SL g4086 ( 
.A1(n_3922),
.A2(n_3415),
.B(n_3453),
.Y(n_4086)
);

AO31x2_ASAP7_75t_L g4087 ( 
.A1(n_3889),
.A2(n_3886),
.A3(n_3966),
.B(n_3927),
.Y(n_4087)
);

OAI21x1_ASAP7_75t_L g4088 ( 
.A1(n_3977),
.A2(n_3431),
.B(n_3428),
.Y(n_4088)
);

AOI21xp5_ASAP7_75t_L g4089 ( 
.A1(n_3919),
.A2(n_3560),
.B(n_3473),
.Y(n_4089)
);

O2A1O1Ixp33_ASAP7_75t_SL g4090 ( 
.A1(n_3909),
.A2(n_3452),
.B(n_3565),
.C(n_3584),
.Y(n_4090)
);

CKINVDCx5p33_ASAP7_75t_R g4091 ( 
.A(n_3738),
.Y(n_4091)
);

NAND2x1p5_ASAP7_75t_L g4092 ( 
.A(n_3707),
.B(n_3434),
.Y(n_4092)
);

AO21x2_ASAP7_75t_L g4093 ( 
.A1(n_3975),
.A2(n_3449),
.B(n_3587),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3905),
.Y(n_4094)
);

OR2x2_ASAP7_75t_L g4095 ( 
.A(n_3708),
.B(n_591),
.Y(n_4095)
);

OAI22xp5_ASAP7_75t_L g4096 ( 
.A1(n_3861),
.A2(n_3547),
.B1(n_3635),
.B2(n_3615),
.Y(n_4096)
);

INVx4_ASAP7_75t_L g4097 ( 
.A(n_3696),
.Y(n_4097)
);

AOI21xp5_ASAP7_75t_L g4098 ( 
.A1(n_4006),
.A2(n_3468),
.B(n_3563),
.Y(n_4098)
);

BUFx2_ASAP7_75t_L g4099 ( 
.A(n_3672),
.Y(n_4099)
);

BUFx5_ASAP7_75t_L g4100 ( 
.A(n_3887),
.Y(n_4100)
);

NAND2x1p5_ASAP7_75t_L g4101 ( 
.A(n_3691),
.B(n_3520),
.Y(n_4101)
);

BUFx6f_ASAP7_75t_L g4102 ( 
.A(n_3677),
.Y(n_4102)
);

INVx4_ASAP7_75t_SL g4103 ( 
.A(n_3676),
.Y(n_4103)
);

AND2x4_ASAP7_75t_L g4104 ( 
.A(n_3828),
.B(n_3619),
.Y(n_4104)
);

OAI21x1_ASAP7_75t_L g4105 ( 
.A1(n_3997),
.A2(n_3702),
.B(n_3987),
.Y(n_4105)
);

OAI21x1_ASAP7_75t_L g4106 ( 
.A1(n_3723),
.A2(n_3558),
.B(n_3555),
.Y(n_4106)
);

OAI21x1_ASAP7_75t_SL g4107 ( 
.A1(n_3859),
.A2(n_3385),
.B(n_3370),
.Y(n_4107)
);

OAI21x1_ASAP7_75t_L g4108 ( 
.A1(n_3868),
.A2(n_3559),
.B(n_3567),
.Y(n_4108)
);

AOI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_4006),
.A2(n_3357),
.B(n_3631),
.Y(n_4109)
);

OA21x2_ASAP7_75t_L g4110 ( 
.A1(n_3890),
.A2(n_3634),
.B(n_3599),
.Y(n_4110)
);

AO31x2_ASAP7_75t_L g4111 ( 
.A1(n_3966),
.A2(n_593),
.A3(n_591),
.B(n_592),
.Y(n_4111)
);

NOR2x1_ASAP7_75t_R g4112 ( 
.A(n_3729),
.B(n_3692),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3911),
.Y(n_4113)
);

INVx2_ASAP7_75t_L g4114 ( 
.A(n_3762),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_3731),
.B(n_594),
.Y(n_4115)
);

AO31x2_ASAP7_75t_L g4116 ( 
.A1(n_3959),
.A2(n_3978),
.A3(n_3934),
.B(n_3924),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_3773),
.Y(n_4117)
);

AO21x2_ASAP7_75t_L g4118 ( 
.A1(n_3970),
.A2(n_595),
.B(n_596),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3848),
.Y(n_4119)
);

OA21x2_ASAP7_75t_L g4120 ( 
.A1(n_3939),
.A2(n_595),
.B(n_596),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3710),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3716),
.Y(n_4122)
);

OAI21x1_ASAP7_75t_L g4123 ( 
.A1(n_3763),
.A2(n_742),
.B(n_740),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3725),
.Y(n_4124)
);

OAI21x1_ASAP7_75t_L g4125 ( 
.A1(n_3766),
.A2(n_745),
.B(n_743),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3726),
.Y(n_4126)
);

OAI21x1_ASAP7_75t_L g4127 ( 
.A1(n_3767),
.A2(n_748),
.B(n_746),
.Y(n_4127)
);

AO31x2_ASAP7_75t_L g4128 ( 
.A1(n_3924),
.A2(n_599),
.A3(n_597),
.B(n_598),
.Y(n_4128)
);

AND2x2_ASAP7_75t_L g4129 ( 
.A(n_4005),
.B(n_599),
.Y(n_4129)
);

OR2x6_ASAP7_75t_L g4130 ( 
.A(n_3664),
.B(n_600),
.Y(n_4130)
);

OAI21x1_ASAP7_75t_L g4131 ( 
.A1(n_3950),
.A2(n_750),
.B(n_749),
.Y(n_4131)
);

AND2x4_ASAP7_75t_L g4132 ( 
.A(n_3698),
.B(n_600),
.Y(n_4132)
);

AOI21xp5_ASAP7_75t_L g4133 ( 
.A1(n_4008),
.A2(n_601),
.B(n_602),
.Y(n_4133)
);

OA21x2_ASAP7_75t_L g4134 ( 
.A1(n_4009),
.A2(n_602),
.B(n_603),
.Y(n_4134)
);

OAI21x1_ASAP7_75t_L g4135 ( 
.A1(n_3964),
.A2(n_751),
.B(n_750),
.Y(n_4135)
);

NAND2x1p5_ASAP7_75t_L g4136 ( 
.A(n_3699),
.B(n_603),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3750),
.Y(n_4137)
);

AO21x1_ASAP7_75t_L g4138 ( 
.A1(n_3810),
.A2(n_604),
.B(n_605),
.Y(n_4138)
);

OA21x2_ASAP7_75t_L g4139 ( 
.A1(n_4008),
.A2(n_3934),
.B(n_3965),
.Y(n_4139)
);

OAI21x1_ASAP7_75t_L g4140 ( 
.A1(n_3713),
.A2(n_753),
.B(n_752),
.Y(n_4140)
);

AND2x4_ASAP7_75t_SL g4141 ( 
.A(n_3820),
.B(n_604),
.Y(n_4141)
);

OAI21x1_ASAP7_75t_L g4142 ( 
.A1(n_3801),
.A2(n_3999),
.B(n_3995),
.Y(n_4142)
);

OAI21x1_ASAP7_75t_L g4143 ( 
.A1(n_3666),
.A2(n_754),
.B(n_753),
.Y(n_4143)
);

OAI222xp33_ASAP7_75t_L g4144 ( 
.A1(n_3822),
.A2(n_607),
.B1(n_609),
.B2(n_605),
.C1(n_606),
.C2(n_608),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3833),
.B(n_606),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3839),
.Y(n_4146)
);

AOI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_3957),
.A2(n_606),
.B(n_607),
.Y(n_4147)
);

OA21x2_ASAP7_75t_L g4148 ( 
.A1(n_3928),
.A2(n_607),
.B(n_608),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_3756),
.B(n_609),
.Y(n_4149)
);

OR2x2_ASAP7_75t_L g4150 ( 
.A(n_3714),
.B(n_609),
.Y(n_4150)
);

AO32x2_ASAP7_75t_L g4151 ( 
.A1(n_3910),
.A2(n_612),
.A3(n_610),
.B1(n_611),
.B2(n_613),
.Y(n_4151)
);

AO21x2_ASAP7_75t_L g4152 ( 
.A1(n_3914),
.A2(n_611),
.B(n_612),
.Y(n_4152)
);

OA21x2_ASAP7_75t_L g4153 ( 
.A1(n_3928),
.A2(n_612),
.B(n_613),
.Y(n_4153)
);

AO21x2_ASAP7_75t_L g4154 ( 
.A1(n_3914),
.A2(n_614),
.B(n_615),
.Y(n_4154)
);

OR2x2_ASAP7_75t_L g4155 ( 
.A(n_3722),
.B(n_615),
.Y(n_4155)
);

BUFx6f_ASAP7_75t_L g4156 ( 
.A(n_3677),
.Y(n_4156)
);

AO31x2_ASAP7_75t_L g4157 ( 
.A1(n_3945),
.A2(n_3754),
.A3(n_3770),
.B(n_3739),
.Y(n_4157)
);

OAI21x1_ASAP7_75t_L g4158 ( 
.A1(n_3982),
.A2(n_755),
.B(n_754),
.Y(n_4158)
);

AO31x2_ASAP7_75t_L g4159 ( 
.A1(n_3739),
.A2(n_618),
.A3(n_616),
.B(n_617),
.Y(n_4159)
);

OAI21x1_ASAP7_75t_L g4160 ( 
.A1(n_3829),
.A2(n_756),
.B(n_755),
.Y(n_4160)
);

NAND3xp33_ASAP7_75t_L g4161 ( 
.A(n_3923),
.B(n_619),
.C(n_620),
.Y(n_4161)
);

AO21x2_ASAP7_75t_L g4162 ( 
.A1(n_3923),
.A2(n_620),
.B(n_621),
.Y(n_4162)
);

AOI21xp5_ASAP7_75t_L g4163 ( 
.A1(n_3957),
.A2(n_621),
.B(n_622),
.Y(n_4163)
);

BUFx3_ASAP7_75t_L g4164 ( 
.A(n_3701),
.Y(n_4164)
);

OA21x2_ASAP7_75t_L g4165 ( 
.A1(n_3940),
.A2(n_622),
.B(n_623),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3790),
.B(n_624),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_3949),
.B(n_624),
.Y(n_4167)
);

HB1xp67_ASAP7_75t_L g4168 ( 
.A(n_3712),
.Y(n_4168)
);

OAI21x1_ASAP7_75t_L g4169 ( 
.A1(n_3851),
.A2(n_757),
.B(n_756),
.Y(n_4169)
);

OAI21x1_ASAP7_75t_L g4170 ( 
.A1(n_4010),
.A2(n_759),
.B(n_758),
.Y(n_4170)
);

OAI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_3796),
.A2(n_3830),
.B1(n_3765),
.B2(n_3879),
.Y(n_4171)
);

OR2x2_ASAP7_75t_L g4172 ( 
.A(n_3815),
.B(n_625),
.Y(n_4172)
);

OAI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_3879),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_4173)
);

OAI21xp33_ASAP7_75t_SL g4174 ( 
.A1(n_3822),
.A2(n_626),
.B(n_627),
.Y(n_4174)
);

INVx4_ASAP7_75t_L g4175 ( 
.A(n_3718),
.Y(n_4175)
);

AO21x2_ASAP7_75t_L g4176 ( 
.A1(n_3735),
.A2(n_628),
.B(n_629),
.Y(n_4176)
);

OR2x2_ASAP7_75t_L g4177 ( 
.A(n_3864),
.B(n_3688),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_3688),
.B(n_628),
.Y(n_4178)
);

OAI21x1_ASAP7_75t_L g4179 ( 
.A1(n_4011),
.A2(n_761),
.B(n_760),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3715),
.B(n_630),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_3849),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_3806),
.B(n_630),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_3857),
.Y(n_4183)
);

OAI21xp5_ASAP7_75t_L g4184 ( 
.A1(n_3788),
.A2(n_632),
.B(n_633),
.Y(n_4184)
);

OR2x6_ASAP7_75t_L g4185 ( 
.A(n_3665),
.B(n_632),
.Y(n_4185)
);

BUFx6f_ASAP7_75t_L g4186 ( 
.A(n_3680),
.Y(n_4186)
);

AO21x2_ASAP7_75t_L g4187 ( 
.A1(n_3814),
.A2(n_3968),
.B(n_3949),
.Y(n_4187)
);

OA21x2_ASAP7_75t_L g4188 ( 
.A1(n_3728),
.A2(n_633),
.B(n_634),
.Y(n_4188)
);

AOI22xp33_ASAP7_75t_L g4189 ( 
.A1(n_3782),
.A2(n_636),
.B1(n_634),
.B2(n_635),
.Y(n_4189)
);

OAI21x1_ASAP7_75t_L g4190 ( 
.A1(n_4012),
.A2(n_762),
.B(n_761),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_3870),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_3728),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3784),
.Y(n_4193)
);

INVx2_ASAP7_75t_SL g4194 ( 
.A(n_3674),
.Y(n_4194)
);

AOI22xp33_ASAP7_75t_L g4195 ( 
.A1(n_3834),
.A2(n_637),
.B1(n_635),
.B2(n_636),
.Y(n_4195)
);

OAI22xp33_ASAP7_75t_L g4196 ( 
.A1(n_3969),
.A2(n_638),
.B1(n_635),
.B2(n_637),
.Y(n_4196)
);

BUFx2_ASAP7_75t_L g4197 ( 
.A(n_3680),
.Y(n_4197)
);

OAI21xp5_ASAP7_75t_L g4198 ( 
.A1(n_3974),
.A2(n_639),
.B(n_640),
.Y(n_4198)
);

AO21x2_ASAP7_75t_L g4199 ( 
.A1(n_3936),
.A2(n_639),
.B(n_640),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3745),
.Y(n_4200)
);

OAI21x1_ASAP7_75t_L g4201 ( 
.A1(n_3963),
.A2(n_767),
.B(n_766),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_3745),
.Y(n_4202)
);

NAND2x1p5_ASAP7_75t_L g4203 ( 
.A(n_3727),
.B(n_641),
.Y(n_4203)
);

INVx2_ASAP7_75t_SL g4204 ( 
.A(n_3661),
.Y(n_4204)
);

AO21x2_ASAP7_75t_L g4205 ( 
.A1(n_3662),
.A2(n_643),
.B(n_644),
.Y(n_4205)
);

INVx4_ASAP7_75t_SL g4206 ( 
.A(n_3711),
.Y(n_4206)
);

AO21x2_ASAP7_75t_L g4207 ( 
.A1(n_3768),
.A2(n_644),
.B(n_645),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_3793),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3793),
.Y(n_4209)
);

BUFx2_ASAP7_75t_L g4210 ( 
.A(n_3695),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3876),
.Y(n_4211)
);

NAND2x1p5_ASAP7_75t_L g4212 ( 
.A(n_3671),
.B(n_645),
.Y(n_4212)
);

AO31x2_ASAP7_75t_L g4213 ( 
.A1(n_3754),
.A2(n_648),
.A3(n_646),
.B(n_647),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_3808),
.Y(n_4214)
);

NAND2x1p5_ASAP7_75t_L g4215 ( 
.A(n_3845),
.B(n_647),
.Y(n_4215)
);

OR2x6_ASAP7_75t_L g4216 ( 
.A(n_3752),
.B(n_648),
.Y(n_4216)
);

OAI21x1_ASAP7_75t_L g4217 ( 
.A1(n_4002),
.A2(n_769),
.B(n_766),
.Y(n_4217)
);

INVx2_ASAP7_75t_L g4218 ( 
.A(n_3808),
.Y(n_4218)
);

OAI21x1_ASAP7_75t_L g4219 ( 
.A1(n_3937),
.A2(n_3838),
.B(n_3741),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_3836),
.B(n_3856),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3825),
.Y(n_4221)
);

OAI21x1_ASAP7_75t_L g4222 ( 
.A1(n_3730),
.A2(n_770),
.B(n_769),
.Y(n_4222)
);

HB1xp67_ASAP7_75t_L g4223 ( 
.A(n_3736),
.Y(n_4223)
);

AOI22xp33_ASAP7_75t_L g4224 ( 
.A1(n_3953),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.Y(n_4224)
);

OR2x6_ASAP7_75t_L g4225 ( 
.A(n_3752),
.B(n_649),
.Y(n_4225)
);

O2A1O1Ixp33_ASAP7_75t_SL g4226 ( 
.A1(n_3795),
.A2(n_653),
.B(n_651),
.C(n_652),
.Y(n_4226)
);

OAI21x1_ASAP7_75t_L g4227 ( 
.A1(n_3732),
.A2(n_771),
.B(n_770),
.Y(n_4227)
);

OAI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_3929),
.A2(n_652),
.B(n_653),
.Y(n_4228)
);

OAI21x1_ASAP7_75t_L g4229 ( 
.A1(n_3737),
.A2(n_772),
.B(n_771),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3994),
.Y(n_4230)
);

INVx3_ASAP7_75t_L g4231 ( 
.A(n_3695),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_3825),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_3832),
.Y(n_4233)
);

NOR2xp33_ASAP7_75t_L g4234 ( 
.A(n_3855),
.B(n_654),
.Y(n_4234)
);

AND2x4_ASAP7_75t_L g4235 ( 
.A(n_3761),
.B(n_654),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_3844),
.B(n_654),
.Y(n_4236)
);

NOR2xp67_ASAP7_75t_SL g4237 ( 
.A(n_3809),
.B(n_655),
.Y(n_4237)
);

OAI21x1_ASAP7_75t_L g4238 ( 
.A1(n_3811),
.A2(n_775),
.B(n_774),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3854),
.B(n_655),
.Y(n_4239)
);

OR2x2_ASAP7_75t_L g4240 ( 
.A(n_3842),
.B(n_655),
.Y(n_4240)
);

OR2x6_ASAP7_75t_L g4241 ( 
.A(n_3847),
.B(n_656),
.Y(n_4241)
);

AND2x4_ASAP7_75t_L g4242 ( 
.A(n_3742),
.B(n_656),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_SL g4243 ( 
.A(n_3757),
.B(n_657),
.Y(n_4243)
);

HB1xp67_ASAP7_75t_L g4244 ( 
.A(n_3736),
.Y(n_4244)
);

BUFx3_ASAP7_75t_L g4245 ( 
.A(n_3703),
.Y(n_4245)
);

OAI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_3915),
.A2(n_658),
.B(n_659),
.Y(n_4246)
);

INVx8_ASAP7_75t_L g4247 ( 
.A(n_3841),
.Y(n_4247)
);

OA21x2_ASAP7_75t_L g4248 ( 
.A1(n_3717),
.A2(n_659),
.B(n_660),
.Y(n_4248)
);

CKINVDCx6p67_ASAP7_75t_R g4249 ( 
.A(n_3721),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4020),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_4116),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4023),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4032),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4116),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_4192),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4119),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4076),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4078),
.Y(n_4258)
);

AND2x4_ASAP7_75t_L g4259 ( 
.A(n_4057),
.B(n_3880),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4035),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4018),
.Y(n_4261)
);

BUFx3_ASAP7_75t_L g4262 ( 
.A(n_4164),
.Y(n_4262)
);

AOI22xp33_ASAP7_75t_L g4263 ( 
.A1(n_4019),
.A2(n_4004),
.B1(n_3872),
.B2(n_3896),
.Y(n_4263)
);

A2O1A1Ixp33_ASAP7_75t_L g4264 ( 
.A1(n_4174),
.A2(n_3956),
.B(n_3961),
.C(n_3684),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_4022),
.Y(n_4265)
);

INVx3_ASAP7_75t_L g4266 ( 
.A(n_4097),
.Y(n_4266)
);

BUFx12f_ASAP7_75t_L g4267 ( 
.A(n_4033),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4046),
.Y(n_4268)
);

HB1xp67_ASAP7_75t_L g4269 ( 
.A(n_4223),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_4041),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4049),
.Y(n_4271)
);

AND2x4_ASAP7_75t_L g4272 ( 
.A(n_4057),
.B(n_3880),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4056),
.Y(n_4273)
);

OR2x6_ASAP7_75t_L g4274 ( 
.A(n_4247),
.B(n_3874),
.Y(n_4274)
);

BUFx6f_ASAP7_75t_L g4275 ( 
.A(n_4047),
.Y(n_4275)
);

BUFx2_ASAP7_75t_L g4276 ( 
.A(n_4157),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4050),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_4064),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4052),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4054),
.Y(n_4280)
);

OR2x2_ASAP7_75t_L g4281 ( 
.A(n_4177),
.B(n_3705),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4058),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_4068),
.Y(n_4283)
);

INVx2_ASAP7_75t_L g4284 ( 
.A(n_4070),
.Y(n_4284)
);

BUFx6f_ASAP7_75t_L g4285 ( 
.A(n_4102),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_4074),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_4114),
.Y(n_4287)
);

AO21x2_ASAP7_75t_L g4288 ( 
.A1(n_4024),
.A2(n_3941),
.B(n_3852),
.Y(n_4288)
);

BUFx2_ASAP7_75t_L g4289 ( 
.A(n_4157),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4137),
.Y(n_4290)
);

BUFx3_ASAP7_75t_L g4291 ( 
.A(n_4080),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4117),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4081),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4082),
.Y(n_4294)
);

INVx3_ASAP7_75t_L g4295 ( 
.A(n_4249),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4094),
.Y(n_4296)
);

OAI21x1_ASAP7_75t_L g4297 ( 
.A1(n_4026),
.A2(n_3863),
.B(n_3835),
.Y(n_4297)
);

INVx2_ASAP7_75t_L g4298 ( 
.A(n_4113),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4230),
.Y(n_4299)
);

AO21x1_ASAP7_75t_SL g4300 ( 
.A1(n_4211),
.A2(n_3791),
.B(n_3757),
.Y(n_4300)
);

AND2x2_ASAP7_75t_L g4301 ( 
.A(n_4220),
.B(n_3926),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4121),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4122),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4124),
.Y(n_4304)
);

BUFx2_ASAP7_75t_SL g4305 ( 
.A(n_4100),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4126),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4146),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4168),
.Y(n_4308)
);

INVx4_ASAP7_75t_L g4309 ( 
.A(n_4103),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_L g4310 ( 
.A(n_4048),
.B(n_3866),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4045),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_4244),
.Y(n_4312)
);

OR2x6_ASAP7_75t_L g4313 ( 
.A(n_4216),
.B(n_3847),
.Y(n_4313)
);

BUFx6f_ASAP7_75t_L g4314 ( 
.A(n_4102),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4193),
.Y(n_4315)
);

AOI22xp33_ASAP7_75t_L g4316 ( 
.A1(n_4084),
.A2(n_3882),
.B1(n_4062),
.B2(n_4029),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_4187),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4030),
.Y(n_4318)
);

HB1xp67_ASAP7_75t_L g4319 ( 
.A(n_4181),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4025),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4183),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4200),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4202),
.Y(n_4323)
);

OAI21x1_ASAP7_75t_L g4324 ( 
.A1(n_4028),
.A2(n_3823),
.B(n_3881),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4208),
.Y(n_4325)
);

BUFx3_ASAP7_75t_L g4326 ( 
.A(n_4080),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_4191),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4139),
.Y(n_4328)
);

INVx1_ASAP7_75t_SL g4329 ( 
.A(n_4021),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4209),
.B(n_3926),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4095),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4214),
.Y(n_4332)
);

OAI21x1_ASAP7_75t_L g4333 ( 
.A1(n_4013),
.A2(n_3883),
.B(n_3858),
.Y(n_4333)
);

HB1xp67_ASAP7_75t_L g4334 ( 
.A(n_4129),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4218),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4077),
.Y(n_4336)
);

AOI22xp33_ASAP7_75t_L g4337 ( 
.A1(n_4225),
.A2(n_3955),
.B1(n_3930),
.B2(n_3956),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4221),
.Y(n_4338)
);

NOR2x1_ASAP7_75t_SL g4339 ( 
.A(n_4225),
.B(n_3743),
.Y(n_4339)
);

BUFx6f_ASAP7_75t_L g4340 ( 
.A(n_4156),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4232),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4150),
.Y(n_4342)
);

INVx2_ASAP7_75t_SL g4343 ( 
.A(n_4103),
.Y(n_4343)
);

BUFx6f_ASAP7_75t_L g4344 ( 
.A(n_4156),
.Y(n_4344)
);

AOI21x1_ASAP7_75t_L g4345 ( 
.A1(n_4037),
.A2(n_3771),
.B(n_3770),
.Y(n_4345)
);

OA21x2_ASAP7_75t_L g4346 ( 
.A1(n_4219),
.A2(n_3836),
.B(n_3777),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4233),
.Y(n_4347)
);

AOI22xp33_ASAP7_75t_SL g4348 ( 
.A1(n_4171),
.A2(n_3757),
.B1(n_3758),
.B2(n_3947),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4155),
.Y(n_4349)
);

AOI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_4085),
.A2(n_4007),
.B1(n_3898),
.B2(n_3772),
.Y(n_4350)
);

NOR2xp67_ASAP7_75t_L g4351 ( 
.A(n_4175),
.B(n_3780),
.Y(n_4351)
);

BUFx2_ASAP7_75t_L g4352 ( 
.A(n_4071),
.Y(n_4352)
);

OAI21x1_ASAP7_75t_L g4353 ( 
.A1(n_4036),
.A2(n_3888),
.B(n_3885),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4167),
.B(n_3980),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4099),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_4197),
.Y(n_4356)
);

CKINVDCx20_ASAP7_75t_R g4357 ( 
.A(n_4072),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_4210),
.Y(n_4358)
);

OAI21x1_ASAP7_75t_L g4359 ( 
.A1(n_4016),
.A2(n_3878),
.B(n_3871),
.Y(n_4359)
);

INVx3_ASAP7_75t_L g4360 ( 
.A(n_4130),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4053),
.Y(n_4361)
);

BUFx6f_ASAP7_75t_L g4362 ( 
.A(n_4186),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4167),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_4109),
.A2(n_3749),
.B(n_3771),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4039),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4105),
.Y(n_4366)
);

BUFx2_ASAP7_75t_L g4367 ( 
.A(n_4245),
.Y(n_4367)
);

OR2x6_ASAP7_75t_L g4368 ( 
.A(n_4130),
.B(n_3711),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4166),
.Y(n_4369)
);

AND2x2_ASAP7_75t_L g4370 ( 
.A(n_4182),
.B(n_3843),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4087),
.Y(n_4371)
);

INVx2_ASAP7_75t_SL g4372 ( 
.A(n_4091),
.Y(n_4372)
);

OAI21x1_ASAP7_75t_L g4373 ( 
.A1(n_4142),
.A2(n_3906),
.B(n_3903),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4061),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4087),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4165),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4043),
.Y(n_4377)
);

OAI21x1_ASAP7_75t_L g4378 ( 
.A1(n_4069),
.A2(n_3925),
.B(n_3920),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_4188),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4111),
.Y(n_4380)
);

NAND4xp25_ASAP7_75t_L g4381 ( 
.A(n_4264),
.B(n_4031),
.C(n_4027),
.D(n_4234),
.Y(n_4381)
);

BUFx6f_ASAP7_75t_L g4382 ( 
.A(n_4275),
.Y(n_4382)
);

NOR2x1p5_ASAP7_75t_L g4383 ( 
.A(n_4309),
.B(n_4240),
.Y(n_4383)
);

AND2x4_ASAP7_75t_L g4384 ( 
.A(n_4259),
.B(n_4206),
.Y(n_4384)
);

BUFx8_ASAP7_75t_L g4385 ( 
.A(n_4267),
.Y(n_4385)
);

NOR2xp33_ASAP7_75t_L g4386 ( 
.A(n_4329),
.B(n_4112),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4252),
.Y(n_4387)
);

CKINVDCx16_ASAP7_75t_R g4388 ( 
.A(n_4291),
.Y(n_4388)
);

CKINVDCx5p33_ASAP7_75t_R g4389 ( 
.A(n_4326),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_4352),
.Y(n_4390)
);

CKINVDCx5p33_ASAP7_75t_R g4391 ( 
.A(n_4357),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4301),
.B(n_4059),
.Y(n_4392)
);

OR2x6_ASAP7_75t_L g4393 ( 
.A(n_4274),
.B(n_4185),
.Y(n_4393)
);

CKINVDCx16_ASAP7_75t_R g4394 ( 
.A(n_4262),
.Y(n_4394)
);

HB1xp67_ASAP7_75t_L g4395 ( 
.A(n_4269),
.Y(n_4395)
);

BUFx3_ASAP7_75t_L g4396 ( 
.A(n_4275),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4253),
.Y(n_4397)
);

INVxp67_ASAP7_75t_L g4398 ( 
.A(n_4352),
.Y(n_4398)
);

AND2x2_ASAP7_75t_L g4399 ( 
.A(n_4377),
.B(n_4194),
.Y(n_4399)
);

BUFx6f_ASAP7_75t_L g4400 ( 
.A(n_4285),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4334),
.B(n_3719),
.Y(n_4401)
);

AO32x1_ASAP7_75t_L g4402 ( 
.A1(n_4343),
.A2(n_4173),
.A3(n_4141),
.B1(n_4204),
.B2(n_3960),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4257),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4258),
.Y(n_4404)
);

NOR2xp33_ASAP7_75t_R g4405 ( 
.A(n_4266),
.B(n_3760),
.Y(n_4405)
);

CKINVDCx5p33_ASAP7_75t_R g4406 ( 
.A(n_4295),
.Y(n_4406)
);

INVx3_ASAP7_75t_L g4407 ( 
.A(n_4368),
.Y(n_4407)
);

OR2x6_ASAP7_75t_L g4408 ( 
.A(n_4313),
.B(n_4305),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_4319),
.B(n_4311),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4260),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4261),
.Y(n_4411)
);

BUFx6f_ASAP7_75t_L g4412 ( 
.A(n_4285),
.Y(n_4412)
);

NOR2x1p5_ASAP7_75t_L g4413 ( 
.A(n_4360),
.B(n_4172),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4268),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_4308),
.B(n_4017),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4277),
.Y(n_4416)
);

AO31x2_ASAP7_75t_L g4417 ( 
.A1(n_4276),
.A2(n_4138),
.A3(n_3800),
.B(n_4145),
.Y(n_4417)
);

AO22x1_ASAP7_75t_L g4418 ( 
.A1(n_4259),
.A2(n_3812),
.B1(n_4132),
.B2(n_4198),
.Y(n_4418)
);

HB1xp67_ASAP7_75t_L g4419 ( 
.A(n_4312),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_L g4420 ( 
.A(n_4320),
.B(n_4152),
.Y(n_4420)
);

HB1xp67_ASAP7_75t_L g4421 ( 
.A(n_4255),
.Y(n_4421)
);

NOR3xp33_ASAP7_75t_SL g4422 ( 
.A(n_4310),
.B(n_4196),
.C(n_4144),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4279),
.Y(n_4423)
);

CKINVDCx20_ASAP7_75t_R g4424 ( 
.A(n_4372),
.Y(n_4424)
);

AND2x2_ASAP7_75t_L g4425 ( 
.A(n_4355),
.B(n_4044),
.Y(n_4425)
);

NOR2xp33_ASAP7_75t_R g4426 ( 
.A(n_4367),
.B(n_4100),
.Y(n_4426)
);

HB1xp67_ASAP7_75t_L g4427 ( 
.A(n_4367),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_4265),
.Y(n_4428)
);

OR2x2_ASAP7_75t_L g4429 ( 
.A(n_4363),
.B(n_4178),
.Y(n_4429)
);

BUFx6f_ASAP7_75t_L g4430 ( 
.A(n_4314),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_4318),
.B(n_4154),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4270),
.Y(n_4432)
);

AND2x2_ASAP7_75t_L g4433 ( 
.A(n_4356),
.B(n_4115),
.Y(n_4433)
);

AND2x2_ASAP7_75t_L g4434 ( 
.A(n_4358),
.B(n_4149),
.Y(n_4434)
);

NOR2xp33_ASAP7_75t_R g4435 ( 
.A(n_4370),
.B(n_4100),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4330),
.B(n_4015),
.Y(n_4436)
);

OAI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_4337),
.A2(n_4241),
.B1(n_4040),
.B2(n_3867),
.Y(n_4437)
);

OR2x2_ASAP7_75t_L g4438 ( 
.A(n_4361),
.B(n_3831),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4280),
.Y(n_4439)
);

OR2x6_ASAP7_75t_L g4440 ( 
.A(n_4272),
.B(n_4136),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_4374),
.B(n_4162),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_4281),
.B(n_4321),
.Y(n_4442)
);

INVx1_ASAP7_75t_L g4443 ( 
.A(n_4282),
.Y(n_4443)
);

NAND2xp33_ASAP7_75t_SL g4444 ( 
.A(n_4272),
.B(n_4237),
.Y(n_4444)
);

AOI22xp33_ASAP7_75t_SL g4445 ( 
.A1(n_4339),
.A2(n_4104),
.B1(n_4153),
.B2(n_4148),
.Y(n_4445)
);

OAI21xp5_ASAP7_75t_SL g4446 ( 
.A1(n_4348),
.A2(n_4215),
.B(n_4203),
.Y(n_4446)
);

NOR2xp33_ASAP7_75t_R g4447 ( 
.A(n_4300),
.B(n_4100),
.Y(n_4447)
);

CKINVDCx5p33_ASAP7_75t_R g4448 ( 
.A(n_4314),
.Y(n_4448)
);

AOI22xp33_ASAP7_75t_L g4449 ( 
.A1(n_4263),
.A2(n_4007),
.B1(n_4107),
.B2(n_4051),
.Y(n_4449)
);

NAND3xp33_ASAP7_75t_L g4450 ( 
.A(n_4317),
.B(n_4034),
.C(n_3976),
.Y(n_4450)
);

OAI22xp5_ASAP7_75t_L g4451 ( 
.A1(n_4316),
.A2(n_4055),
.B1(n_4161),
.B2(n_4101),
.Y(n_4451)
);

CKINVDCx5p33_ASAP7_75t_R g4452 ( 
.A(n_4340),
.Y(n_4452)
);

AND2x2_ASAP7_75t_L g4453 ( 
.A(n_4327),
.B(n_3971),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4306),
.Y(n_4454)
);

NOR2x1_ASAP7_75t_SL g4455 ( 
.A(n_4345),
.B(n_4243),
.Y(n_4455)
);

AND2x4_ASAP7_75t_L g4456 ( 
.A(n_4336),
.B(n_4206),
.Y(n_4456)
);

OAI21xp5_ASAP7_75t_L g4457 ( 
.A1(n_4364),
.A2(n_4163),
.B(n_4147),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4342),
.B(n_4060),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4349),
.B(n_3894),
.Y(n_4459)
);

NAND2xp33_ASAP7_75t_SL g4460 ( 
.A(n_4376),
.B(n_3869),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_4369),
.B(n_3983),
.Y(n_4461)
);

CKINVDCx5p33_ASAP7_75t_R g4462 ( 
.A(n_4340),
.Y(n_4462)
);

AND2x4_ASAP7_75t_L g4463 ( 
.A(n_4322),
.B(n_4231),
.Y(n_4463)
);

INVx8_ASAP7_75t_L g4464 ( 
.A(n_4344),
.Y(n_4464)
);

AO31x2_ASAP7_75t_L g4465 ( 
.A1(n_4276),
.A2(n_3777),
.A3(n_3667),
.B(n_4098),
.Y(n_4465)
);

NAND3xp33_ASAP7_75t_SL g4466 ( 
.A(n_4350),
.B(n_4228),
.C(n_4212),
.Y(n_4466)
);

OR2x2_ASAP7_75t_SL g4467 ( 
.A(n_4346),
.B(n_4248),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4302),
.Y(n_4468)
);

CKINVDCx5p33_ASAP7_75t_R g4469 ( 
.A(n_4344),
.Y(n_4469)
);

INVx2_ASAP7_75t_L g4470 ( 
.A(n_4271),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4250),
.B(n_4307),
.Y(n_4471)
);

NOR2xp33_ASAP7_75t_L g4472 ( 
.A(n_4331),
.B(n_3899),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4303),
.Y(n_4473)
);

AOI22xp33_ASAP7_75t_L g4474 ( 
.A1(n_4288),
.A2(n_3952),
.B1(n_3958),
.B2(n_4096),
.Y(n_4474)
);

AOI22xp33_ASAP7_75t_L g4475 ( 
.A1(n_4466),
.A2(n_4379),
.B1(n_3979),
.B2(n_3962),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4468),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_4427),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4473),
.Y(n_4478)
);

INVx3_ASAP7_75t_L g4479 ( 
.A(n_4408),
.Y(n_4479)
);

HB1xp67_ASAP7_75t_L g4480 ( 
.A(n_4395),
.Y(n_4480)
);

BUFx2_ASAP7_75t_L g4481 ( 
.A(n_4447),
.Y(n_4481)
);

INVx2_ASAP7_75t_L g4482 ( 
.A(n_4411),
.Y(n_4482)
);

INVx1_ASAP7_75t_SL g4483 ( 
.A(n_4394),
.Y(n_4483)
);

OR2x2_ASAP7_75t_L g4484 ( 
.A(n_4419),
.B(n_4421),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4436),
.B(n_4256),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4428),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4458),
.B(n_4315),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4442),
.B(n_4289),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4401),
.B(n_4289),
.Y(n_4489)
);

OR2x2_ASAP7_75t_L g4490 ( 
.A(n_4429),
.B(n_4290),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4390),
.B(n_4409),
.Y(n_4491)
);

NOR2xp33_ASAP7_75t_SL g4492 ( 
.A(n_4388),
.B(n_3697),
.Y(n_4492)
);

BUFx3_ASAP7_75t_L g4493 ( 
.A(n_4385),
.Y(n_4493)
);

INVx2_ASAP7_75t_SL g4494 ( 
.A(n_4396),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4432),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_4420),
.B(n_4323),
.Y(n_4496)
);

OR2x2_ASAP7_75t_L g4497 ( 
.A(n_4470),
.B(n_4354),
.Y(n_4497)
);

BUFx6f_ASAP7_75t_L g4498 ( 
.A(n_4382),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4387),
.Y(n_4499)
);

HB1xp67_ASAP7_75t_L g4500 ( 
.A(n_4398),
.Y(n_4500)
);

BUFx3_ASAP7_75t_L g4501 ( 
.A(n_4389),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_4425),
.B(n_4325),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4438),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_4453),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4433),
.B(n_4332),
.Y(n_4505)
);

BUFx3_ASAP7_75t_L g4506 ( 
.A(n_4424),
.Y(n_4506)
);

INVx2_ASAP7_75t_L g4507 ( 
.A(n_4397),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4434),
.B(n_4335),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4399),
.B(n_4407),
.Y(n_4509)
);

BUFx2_ASAP7_75t_L g4510 ( 
.A(n_4426),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4403),
.Y(n_4511)
);

BUFx2_ASAP7_75t_L g4512 ( 
.A(n_4435),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4404),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4410),
.Y(n_4514)
);

OAI22xp5_ASAP7_75t_L g4515 ( 
.A1(n_4383),
.A2(n_4351),
.B1(n_3816),
.B2(n_4298),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4415),
.B(n_4338),
.Y(n_4516)
);

INVx2_ASAP7_75t_L g4517 ( 
.A(n_4414),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4392),
.B(n_4341),
.Y(n_4518)
);

OR2x2_ASAP7_75t_L g4519 ( 
.A(n_4431),
.B(n_4273),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4416),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4423),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_4439),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4443),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4454),
.Y(n_4524)
);

AND2x2_ASAP7_75t_L g4525 ( 
.A(n_4459),
.B(n_4347),
.Y(n_4525)
);

AND2x4_ASAP7_75t_L g4526 ( 
.A(n_4408),
.B(n_4333),
.Y(n_4526)
);

BUFx2_ASAP7_75t_L g4527 ( 
.A(n_4393),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4441),
.B(n_4471),
.Y(n_4528)
);

INVx2_ASAP7_75t_L g4529 ( 
.A(n_4467),
.Y(n_4529)
);

AND2x6_ASAP7_75t_L g4530 ( 
.A(n_4384),
.B(n_4380),
.Y(n_4530)
);

AND2x2_ASAP7_75t_L g4531 ( 
.A(n_4413),
.B(n_4463),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4456),
.B(n_4251),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4461),
.B(n_4254),
.Y(n_4533)
);

AND2x2_ASAP7_75t_L g4534 ( 
.A(n_4474),
.B(n_4304),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4450),
.Y(n_4535)
);

AND2x2_ASAP7_75t_L g4536 ( 
.A(n_4472),
.B(n_4328),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4386),
.B(n_4278),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4465),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4465),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4445),
.B(n_4380),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4455),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4400),
.B(n_4283),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4400),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4412),
.Y(n_4544)
);

INVx1_ASAP7_75t_SL g4545 ( 
.A(n_4391),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4412),
.B(n_4284),
.Y(n_4546)
);

OAI21xp5_ASAP7_75t_L g4547 ( 
.A1(n_4444),
.A2(n_4324),
.B(n_4297),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4417),
.B(n_4299),
.Y(n_4548)
);

NOR2xp33_ASAP7_75t_L g4549 ( 
.A(n_4406),
.B(n_3675),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_4430),
.Y(n_4550)
);

OAI21x1_ASAP7_75t_L g4551 ( 
.A1(n_4479),
.A2(n_4345),
.B(n_4371),
.Y(n_4551)
);

AOI211xp5_ASAP7_75t_L g4552 ( 
.A1(n_4515),
.A2(n_4446),
.B(n_4418),
.C(n_4381),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4519),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4527),
.B(n_4430),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4535),
.B(n_4293),
.Y(n_4555)
);

NOR2x1_ASAP7_75t_L g4556 ( 
.A(n_4481),
.B(n_4512),
.Y(n_4556)
);

HB1xp67_ASAP7_75t_L g4557 ( 
.A(n_4480),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4484),
.Y(n_4558)
);

AOI21xp5_ASAP7_75t_L g4559 ( 
.A1(n_4510),
.A2(n_4402),
.B(n_4460),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4479),
.B(n_4449),
.Y(n_4560)
);

INVx2_ASAP7_75t_L g4561 ( 
.A(n_4477),
.Y(n_4561)
);

INVx2_ASAP7_75t_L g4562 ( 
.A(n_4482),
.Y(n_4562)
);

OAI211xp5_ASAP7_75t_L g4563 ( 
.A1(n_4475),
.A2(n_4405),
.B(n_4422),
.C(n_4437),
.Y(n_4563)
);

CKINVDCx5p33_ASAP7_75t_R g4564 ( 
.A(n_4493),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4476),
.Y(n_4565)
);

AO31x2_ASAP7_75t_L g4566 ( 
.A1(n_4529),
.A2(n_4451),
.A3(n_4375),
.B(n_4294),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4478),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4478),
.Y(n_4568)
);

AO21x2_ASAP7_75t_L g4569 ( 
.A1(n_4547),
.A2(n_4457),
.B(n_4373),
.Y(n_4569)
);

INVx3_ASAP7_75t_L g4570 ( 
.A(n_4506),
.Y(n_4570)
);

AND2x2_ASAP7_75t_L g4571 ( 
.A(n_4489),
.B(n_4448),
.Y(n_4571)
);

NOR2xp67_ASAP7_75t_L g4572 ( 
.A(n_4526),
.B(n_4452),
.Y(n_4572)
);

NOR2xp33_ASAP7_75t_R g4573 ( 
.A(n_4492),
.B(n_4462),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4486),
.Y(n_4574)
);

OR2x2_ASAP7_75t_L g4575 ( 
.A(n_4528),
.B(n_4286),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4499),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4499),
.Y(n_4577)
);

INVxp67_ASAP7_75t_SL g4578 ( 
.A(n_4500),
.Y(n_4578)
);

INVx3_ASAP7_75t_L g4579 ( 
.A(n_4501),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4495),
.Y(n_4580)
);

BUFx2_ASAP7_75t_L g4581 ( 
.A(n_4530),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_4513),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4513),
.Y(n_4583)
);

OA21x2_ASAP7_75t_L g4584 ( 
.A1(n_4540),
.A2(n_4378),
.B(n_4359),
.Y(n_4584)
);

HB1xp67_ASAP7_75t_L g4585 ( 
.A(n_4514),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_4507),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4514),
.Y(n_4587)
);

OAI21x1_ASAP7_75t_L g4588 ( 
.A1(n_4548),
.A2(n_4346),
.B(n_4366),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4511),
.Y(n_4589)
);

NOR2x1_ASAP7_75t_L g4590 ( 
.A(n_4483),
.B(n_4440),
.Y(n_4590)
);

OA21x2_ASAP7_75t_L g4591 ( 
.A1(n_4541),
.A2(n_4353),
.B(n_4365),
.Y(n_4591)
);

NOR2xp33_ASAP7_75t_L g4592 ( 
.A(n_4545),
.B(n_4469),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4496),
.B(n_4296),
.Y(n_4593)
);

AO21x2_ASAP7_75t_L g4594 ( 
.A1(n_4538),
.A2(n_4133),
.B(n_4236),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4520),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_4517),
.Y(n_4596)
);

AOI21xp5_ASAP7_75t_L g4597 ( 
.A1(n_4526),
.A2(n_4464),
.B(n_4226),
.Y(n_4597)
);

HB1xp67_ASAP7_75t_L g4598 ( 
.A(n_4524),
.Y(n_4598)
);

INVx2_ASAP7_75t_L g4599 ( 
.A(n_4521),
.Y(n_4599)
);

OR2x2_ASAP7_75t_L g4600 ( 
.A(n_4497),
.B(n_4287),
.Y(n_4600)
);

INVxp67_ASAP7_75t_L g4601 ( 
.A(n_4494),
.Y(n_4601)
);

AND2x6_ASAP7_75t_L g4602 ( 
.A(n_4531),
.B(n_4235),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4524),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4488),
.B(n_4292),
.Y(n_4604)
);

AOI22xp33_ASAP7_75t_L g4605 ( 
.A1(n_4536),
.A2(n_3972),
.B1(n_3984),
.B2(n_3981),
.Y(n_4605)
);

BUFx2_ASAP7_75t_L g4606 ( 
.A(n_4530),
.Y(n_4606)
);

NAND3xp33_ASAP7_75t_SL g4607 ( 
.A(n_4539),
.B(n_4224),
.C(n_4014),
.Y(n_4607)
);

AND2x2_ASAP7_75t_L g4608 ( 
.A(n_4485),
.B(n_4362),
.Y(n_4608)
);

NAND4xp25_ASAP7_75t_L g4609 ( 
.A(n_4549),
.B(n_4189),
.C(n_4195),
.D(n_4038),
.Y(n_4609)
);

HB1xp67_ASAP7_75t_L g4610 ( 
.A(n_4557),
.Y(n_4610)
);

INVx5_ASAP7_75t_L g4611 ( 
.A(n_4602),
.Y(n_4611)
);

INVx2_ASAP7_75t_L g4612 ( 
.A(n_4558),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4578),
.Y(n_4613)
);

AOI22xp5_ASAP7_75t_L g4614 ( 
.A1(n_4552),
.A2(n_4530),
.B1(n_4534),
.B2(n_4537),
.Y(n_4614)
);

INVx2_ASAP7_75t_L g4615 ( 
.A(n_4562),
.Y(n_4615)
);

INVx3_ASAP7_75t_L g4616 ( 
.A(n_4581),
.Y(n_4616)
);

INVx2_ASAP7_75t_L g4617 ( 
.A(n_4574),
.Y(n_4617)
);

AND2x2_ASAP7_75t_L g4618 ( 
.A(n_4560),
.B(n_4532),
.Y(n_4618)
);

AND2x2_ASAP7_75t_L g4619 ( 
.A(n_4590),
.B(n_4556),
.Y(n_4619)
);

INVxp67_ASAP7_75t_L g4620 ( 
.A(n_4570),
.Y(n_4620)
);

INVx1_ASAP7_75t_L g4621 ( 
.A(n_4582),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4585),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_L g4623 ( 
.A(n_4553),
.B(n_4533),
.Y(n_4623)
);

HB1xp67_ASAP7_75t_L g4624 ( 
.A(n_4598),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4555),
.Y(n_4625)
);

AND2x2_ASAP7_75t_L g4626 ( 
.A(n_4554),
.B(n_4509),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4576),
.Y(n_4627)
);

INVx4_ASAP7_75t_L g4628 ( 
.A(n_4564),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4594),
.B(n_4593),
.Y(n_4629)
);

INVx1_ASAP7_75t_SL g4630 ( 
.A(n_4579),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4581),
.B(n_4542),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4580),
.Y(n_4632)
);

BUFx2_ASAP7_75t_L g4633 ( 
.A(n_4602),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4606),
.B(n_4572),
.Y(n_4634)
);

OAI31xp33_ASAP7_75t_L g4635 ( 
.A1(n_4563),
.A2(n_4543),
.A3(n_4544),
.B(n_4092),
.Y(n_4635)
);

NOR3xp33_ASAP7_75t_SL g4636 ( 
.A(n_4607),
.B(n_4184),
.C(n_4246),
.Y(n_4636)
);

OR2x2_ASAP7_75t_L g4637 ( 
.A(n_4600),
.B(n_4490),
.Y(n_4637)
);

OAI22xp5_ASAP7_75t_L g4638 ( 
.A1(n_4606),
.A2(n_4504),
.B1(n_4503),
.B2(n_4550),
.Y(n_4638)
);

INVx2_ASAP7_75t_L g4639 ( 
.A(n_4586),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4571),
.B(n_4546),
.Y(n_4640)
);

AND2x2_ASAP7_75t_L g4641 ( 
.A(n_4601),
.B(n_4608),
.Y(n_4641)
);

AND2x2_ASAP7_75t_L g4642 ( 
.A(n_4602),
.B(n_4604),
.Y(n_4642)
);

AND2x4_ASAP7_75t_L g4643 ( 
.A(n_4597),
.B(n_4498),
.Y(n_4643)
);

INVx1_ASAP7_75t_SL g4644 ( 
.A(n_4573),
.Y(n_4644)
);

HB1xp67_ASAP7_75t_L g4645 ( 
.A(n_4565),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4577),
.B(n_4502),
.Y(n_4646)
);

OAI222xp33_ASAP7_75t_L g4647 ( 
.A1(n_4559),
.A2(n_4491),
.B1(n_4487),
.B2(n_4516),
.C1(n_4518),
.C2(n_4508),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4583),
.Y(n_4648)
);

AND2x2_ASAP7_75t_L g4649 ( 
.A(n_4566),
.B(n_4498),
.Y(n_4649)
);

OAI21x1_ASAP7_75t_L g4650 ( 
.A1(n_4551),
.A2(n_4523),
.B(n_4522),
.Y(n_4650)
);

AND2x2_ASAP7_75t_L g4651 ( 
.A(n_4566),
.B(n_4525),
.Y(n_4651)
);

HB1xp67_ASAP7_75t_L g4652 ( 
.A(n_4567),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_4587),
.B(n_4505),
.Y(n_4653)
);

AOI22xp33_ASAP7_75t_L g4654 ( 
.A1(n_4609),
.A2(n_4569),
.B1(n_4591),
.B2(n_4605),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4595),
.Y(n_4655)
);

INVxp67_ASAP7_75t_L g4656 ( 
.A(n_4592),
.Y(n_4656)
);

OR2x2_ASAP7_75t_L g4657 ( 
.A(n_4575),
.B(n_4128),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4603),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4568),
.B(n_4128),
.Y(n_4659)
);

AOI22xp33_ASAP7_75t_SL g4660 ( 
.A1(n_4591),
.A2(n_4584),
.B1(n_4464),
.B2(n_4561),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4589),
.Y(n_4661)
);

NOR2x1_ASAP7_75t_L g4662 ( 
.A(n_4596),
.B(n_4134),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4599),
.B(n_4362),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4637),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4613),
.B(n_4588),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4610),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4619),
.B(n_3904),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4624),
.Y(n_4668)
);

BUFx2_ASAP7_75t_L g4669 ( 
.A(n_4643),
.Y(n_4669)
);

AND2x2_ASAP7_75t_L g4670 ( 
.A(n_4611),
.B(n_3917),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4646),
.Y(n_4671)
);

HB1xp67_ASAP7_75t_L g4672 ( 
.A(n_4621),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4622),
.Y(n_4673)
);

NAND2x1p5_ASAP7_75t_L g4674 ( 
.A(n_4628),
.B(n_4242),
.Y(n_4674)
);

AND2x2_ASAP7_75t_L g4675 ( 
.A(n_4634),
.B(n_3935),
.Y(n_4675)
);

AND2x4_ASAP7_75t_L g4676 ( 
.A(n_4630),
.B(n_3748),
.Y(n_4676)
);

NAND5xp2_ASAP7_75t_L g4677 ( 
.A(n_4635),
.B(n_4089),
.C(n_3744),
.D(n_4090),
.E(n_3862),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4643),
.B(n_4633),
.Y(n_4678)
);

INVx2_ASAP7_75t_L g4679 ( 
.A(n_4612),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4645),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4625),
.B(n_4118),
.Y(n_4681)
);

OR2x2_ASAP7_75t_L g4682 ( 
.A(n_4657),
.B(n_4659),
.Y(n_4682)
);

OR2x2_ASAP7_75t_L g4683 ( 
.A(n_4629),
.B(n_4159),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4652),
.Y(n_4684)
);

INVx1_ASAP7_75t_SL g4685 ( 
.A(n_4644),
.Y(n_4685)
);

AND2x2_ASAP7_75t_L g4686 ( 
.A(n_4642),
.B(n_3993),
.Y(n_4686)
);

AND2x2_ASAP7_75t_L g4687 ( 
.A(n_4618),
.B(n_3996),
.Y(n_4687)
);

OR2x2_ASAP7_75t_L g4688 ( 
.A(n_4616),
.B(n_4159),
.Y(n_4688)
);

INVx2_ASAP7_75t_L g4689 ( 
.A(n_4615),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4620),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4653),
.Y(n_4691)
);

AND2x2_ASAP7_75t_L g4692 ( 
.A(n_4631),
.B(n_4079),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4623),
.Y(n_4693)
);

AND2x2_ASAP7_75t_L g4694 ( 
.A(n_4641),
.B(n_4120),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4627),
.Y(n_4695)
);

INVx5_ASAP7_75t_L g4696 ( 
.A(n_4628),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4648),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4655),
.Y(n_4698)
);

BUFx3_ASAP7_75t_L g4699 ( 
.A(n_4663),
.Y(n_4699)
);

OR2x2_ASAP7_75t_L g4700 ( 
.A(n_4666),
.B(n_4616),
.Y(n_4700)
);

OR2x2_ASAP7_75t_L g4701 ( 
.A(n_4664),
.B(n_4638),
.Y(n_4701)
);

INVx2_ASAP7_75t_L g4702 ( 
.A(n_4690),
.Y(n_4702)
);

OR2x2_ASAP7_75t_L g4703 ( 
.A(n_4668),
.B(n_4681),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4672),
.Y(n_4704)
);

NAND2x1_ASAP7_75t_L g4705 ( 
.A(n_4669),
.B(n_4676),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4678),
.B(n_4656),
.Y(n_4706)
);

OR2x2_ASAP7_75t_L g4707 ( 
.A(n_4679),
.B(n_4614),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4680),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4680),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4693),
.B(n_4636),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4685),
.B(n_4654),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4699),
.B(n_4626),
.Y(n_4712)
);

INVxp67_ASAP7_75t_L g4713 ( 
.A(n_4676),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4689),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4684),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4673),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4674),
.Y(n_4717)
);

INVx2_ASAP7_75t_L g4718 ( 
.A(n_4675),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4695),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_4696),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4691),
.Y(n_4721)
);

INVx3_ASAP7_75t_L g4722 ( 
.A(n_4696),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4671),
.B(n_4662),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4694),
.B(n_4640),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4696),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4695),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4697),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_4667),
.B(n_4670),
.Y(n_4728)
);

INVx1_ASAP7_75t_SL g4729 ( 
.A(n_4686),
.Y(n_4729)
);

INVx2_ASAP7_75t_L g4730 ( 
.A(n_4697),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4698),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4698),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_4706),
.B(n_4665),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4704),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_4712),
.B(n_4692),
.Y(n_4735)
);

NOR2x1_ASAP7_75t_L g4736 ( 
.A(n_4722),
.B(n_4677),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4702),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4700),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4701),
.Y(n_4739)
);

AOI22xp5_ASAP7_75t_L g4740 ( 
.A1(n_4713),
.A2(n_4687),
.B1(n_4683),
.B2(n_4660),
.Y(n_4740)
);

NAND3x1_ASAP7_75t_L g4741 ( 
.A(n_4711),
.B(n_4649),
.C(n_4651),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4728),
.B(n_4682),
.Y(n_4742)
);

OR2x2_ASAP7_75t_L g4743 ( 
.A(n_4710),
.B(n_4688),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4720),
.B(n_4725),
.Y(n_4744)
);

OR2x2_ASAP7_75t_L g4745 ( 
.A(n_4714),
.B(n_4661),
.Y(n_4745)
);

HB1xp67_ASAP7_75t_L g4746 ( 
.A(n_4708),
.Y(n_4746)
);

AOI22xp33_ASAP7_75t_L g4747 ( 
.A1(n_4717),
.A2(n_4707),
.B1(n_4705),
.B2(n_4718),
.Y(n_4747)
);

INVx2_ASAP7_75t_SL g4748 ( 
.A(n_4729),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4709),
.Y(n_4749)
);

AND2x2_ASAP7_75t_L g4750 ( 
.A(n_4724),
.B(n_4658),
.Y(n_4750)
);

INVx2_ASAP7_75t_SL g4751 ( 
.A(n_4715),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4730),
.Y(n_4752)
);

OR2x2_ASAP7_75t_L g4753 ( 
.A(n_4703),
.B(n_4639),
.Y(n_4753)
);

INVx1_ASAP7_75t_SL g4754 ( 
.A(n_4723),
.Y(n_4754)
);

BUFx3_ASAP7_75t_L g4755 ( 
.A(n_4721),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4719),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4719),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4731),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4731),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4732),
.Y(n_4760)
);

AND2x2_ASAP7_75t_L g4761 ( 
.A(n_4716),
.B(n_4617),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4726),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4727),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4706),
.Y(n_4764)
);

AND2x4_ASAP7_75t_L g4765 ( 
.A(n_4713),
.B(n_4632),
.Y(n_4765)
);

NAND2x1_ASAP7_75t_L g4766 ( 
.A(n_4722),
.B(n_4647),
.Y(n_4766)
);

INVx1_ASAP7_75t_SL g4767 ( 
.A(n_4705),
.Y(n_4767)
);

NOR2x1_ASAP7_75t_L g4768 ( 
.A(n_4736),
.B(n_4744),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4735),
.B(n_4650),
.Y(n_4769)
);

HB1xp67_ASAP7_75t_L g4770 ( 
.A(n_4764),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4739),
.Y(n_4771)
);

OR2x2_ASAP7_75t_L g4772 ( 
.A(n_4748),
.B(n_660),
.Y(n_4772)
);

INVxp67_ASAP7_75t_L g4773 ( 
.A(n_4767),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4747),
.B(n_4742),
.Y(n_4774)
);

INVx1_ASAP7_75t_SL g4775 ( 
.A(n_4765),
.Y(n_4775)
);

INVxp33_ASAP7_75t_L g4776 ( 
.A(n_4765),
.Y(n_4776)
);

INVx1_ASAP7_75t_SL g4777 ( 
.A(n_4755),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4738),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4753),
.Y(n_4779)
);

AND2x2_ASAP7_75t_L g4780 ( 
.A(n_4750),
.B(n_4151),
.Y(n_4780)
);

BUFx2_ASAP7_75t_L g4781 ( 
.A(n_4737),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4745),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_4754),
.B(n_4205),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4740),
.B(n_4761),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4733),
.B(n_4207),
.Y(n_4785)
);

INVx2_ASAP7_75t_L g4786 ( 
.A(n_4752),
.Y(n_4786)
);

NAND4xp25_ASAP7_75t_L g4787 ( 
.A(n_4743),
.B(n_4003),
.C(n_3992),
.D(n_3798),
.Y(n_4787)
);

OR2x2_ASAP7_75t_L g4788 ( 
.A(n_4751),
.B(n_661),
.Y(n_4788)
);

INVx2_ASAP7_75t_L g4789 ( 
.A(n_4734),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_4746),
.B(n_3948),
.Y(n_4790)
);

AND2x2_ASAP7_75t_L g4791 ( 
.A(n_4766),
.B(n_4151),
.Y(n_4791)
);

OAI22xp33_ASAP7_75t_L g4792 ( 
.A1(n_4749),
.A2(n_3989),
.B1(n_3942),
.B2(n_3986),
.Y(n_4792)
);

OR2x2_ASAP7_75t_L g4793 ( 
.A(n_4762),
.B(n_661),
.Y(n_4793)
);

NOR2x1p5_ASAP7_75t_L g4794 ( 
.A(n_4763),
.B(n_4239),
.Y(n_4794)
);

INVx3_ASAP7_75t_L g4795 ( 
.A(n_4741),
.Y(n_4795)
);

OR2x2_ASAP7_75t_L g4796 ( 
.A(n_4760),
.B(n_662),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4756),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4757),
.Y(n_4798)
);

AND2x2_ASAP7_75t_L g4799 ( 
.A(n_4758),
.B(n_3931),
.Y(n_4799)
);

INVx2_ASAP7_75t_SL g4800 ( 
.A(n_4759),
.Y(n_4800)
);

INVx1_ASAP7_75t_SL g4801 ( 
.A(n_4767),
.Y(n_4801)
);

NOR2x1_ASAP7_75t_L g4802 ( 
.A(n_4736),
.B(n_3967),
.Y(n_4802)
);

HB1xp67_ASAP7_75t_L g4803 ( 
.A(n_4779),
.Y(n_4803)
);

AOI21xp5_ASAP7_75t_L g4804 ( 
.A1(n_4801),
.A2(n_3943),
.B(n_3860),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4772),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4781),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4774),
.B(n_3981),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4770),
.Y(n_4808)
);

INVx2_ASAP7_75t_L g4809 ( 
.A(n_4777),
.Y(n_4809)
);

NOR2xp33_ASAP7_75t_L g4810 ( 
.A(n_4776),
.B(n_4795),
.Y(n_4810)
);

INVx2_ASAP7_75t_L g4811 ( 
.A(n_4786),
.Y(n_4811)
);

OAI21xp5_ASAP7_75t_L g4812 ( 
.A1(n_4768),
.A2(n_4227),
.B(n_4222),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_4782),
.Y(n_4813)
);

AOI31xp33_ASAP7_75t_L g4814 ( 
.A1(n_4771),
.A2(n_3967),
.A3(n_3942),
.B(n_3877),
.Y(n_4814)
);

AND2x2_ASAP7_75t_L g4815 ( 
.A(n_4784),
.B(n_4176),
.Y(n_4815)
);

HB1xp67_ASAP7_75t_L g4816 ( 
.A(n_4788),
.Y(n_4816)
);

OAI21xp33_ASAP7_75t_L g4817 ( 
.A1(n_4802),
.A2(n_4180),
.B(n_4066),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4769),
.B(n_4799),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4796),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4793),
.Y(n_4820)
);

OAI21xp33_ASAP7_75t_SL g4821 ( 
.A1(n_4795),
.A2(n_4229),
.B(n_4131),
.Y(n_4821)
);

AOI221xp5_ASAP7_75t_SL g4822 ( 
.A1(n_4778),
.A2(n_3819),
.B1(n_4000),
.B2(n_3932),
.C(n_3813),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4789),
.Y(n_4823)
);

O2A1O1Ixp33_ASAP7_75t_L g4824 ( 
.A1(n_4800),
.A2(n_4086),
.B(n_3775),
.C(n_3913),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4783),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4791),
.B(n_663),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4790),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4798),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4798),
.Y(n_4829)
);

OAI33xp33_ASAP7_75t_L g4830 ( 
.A1(n_4797),
.A2(n_665),
.A3(n_667),
.B1(n_663),
.B2(n_664),
.B3(n_666),
.Y(n_4830)
);

NOR2xp33_ASAP7_75t_L g4831 ( 
.A(n_4785),
.B(n_3733),
.Y(n_4831)
);

OAI22xp5_ASAP7_75t_L g4832 ( 
.A1(n_4780),
.A2(n_3891),
.B1(n_3954),
.B2(n_4083),
.Y(n_4832)
);

OAI22xp5_ASAP7_75t_L g4833 ( 
.A1(n_4794),
.A2(n_3973),
.B1(n_4073),
.B2(n_3895),
.Y(n_4833)
);

OAI21xp5_ASAP7_75t_SL g4834 ( 
.A1(n_4787),
.A2(n_3946),
.B(n_3944),
.Y(n_4834)
);

AOI211xp5_ASAP7_75t_L g4835 ( 
.A1(n_4792),
.A2(n_4238),
.B(n_4201),
.C(n_4140),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4779),
.Y(n_4836)
);

O2A1O1Ixp33_ASAP7_75t_L g4837 ( 
.A1(n_4773),
.A2(n_4199),
.B(n_4093),
.C(n_4067),
.Y(n_4837)
);

OR2x2_ASAP7_75t_L g4838 ( 
.A(n_4775),
.B(n_664),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4774),
.B(n_665),
.Y(n_4839)
);

OAI22xp5_ASAP7_75t_L g4840 ( 
.A1(n_4773),
.A2(n_3747),
.B1(n_3916),
.B2(n_3912),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4774),
.B(n_666),
.Y(n_4841)
);

OAI211xp5_ASAP7_75t_SL g4842 ( 
.A1(n_4773),
.A2(n_670),
.B(n_668),
.C(n_669),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4809),
.B(n_668),
.Y(n_4843)
);

INVx2_ASAP7_75t_L g4844 ( 
.A(n_4811),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4838),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4803),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4806),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4818),
.B(n_670),
.Y(n_4848)
);

NAND4xp25_ASAP7_75t_L g4849 ( 
.A(n_4810),
.B(n_673),
.C(n_671),
.D(n_672),
.Y(n_4849)
);

OR2x2_ASAP7_75t_L g4850 ( 
.A(n_4839),
.B(n_672),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4841),
.B(n_672),
.Y(n_4851)
);

OR2x2_ASAP7_75t_L g4852 ( 
.A(n_4808),
.B(n_674),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4816),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4813),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4836),
.Y(n_4855)
);

INVx2_ASAP7_75t_SL g4856 ( 
.A(n_4807),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4804),
.B(n_674),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4823),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4805),
.Y(n_4859)
);

NOR2xp33_ASAP7_75t_L g4860 ( 
.A(n_4830),
.B(n_675),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4815),
.B(n_676),
.Y(n_4861)
);

CKINVDCx11_ASAP7_75t_R g4862 ( 
.A(n_4819),
.Y(n_4862)
);

INVxp67_ASAP7_75t_L g4863 ( 
.A(n_4820),
.Y(n_4863)
);

NAND2xp5_ASAP7_75t_L g4864 ( 
.A(n_4822),
.B(n_677),
.Y(n_4864)
);

INVx2_ASAP7_75t_L g4865 ( 
.A(n_4827),
.Y(n_4865)
);

NOR2xp33_ASAP7_75t_L g4866 ( 
.A(n_4826),
.B(n_677),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4828),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4829),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4814),
.Y(n_4869)
);

A2O1A1Ixp33_ASAP7_75t_L g4870 ( 
.A1(n_4824),
.A2(n_4831),
.B(n_4825),
.C(n_4842),
.Y(n_4870)
);

NAND3xp33_ASAP7_75t_L g4871 ( 
.A(n_4812),
.B(n_677),
.C(n_678),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4817),
.B(n_678),
.Y(n_4872)
);

OAI21xp33_ASAP7_75t_SL g4873 ( 
.A1(n_4832),
.A2(n_4169),
.B(n_4160),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4834),
.B(n_680),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4833),
.Y(n_4875)
);

AND2x2_ASAP7_75t_L g4876 ( 
.A(n_4848),
.B(n_4856),
.Y(n_4876)
);

INVxp67_ASAP7_75t_SL g4877 ( 
.A(n_4843),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4860),
.B(n_4840),
.Y(n_4878)
);

INVx1_ASAP7_75t_SL g4879 ( 
.A(n_4862),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4844),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4853),
.B(n_4821),
.Y(n_4881)
);

INVx1_ASAP7_75t_L g4882 ( 
.A(n_4852),
.Y(n_4882)
);

OR2x2_ASAP7_75t_L g4883 ( 
.A(n_4849),
.B(n_680),
.Y(n_4883)
);

NOR2xp33_ASAP7_75t_L g4884 ( 
.A(n_4871),
.B(n_4854),
.Y(n_4884)
);

NOR2xp33_ASAP7_75t_R g4885 ( 
.A(n_4847),
.B(n_681),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4846),
.B(n_4837),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4845),
.B(n_4835),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4857),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4874),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4858),
.Y(n_4890)
);

NAND2x1p5_ASAP7_75t_L g4891 ( 
.A(n_4865),
.B(n_3740),
.Y(n_4891)
);

AND2x2_ASAP7_75t_L g4892 ( 
.A(n_4869),
.B(n_682),
.Y(n_4892)
);

AND2x2_ASAP7_75t_L g4893 ( 
.A(n_4866),
.B(n_682),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4851),
.Y(n_4894)
);

INVx2_ASAP7_75t_L g4895 ( 
.A(n_4859),
.Y(n_4895)
);

NOR2xp33_ASAP7_75t_L g4896 ( 
.A(n_4864),
.B(n_684),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4863),
.B(n_684),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4850),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4872),
.Y(n_4899)
);

OAI21xp33_ASAP7_75t_L g4900 ( 
.A1(n_4870),
.A2(n_4190),
.B(n_4179),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4861),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4855),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4875),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_4867),
.B(n_684),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4868),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4873),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4873),
.B(n_685),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4848),
.B(n_685),
.Y(n_4908)
);

OAI21xp5_ASAP7_75t_L g4909 ( 
.A1(n_4879),
.A2(n_4125),
.B(n_4123),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4876),
.Y(n_4910)
);

NAND4xp25_ASAP7_75t_L g4911 ( 
.A(n_4878),
.B(n_688),
.C(n_686),
.D(n_687),
.Y(n_4911)
);

NOR3xp33_ASAP7_75t_L g4912 ( 
.A(n_4880),
.B(n_687),
.C(n_688),
.Y(n_4912)
);

AOI211xp5_ASAP7_75t_L g4913 ( 
.A1(n_4896),
.A2(n_4127),
.B(n_4170),
.C(n_4158),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4883),
.Y(n_4914)
);

NAND2xp33_ASAP7_75t_L g4915 ( 
.A(n_4903),
.B(n_3703),
.Y(n_4915)
);

NAND3xp33_ASAP7_75t_L g4916 ( 
.A(n_4884),
.B(n_687),
.C(n_689),
.Y(n_4916)
);

OAI221xp5_ASAP7_75t_L g4917 ( 
.A1(n_4900),
.A2(n_3778),
.B1(n_3804),
.B2(n_3792),
.C(n_3797),
.Y(n_4917)
);

NAND4xp25_ASAP7_75t_L g4918 ( 
.A(n_4892),
.B(n_691),
.C(n_689),
.D(n_690),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_4906),
.B(n_689),
.Y(n_4919)
);

AND2x2_ASAP7_75t_L g4920 ( 
.A(n_4893),
.B(n_691),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_SL g4921 ( 
.A(n_4907),
.B(n_3778),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_SL g4922 ( 
.A(n_4881),
.B(n_3804),
.Y(n_4922)
);

INVx1_ASAP7_75t_SL g4923 ( 
.A(n_4891),
.Y(n_4923)
);

NOR3xp33_ASAP7_75t_L g4924 ( 
.A(n_4897),
.B(n_4895),
.C(n_4890),
.Y(n_4924)
);

OAI22xp5_ASAP7_75t_L g4925 ( 
.A1(n_4908),
.A2(n_3884),
.B1(n_4063),
.B2(n_4110),
.Y(n_4925)
);

OAI211xp5_ASAP7_75t_L g4926 ( 
.A1(n_4885),
.A2(n_694),
.B(n_692),
.C(n_693),
.Y(n_4926)
);

AO21x1_ASAP7_75t_L g4927 ( 
.A1(n_4904),
.A2(n_4135),
.B(n_4143),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_L g4928 ( 
.A(n_4890),
.B(n_692),
.Y(n_4928)
);

OR2x2_ASAP7_75t_L g4929 ( 
.A(n_4882),
.B(n_693),
.Y(n_4929)
);

NAND3xp33_ASAP7_75t_L g4930 ( 
.A(n_4905),
.B(n_4902),
.C(n_4889),
.Y(n_4930)
);

NAND4xp25_ASAP7_75t_L g4931 ( 
.A(n_4887),
.B(n_4898),
.C(n_4901),
.D(n_4899),
.Y(n_4931)
);

AOI222xp33_ASAP7_75t_L g4932 ( 
.A1(n_4886),
.A2(n_4217),
.B1(n_3764),
.B2(n_3774),
.C1(n_3781),
.C2(n_3776),
.Y(n_4932)
);

AND2x2_ASAP7_75t_L g4933 ( 
.A(n_4877),
.B(n_695),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4888),
.Y(n_4934)
);

NOR2xp33_ASAP7_75t_SL g4935 ( 
.A(n_4894),
.B(n_3787),
.Y(n_4935)
);

AOI22xp33_ASAP7_75t_L g4936 ( 
.A1(n_4912),
.A2(n_4088),
.B1(n_3803),
.B2(n_3769),
.Y(n_4936)
);

AOI222xp33_ASAP7_75t_L g4937 ( 
.A1(n_4919),
.A2(n_4915),
.B1(n_4910),
.B2(n_4923),
.C1(n_4922),
.C2(n_4914),
.Y(n_4937)
);

AOI211x1_ASAP7_75t_SL g4938 ( 
.A1(n_4931),
.A2(n_4930),
.B(n_4921),
.C(n_4918),
.Y(n_4938)
);

OAI21xp5_ASAP7_75t_L g4939 ( 
.A1(n_4916),
.A2(n_4075),
.B(n_4106),
.Y(n_4939)
);

OAI211xp5_ASAP7_75t_L g4940 ( 
.A1(n_4928),
.A2(n_4933),
.B(n_4924),
.C(n_4929),
.Y(n_4940)
);

NAND4xp75_ASAP7_75t_L g4941 ( 
.A(n_4934),
.B(n_699),
.C(n_697),
.D(n_698),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_L g4942 ( 
.A(n_4920),
.B(n_699),
.Y(n_4942)
);

AOI211xp5_ASAP7_75t_L g4943 ( 
.A1(n_4909),
.A2(n_4935),
.B(n_4927),
.C(n_4917),
.Y(n_4943)
);

AOI221xp5_ASAP7_75t_L g4944 ( 
.A1(n_4925),
.A2(n_702),
.B1(n_700),
.B2(n_701),
.C(n_703),
.Y(n_4944)
);

OAI21xp33_ASAP7_75t_SL g4945 ( 
.A1(n_4932),
.A2(n_4913),
.B(n_4108),
.Y(n_4945)
);

AOI211xp5_ASAP7_75t_L g4946 ( 
.A1(n_4926),
.A2(n_703),
.B(n_701),
.C(n_702),
.Y(n_4946)
);

AOI21xp5_ASAP7_75t_L g4947 ( 
.A1(n_4919),
.A2(n_701),
.B(n_703),
.Y(n_4947)
);

NAND3xp33_ASAP7_75t_SL g4948 ( 
.A(n_4912),
.B(n_704),
.C(n_705),
.Y(n_4948)
);

AOI211xp5_ASAP7_75t_SL g4949 ( 
.A1(n_4926),
.A2(n_709),
.B(n_706),
.C(n_708),
.Y(n_4949)
);

AOI221xp5_ASAP7_75t_L g4950 ( 
.A1(n_4911),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.C(n_711),
.Y(n_4950)
);

AOI221xp5_ASAP7_75t_L g4951 ( 
.A1(n_4911),
.A2(n_712),
.B1(n_710),
.B2(n_711),
.C(n_713),
.Y(n_4951)
);

AOI22xp33_ASAP7_75t_L g4952 ( 
.A1(n_4912),
.A2(n_4065),
.B1(n_3985),
.B2(n_3894),
.Y(n_4952)
);

AOI22xp5_ASAP7_75t_L g4953 ( 
.A1(n_4910),
.A2(n_3985),
.B1(n_3759),
.B2(n_4042),
.Y(n_4953)
);

AOI221x1_ASAP7_75t_L g4954 ( 
.A1(n_4947),
.A2(n_715),
.B1(n_712),
.B2(n_714),
.C(n_716),
.Y(n_4954)
);

NAND5xp2_ASAP7_75t_L g4955 ( 
.A(n_4949),
.B(n_716),
.C(n_714),
.D(n_715),
.E(n_774),
.Y(n_4955)
);

NAND3xp33_ASAP7_75t_L g4956 ( 
.A(n_4946),
.B(n_714),
.C(n_715),
.Y(n_4956)
);

XNOR2xp5_ASAP7_75t_L g4957 ( 
.A(n_4938),
.B(n_775),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4941),
.Y(n_4958)
);

BUFx2_ASAP7_75t_L g4959 ( 
.A(n_4945),
.Y(n_4959)
);

NAND4xp25_ASAP7_75t_L g4960 ( 
.A(n_4937),
.B(n_781),
.C(n_779),
.D(n_780),
.Y(n_4960)
);

AND2x2_ASAP7_75t_L g4961 ( 
.A(n_4942),
.B(n_4213),
.Y(n_4961)
);

AOI22xp5_ASAP7_75t_L g4962 ( 
.A1(n_4948),
.A2(n_4951),
.B1(n_4950),
.B2(n_4940),
.Y(n_4962)
);

AOI221xp5_ASAP7_75t_L g4963 ( 
.A1(n_4944),
.A2(n_786),
.B1(n_784),
.B2(n_785),
.C(n_787),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4943),
.B(n_786),
.Y(n_4964)
);

OR3x2_ASAP7_75t_L g4965 ( 
.A(n_4955),
.B(n_4960),
.C(n_4958),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4957),
.Y(n_4966)
);

NOR2x1_ASAP7_75t_L g4967 ( 
.A(n_4956),
.B(n_4939),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4964),
.B(n_4959),
.Y(n_4968)
);

AND4x1_ASAP7_75t_L g4969 ( 
.A(n_4962),
.B(n_4936),
.C(n_4952),
.D(n_4953),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4954),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4961),
.B(n_790),
.Y(n_4971)
);

NAND3xp33_ASAP7_75t_SL g4972 ( 
.A(n_4963),
.B(n_790),
.C(n_791),
.Y(n_4972)
);

NAND3x1_ASAP7_75t_L g4973 ( 
.A(n_4967),
.B(n_793),
.C(n_794),
.Y(n_4973)
);

HB1xp67_ASAP7_75t_L g4974 ( 
.A(n_4965),
.Y(n_4974)
);

NOR3xp33_ASAP7_75t_L g4975 ( 
.A(n_4968),
.B(n_4966),
.C(n_4970),
.Y(n_4975)
);

NOR3xp33_ASAP7_75t_SL g4976 ( 
.A(n_4972),
.B(n_799),
.C(n_800),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4971),
.Y(n_4977)
);

INVx2_ASAP7_75t_SL g4978 ( 
.A(n_4969),
.Y(n_4978)
);

CKINVDCx20_ASAP7_75t_R g4979 ( 
.A(n_4974),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4978),
.B(n_4975),
.Y(n_4980)
);

BUFx2_ASAP7_75t_L g4981 ( 
.A(n_4973),
.Y(n_4981)
);

CKINVDCx5p33_ASAP7_75t_R g4982 ( 
.A(n_4976),
.Y(n_4982)
);

CKINVDCx20_ASAP7_75t_R g4983 ( 
.A(n_4977),
.Y(n_4983)
);

AOI21xp5_ASAP7_75t_L g4984 ( 
.A1(n_4980),
.A2(n_803),
.B(n_804),
.Y(n_4984)
);

BUFx2_ASAP7_75t_L g4985 ( 
.A(n_4979),
.Y(n_4985)
);

OAI22x1_ASAP7_75t_L g4986 ( 
.A1(n_4982),
.A2(n_810),
.B1(n_805),
.B2(n_807),
.Y(n_4986)
);

XNOR2xp5_ASAP7_75t_L g4987 ( 
.A(n_4983),
.B(n_812),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4981),
.Y(n_4988)
);

INVx2_ASAP7_75t_L g4989 ( 
.A(n_4985),
.Y(n_4989)
);

AOI22xp5_ASAP7_75t_L g4990 ( 
.A1(n_4988),
.A2(n_3985),
.B1(n_814),
.B2(n_812),
.Y(n_4990)
);

INVx2_ASAP7_75t_SL g4991 ( 
.A(n_4989),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4991),
.B(n_4987),
.Y(n_4992)
);

INVx3_ASAP7_75t_L g4993 ( 
.A(n_4992),
.Y(n_4993)
);

INVx1_ASAP7_75t_SL g4994 ( 
.A(n_4993),
.Y(n_4994)
);

AOI22xp33_ASAP7_75t_L g4995 ( 
.A1(n_4994),
.A2(n_4986),
.B1(n_4984),
.B2(n_4990),
.Y(n_4995)
);

AOI22xp33_ASAP7_75t_SL g4996 ( 
.A1(n_4995),
.A2(n_818),
.B1(n_815),
.B2(n_816),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_SL g4997 ( 
.A(n_4996),
.B(n_821),
.Y(n_4997)
);

AOI21xp5_ASAP7_75t_L g4998 ( 
.A1(n_4997),
.A2(n_823),
.B(n_824),
.Y(n_4998)
);

AOI22xp5_ASAP7_75t_L g4999 ( 
.A1(n_4998),
.A2(n_829),
.B1(n_825),
.B2(n_827),
.Y(n_4999)
);


endmodule