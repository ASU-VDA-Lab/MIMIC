module fake_jpeg_19396_n_165 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_2),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_35),
.A3(n_39),
.B1(n_37),
.B2(n_42),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_52),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_55),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_54),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_62),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_2),
.Y(n_80)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_27),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_64),
.B(n_63),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_34),
.B1(n_16),
.B2(n_23),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_73),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_18),
.B1(n_25),
.B2(n_19),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_15),
.B(n_2),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_72),
.B(n_74),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_18),
.B1(n_19),
.B2(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_75),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_27),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_16),
.B1(n_26),
.B2(n_23),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_82),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_10),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_14),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_48),
.B1(n_59),
.B2(n_11),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_100),
.B1(n_90),
.B2(n_109),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_95),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_72),
.B(n_74),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_104),
.B(n_106),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_73),
.B(n_70),
.Y(n_121)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_85),
.B1(n_76),
.B2(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_118),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_117),
.B(n_124),
.Y(n_133)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_112),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_84),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_92),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_118),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_124),
.B1(n_114),
.B2(n_111),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_108),
.B1(n_107),
.B2(n_95),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_107),
.A3(n_96),
.B1(n_103),
.B2(n_89),
.C1(n_92),
.C2(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_128),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_130),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_89),
.B(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_131),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_120),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_122),
.C(n_115),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_138),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_134),
.Y(n_146)
);

INVxp33_ASAP7_75t_SL g144 ( 
.A(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_141),
.A2(n_133),
.B1(n_129),
.B2(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_126),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_148),
.B(n_137),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_133),
.B(n_116),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_136),
.Y(n_154)
);

NOR2x1_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_144),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_155),
.B(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_149),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_156),
.B(n_150),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_156),
.B(n_138),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_160),
.C(n_145),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);


endmodule