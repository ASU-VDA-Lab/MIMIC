module real_jpeg_12883_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_4),
.A2(n_37),
.B1(n_38),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_4),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_84),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_84),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_6),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_6),
.A2(n_41),
.B1(n_66),
.B2(n_67),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_8),
.A2(n_48),
.B1(n_66),
.B2(n_67),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_70),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_12),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_12),
.A2(n_37),
.B1(n_38),
.B2(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_13),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_13),
.B(n_140),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_104),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_13),
.B(n_67),
.C(n_87),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_13),
.B(n_36),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_13),
.A2(n_71),
.B(n_168),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_13),
.A2(n_27),
.B(n_35),
.C(n_195),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_104),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_14),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_14),
.A2(n_30),
.B1(n_66),
.B2(n_67),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_14),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_15),
.A2(n_66),
.B1(n_67),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_15),
.Y(n_116)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_106),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_92),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_21),
.A2(n_22),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_58),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_24),
.B(n_58),
.C(n_59),
.Y(n_125)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_26),
.A2(n_31),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_28),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AOI32xp33_ASAP7_75t_L g61 ( 
.A1(n_27),
.A2(n_45),
.A3(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_28),
.B(n_50),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_31),
.A2(n_39),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_32),
.B(n_40),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_34),
.A2(n_37),
.B(n_104),
.Y(n_195)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_37),
.A2(n_38),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_38),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_49),
.B(n_52),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_43),
.A2(n_49),
.B1(n_54),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_54),
.B(n_104),
.C(n_105),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_49),
.Y(n_140)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_71),
.B1(n_74),
.B2(n_77),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_65),
.A2(n_71),
.B1(n_77),
.B2(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_66),
.B(n_73),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_67),
.B1(n_87),
.B2(n_88),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_66),
.B(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_77),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_71),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_72),
.A2(n_73),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_72),
.B(n_169),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_73),
.B(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_77),
.A2(n_174),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_77),
.B(n_104),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_77),
.A2(n_142),
.B(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_78),
.B(n_92),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_82),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_85),
.A2(n_91),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_89),
.A2(n_95),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_89),
.B(n_104),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_91),
.B(n_96),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_100),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_97),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_99),
.B(n_123),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_101),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_125),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_117),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_146),
.B(n_226),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_143),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_130),
.B(n_143),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_136),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_131),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_134),
.B(n_136),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_141),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_137),
.B(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_221),
.B(n_225),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_206),
.B(n_220),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_190),
.B(n_205),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_170),
.B(n_189),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_159),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_157),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_152),
.A2(n_153),
.B1(n_157),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B(n_156),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_154),
.A2(n_156),
.B(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_167),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_178),
.B(n_188),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_172),
.B(n_176),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_183),
.B(n_187),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_180),
.B(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_192),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_200),
.C(n_204),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_196),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_197)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_208),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_216),
.C(n_218),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);


endmodule