module fake_jpeg_13539_n_68 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_68);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

BUFx10_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx14_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_30),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_10),
.B(n_13),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_18),
.B(n_13),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_20),
.B(n_17),
.C(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_15),
.B1(n_17),
.B2(n_33),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_27),
.B1(n_18),
.B2(n_26),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_18),
.A3(n_23),
.B1(n_29),
.B2(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_48),
.B(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_47),
.C(n_50),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_48),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_59),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_55),
.B1(n_59),
.B2(n_37),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.B(n_62),
.C(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

OAI31xp33_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_35),
.A3(n_38),
.B(n_32),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_38),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_32),
.B1(n_34),
.B2(n_64),
.Y(n_68)
);


endmodule