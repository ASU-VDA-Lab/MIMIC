module fake_jpeg_6128_n_251 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_42),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_12),
.B1(n_23),
.B2(n_22),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_12),
.B1(n_20),
.B2(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_12),
.B1(n_27),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_55),
.B1(n_13),
.B2(n_19),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_43),
.B(n_38),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_16),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_12),
.B1(n_18),
.B2(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_32),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_31),
.B(n_25),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_44),
.B(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_66),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_67),
.B(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_29),
.B1(n_37),
.B2(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_57),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_29),
.B(n_28),
.C(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_41),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_29),
.Y(n_78)
);

OR2x4_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_29),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_82),
.C(n_84),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_66),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_54),
.B1(n_60),
.B2(n_51),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_72),
.B1(n_70),
.B2(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_63),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_40),
.B(n_47),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_64),
.C(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_104),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_79),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_82),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_85),
.B1(n_94),
.B2(n_96),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_109),
.B(n_90),
.Y(n_119)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_64),
.B(n_76),
.C(n_69),
.D(n_63),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_72),
.C(n_76),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_73),
.C(n_71),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_96),
.C(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_80),
.B(n_79),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_130),
.B(n_132),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_85),
.B1(n_80),
.B2(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_117),
.A2(n_127),
.B1(n_131),
.B2(n_58),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_120),
.C(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_108),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_92),
.B1(n_82),
.B2(n_70),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_94),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_112),
.C(n_113),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_92),
.B(n_86),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_81),
.B1(n_67),
.B2(n_61),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_98),
.B(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_105),
.B1(n_104),
.B2(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_102),
.B(n_97),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_148),
.B(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_147),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_143),
.C(n_34),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_106),
.B1(n_58),
.B2(n_91),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_126),
.B1(n_91),
.B2(n_122),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_126),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_67),
.C(n_81),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_108),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_155),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_154),
.B(n_34),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_153),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_40),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_16),
.B(n_17),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_121),
.B1(n_116),
.B2(n_115),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_28),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_163),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_146),
.B1(n_147),
.B2(n_135),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_132),
.B1(n_119),
.B2(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_132),
.B1(n_143),
.B2(n_139),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_R g164 ( 
.A(n_137),
.B(n_130),
.C(n_124),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_154),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_16),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_41),
.B1(n_23),
.B2(n_22),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_31),
.C(n_25),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_37),
.C(n_36),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_37),
.C(n_36),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_34),
.C(n_36),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_152),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_183),
.C(n_184),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_168),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_149),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_41),
.B1(n_20),
.B2(n_22),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_166),
.B1(n_20),
.B2(n_19),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_34),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_28),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_34),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_160),
.B(n_11),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

NAND4xp25_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_164),
.C(n_161),
.D(n_37),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_199),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_24),
.B(n_21),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_171),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_167),
.B1(n_165),
.B2(n_173),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_202),
.B1(n_34),
.B2(n_1),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_165),
.B1(n_175),
.B2(n_166),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_204),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_24),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_34),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_177),
.C(n_183),
.Y(n_209)
);

OAI322xp33_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_28),
.A3(n_34),
.B1(n_24),
.B2(n_21),
.C1(n_14),
.C2(n_11),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_207),
.A2(n_19),
.B(n_28),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_184),
.B1(n_177),
.B2(n_190),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_209),
.C(n_211),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_213),
.B(n_214),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_0),
.B(n_1),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_212),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_1),
.B(n_2),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_218),
.C(n_3),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_24),
.C(n_21),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_206),
.B1(n_201),
.B2(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_2),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_228),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_215),
.B(n_24),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_229),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_24),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_3),
.C(n_4),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_233),
.C(n_5),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_3),
.B(n_5),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_236),
.A2(n_3),
.B(n_5),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_6),
.B(n_7),
.Y(n_246)
);

OAI321xp33_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_21),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_239)
);

OAI211xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_242),
.B(n_243),
.C(n_235),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_237),
.B(n_234),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_244),
.A2(n_246),
.B1(n_9),
.B2(n_10),
.Y(n_249)
);

AOI321xp33_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_6),
.C(n_8),
.Y(n_248)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_249),
.B(n_245),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_250),
.Y(n_251)
);


endmodule