module real_jpeg_5070_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_22),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_1),
.A2(n_36),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_1),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_1),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_1),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_1),
.A2(n_165),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_1),
.A2(n_261),
.B(n_264),
.C(n_267),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_1),
.B(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_1),
.B(n_55),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_1),
.B(n_75),
.C(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_1),
.B(n_112),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_1),
.B(n_108),
.C(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_1),
.B(n_29),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_78),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_2),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_2),
.A2(n_83),
.B1(n_114),
.B2(n_118),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_2),
.A2(n_83),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_3),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_89),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_3),
.A2(n_89),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_89),
.B1(n_204),
.B2(n_208),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_6),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_6),
.Y(n_275)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_9),
.A2(n_24),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_9),
.A2(n_24),
.B1(n_194),
.B2(n_198),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_9),
.A2(n_24),
.B1(n_178),
.B2(n_273),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_10),
.Y(n_269)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_11),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_12),
.Y(n_400)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_396),
.B(n_398),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_145),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_18),
.B(n_127),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_52),
.C(n_84),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_20),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_20),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_20),
.A2(n_129),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_20),
.B(n_152),
.C(n_192),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_20),
.B(n_242),
.C(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_20),
.A2(n_129),
.B1(n_242),
.B2(n_336),
.Y(n_359)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B1(n_48),
.B2(n_51),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_21),
.A2(n_28),
.B1(n_48),
.B2(n_51),
.Y(n_134)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_28),
.A2(n_48),
.B1(n_51),
.B2(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_28),
.A2(n_48),
.B(n_51),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_31),
.Y(n_142)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_36),
.Y(n_266)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_52),
.A2(n_84),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_52),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_52),
.B(n_134),
.C(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_52),
.A2(n_133),
.B1(n_136),
.B2(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_80),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_53),
.B(n_162),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_68),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_54),
.A2(n_68),
.B1(n_155),
.B2(n_161),
.Y(n_154)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_55),
.A2(n_203),
.B(n_209),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_55),
.B(n_156),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_55),
.A2(n_69),
.B1(n_80),
.B2(n_203),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_59),
.B1(n_62),
.B2(n_66),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_60),
.Y(n_179)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_61),
.Y(n_226)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_65),
.Y(n_186)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_69),
.B(n_162),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_72),
.Y(n_164)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_72),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_72),
.Y(n_299)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_91),
.B1(n_112),
.B2(n_113),
.Y(n_84)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_88),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_91),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_103),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_92),
.A2(n_103),
.B1(n_140),
.B2(n_193),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_92),
.A2(n_103),
.B1(n_140),
.B2(n_193),
.Y(n_242)
);

NAND2x1_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_99),
.Y(n_318)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

AOI22x1_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_103)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_106),
.Y(n_320)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_122),
.B(n_139),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.C(n_135),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_128),
.A2(n_134),
.B1(n_254),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_128),
.Y(n_380)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_134),
.B(n_217),
.C(n_230),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_134),
.A2(n_230),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_134),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_134),
.A2(n_254),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_134),
.B(n_192),
.C(n_346),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_134),
.A2(n_254),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_135),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_136),
.Y(n_385)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_141),
.A2(n_262),
.B(n_265),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_376),
.B(n_393),
.Y(n_146)
);

OAI211xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_276),
.B(n_370),
.C(n_375),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_247),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_149),
.A2(n_247),
.B(n_371),
.C(n_374),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_231),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_150),
.B(n_231),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_200),
.C(n_216),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_151),
.B(n_200),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_190),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_170),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_153),
.A2(n_154),
.B1(n_170),
.B2(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_153),
.A2(n_154),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_153),
.A2(n_154),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_154),
.B(n_271),
.C(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_154),
.B(n_328),
.C(n_330),
.Y(n_341)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_170),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_176),
.B1(n_181),
.B2(n_187),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_172),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_176),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_177),
.A2(n_223),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_177),
.A2(n_223),
.B1(n_272),
.B2(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_178),
.Y(n_287)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_184),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_184),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_191),
.A2(n_192),
.B1(n_228),
.B2(n_297),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_191),
.B(n_297),
.C(n_315),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_191),
.A2(n_192),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_211),
.B2(n_215),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_211),
.Y(n_238)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_215),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_211),
.A2(n_237),
.B(n_238),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_212),
.B(n_223),
.Y(n_321)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_228),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_219),
.A2(n_228),
.B1(n_297),
.B2(n_362),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_219),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_228),
.A2(n_297),
.B1(n_298),
.B2(n_302),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_228),
.Y(n_297)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_245),
.B2(n_246),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_239),
.B1(n_240),
.B2(n_244),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_239),
.B(n_244),
.C(n_246),
.Y(n_392)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_242),
.A2(n_332),
.B1(n_333),
.B2(n_336),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_242),
.Y(n_336)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_243),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_243),
.A2(n_382),
.B1(n_386),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_248),
.B(n_250),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_256),
.C(n_258),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_252),
.B(n_256),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_258),
.B(n_369),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_259),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_270),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_260),
.A2(n_270),
.B1(n_271),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_260),
.Y(n_353)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_270),
.A2(n_271),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_271),
.B(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_292),
.Y(n_293)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_355),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_340),
.B(n_354),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_325),
.B(n_339),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_312),
.B(n_324),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_304),
.B(n_311),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_294),
.B(n_303),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_291),
.B(n_293),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_289),
.A2(n_295),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_296),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_295),
.B(n_334),
.C(n_336),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_302),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_298),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_310),
.Y(n_311)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_314),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_321),
.B2(n_322),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_322),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_338),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_338),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_330),
.B1(n_331),
.B2(n_337),
.Y(n_326)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_342),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_348),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_350),
.C(n_351),
.Y(n_364)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_346),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2x1_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_365),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_364),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_364),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_363),
.C(n_367),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_365),
.A2(n_372),
.B(n_373),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_368),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_388),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_377),
.A2(n_394),
.B(n_395),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_381),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_386),
.C(n_387),
.Y(n_381)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_387),
.B(n_390),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_392),
.Y(n_394)
);

INVx8_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_397),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);


endmodule