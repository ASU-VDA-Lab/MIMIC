module fake_jpeg_6930_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_219;
wire n_70;
wire n_130;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_37),
.Y(n_91)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_43),
.Y(n_65)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_17),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_54),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

OR2x4_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_0),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_27),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_53),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_23),
.B1(n_20),
.B2(n_33),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_59),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_93),
.B1(n_2),
.B2(n_5),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_22),
.B1(n_26),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_68),
.B1(n_73),
.B2(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_70),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_23),
.B1(n_28),
.B2(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_31),
.B1(n_28),
.B2(n_32),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_13),
.B(n_8),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_57),
.B1(n_42),
.B2(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_74),
.B(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_40),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_82),
.B(n_85),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_43),
.B(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_49),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_36),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_41),
.A2(n_36),
.B1(n_30),
.B2(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_36),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_104),
.Y(n_141)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_99),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_103),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_113),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

BUFx6f_ASAP7_75t_SL g111 ( 
.A(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_6),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_6),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_6),
.Y(n_116)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_96),
.B1(n_124),
.B2(n_94),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_61),
.B(n_83),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_75),
.B(n_84),
.Y(n_140)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_72),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_79),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_132),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_137),
.B1(n_143),
.B2(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_97),
.B(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_71),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_91),
.C(n_83),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_10),
.C(n_11),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_145),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_74),
.B1(n_75),
.B2(n_86),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_98),
.B1(n_118),
.B2(n_69),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_84),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_87),
.B(n_11),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_56),
.B1(n_69),
.B2(n_90),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_151),
.A2(n_122),
.B(n_111),
.C(n_102),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_119),
.B1(n_113),
.B2(n_105),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_158),
.B1(n_164),
.B2(n_165),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_166),
.B(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_160),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_123),
.B1(n_125),
.B2(n_101),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_120),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_7),
.C(n_8),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_135),
.C(n_150),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_118),
.B1(n_70),
.B2(n_90),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_87),
.B(n_99),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_132),
.C(n_129),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_133),
.B(n_11),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_172),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_151),
.B(n_143),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_173),
.B(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_136),
.B(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_144),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_177),
.A2(n_178),
.B1(n_168),
.B2(n_155),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_185),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_181),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_146),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_153),
.C(n_162),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_189),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_133),
.C(n_146),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_161),
.B1(n_154),
.B2(n_157),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_167),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_198),
.C(n_204),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_177),
.A3(n_181),
.B1(n_188),
.B2(n_186),
.C1(n_156),
.C2(n_191),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_191),
.C(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_201),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_162),
.A3(n_153),
.B1(n_165),
.B2(n_155),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_169),
.C(n_127),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_192),
.C(n_184),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_201),
.C(n_214),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_214),
.C(n_205),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_182),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_195),
.B(n_202),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_199),
.B1(n_195),
.B2(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_198),
.A2(n_176),
.B1(n_190),
.B2(n_131),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_216),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_204),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_220),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_221),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_224),
.B(n_208),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_203),
.C(n_149),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_207),
.B(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_226),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_216),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_128),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_228),
.B(n_130),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_130),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_229),
.C(n_228),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_234),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_237),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_239),
.A2(n_235),
.B(n_238),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_240),
.B(n_237),
.CI(n_236),
.CON(n_241),
.SN(n_241)
);


endmodule