module fake_netlist_6_2215_n_2779 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_797, n_666, n_371, n_795, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_808, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_788, n_325, n_767, n_804, n_329, n_464, n_600, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_2779);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_808;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_788;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2779;

wire n_992;
wire n_2542;
wire n_1671;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_822;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_1591;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_2641;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2345;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2319;
wire n_2519;
wire n_825;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_890;
wire n_2377;
wire n_2178;
wire n_950;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_2767;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_1992;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_2289;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2100;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_1593;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_845;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_1397;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_1900;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1650;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_876;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_1542;
wire n_2587;
wire n_875;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_946;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_2743;
wire n_1973;
wire n_2267;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_800),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_610),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_326),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_359),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_194),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_740),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_69),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_104),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_377),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_731),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_734),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_376),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_737),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_709),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_43),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_84),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_217),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_710),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_192),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_699),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_795),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_425),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_113),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_387),
.Y(n_833)
);

CKINVDCx16_ASAP7_75t_R g834 ( 
.A(n_504),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_331),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_481),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_311),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_783),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_257),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_335),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_729),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_803),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_114),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_507),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_706),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_778),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_135),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_764),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_391),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_672),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_419),
.Y(n_851)
);

CKINVDCx16_ASAP7_75t_R g852 ( 
.A(n_223),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_307),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_619),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_473),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_633),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_773),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_275),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_143),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_335),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_782),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_518),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_350),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_741),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_714),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_102),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_704),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_546),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_53),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_751),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_655),
.Y(n_871)
);

INVxp33_ASAP7_75t_R g872 ( 
.A(n_723),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_485),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_293),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_692),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_725),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_305),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_131),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_808),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_801),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_496),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_269),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_762),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_727),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_562),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_766),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_499),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_152),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_184),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_747),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_785),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_749),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_13),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_302),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_541),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_193),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_744),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_334),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_776),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_739),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_407),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_682),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_746),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_109),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_279),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_6),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_533),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_255),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_799),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_533),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_332),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_428),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_806),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_631),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_598),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_796),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_189),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_618),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_777),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_275),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_417),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_541),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_461),
.Y(n_923)
);

BUFx2_ASAP7_75t_SL g924 ( 
.A(n_56),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_3),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_71),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_605),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_144),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_65),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_186),
.Y(n_930)
);

CKINVDCx14_ASAP7_75t_R g931 ( 
.A(n_798),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_1),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_715),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_257),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_382),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_11),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_105),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_745),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_802),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_212),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_790),
.Y(n_941)
);

BUFx10_ASAP7_75t_L g942 ( 
.A(n_465),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_91),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_59),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_285),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_331),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_187),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_68),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_233),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_404),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_807),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_43),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_641),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_805),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_417),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_647),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_538),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_213),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_46),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_694),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_732),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_466),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_218),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_395),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_357),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_219),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_728),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_488),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_530),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_718),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_791),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_406),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_752),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_322),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_769),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_115),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_388),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_753),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_761),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_305),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_240),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_711),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_121),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_14),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_9),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_253),
.Y(n_986)
);

BUFx2_ASAP7_75t_SL g987 ( 
.A(n_804),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_57),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_788),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_701),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_134),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_579),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_441),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_794),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_722),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_419),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_736),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_754),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_2),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_464),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_263),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_569),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_569),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_757),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_772),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_330),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_684),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_74),
.Y(n_1008)
);

BUFx10_ASAP7_75t_L g1009 ( 
.A(n_68),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_779),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_64),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_56),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_246),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_255),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_386),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_298),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_500),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_742),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_534),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_32),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_792),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_427),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_294),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_112),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_292),
.Y(n_1025)
);

CKINVDCx14_ASAP7_75t_R g1026 ( 
.A(n_448),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_748),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_583),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_750),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_730),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_96),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_789),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_79),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_85),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_705),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_675),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_719),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_144),
.Y(n_1038)
);

BUFx10_ASAP7_75t_L g1039 ( 
.A(n_767),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_797),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_202),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_743),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_267),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_696),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_258),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_465),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_775),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_693),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_770),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_613),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_708),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_716),
.Y(n_1052)
);

BUFx10_ASAP7_75t_L g1053 ( 
.A(n_566),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_195),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_77),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_36),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_676),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_58),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_106),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_691),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_765),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_253),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_662),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_758),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_483),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_774),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_707),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_3),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_179),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_96),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_486),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_114),
.Y(n_1072)
);

CKINVDCx14_ASAP7_75t_R g1073 ( 
.A(n_439),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_759),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_495),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_488),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_446),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_784),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_733),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_763),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_89),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_380),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_167),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_724),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_500),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_222),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_219),
.Y(n_1087)
);

BUFx2_ASAP7_75t_SL g1088 ( 
.A(n_213),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_300),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_316),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_712),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_532),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_548),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_720),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_449),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_395),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_627),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_621),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_307),
.Y(n_1099)
);

CKINVDCx14_ASAP7_75t_R g1100 ( 
.A(n_449),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_193),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_781),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_366),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_786),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_178),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_436),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_612),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_717),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_738),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_609),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_467),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_108),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_726),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_780),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_793),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_426),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_713),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_458),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_243),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_345),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_760),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_735),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_544),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_768),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_401),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_771),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_148),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_189),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_362),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_322),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_279),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_787),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_173),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_473),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_755),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_220),
.Y(n_1136)
);

BUFx10_ASAP7_75t_L g1137 ( 
.A(n_721),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_702),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_614),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_50),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_285),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_61),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_756),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_371),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_247),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_122),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_565),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_916),
.B(n_1),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1026),
.B(n_2),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1073),
.B(n_0),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_917),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_917),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1100),
.B(n_0),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_933),
.B(n_5),
.Y(n_1154)
);

BUFx12f_ASAP7_75t_L g1155 ( 
.A(n_942),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_917),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1039),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_947),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_863),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_856),
.B(n_1030),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_879),
.B(n_4),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_864),
.B(n_4),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_971),
.B(n_6),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_844),
.B(n_5),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_947),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_979),
.B(n_7),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_972),
.B(n_7),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_982),
.B(n_9),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_845),
.B(n_10),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_884),
.B(n_8),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_910),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_931),
.B(n_8),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1027),
.B(n_10),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_900),
.B(n_12),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1057),
.B(n_11),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_942),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_947),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_811),
.B(n_823),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_842),
.B(n_12),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_953),
.B(n_13),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_955),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1149),
.A2(n_834),
.B1(n_852),
.B2(n_829),
.Y(n_1182)
);

AO22x2_ASAP7_75t_L g1183 ( 
.A1(n_1164),
.A2(n_1167),
.B1(n_1166),
.B2(n_1153),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1152),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1151),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1171),
.B(n_1141),
.Y(n_1186)
);

OAI22xp33_ASAP7_75t_SL g1187 ( 
.A1(n_1150),
.A2(n_934),
.B1(n_1083),
.B2(n_922),
.Y(n_1187)
);

NAND3x1_ASAP7_75t_L g1188 ( 
.A(n_1148),
.B(n_824),
.C(n_814),
.Y(n_1188)
);

CKINVDCx6p67_ASAP7_75t_R g1189 ( 
.A(n_1155),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1180),
.A2(n_830),
.B1(n_871),
.B2(n_822),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1171),
.B(n_985),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1172),
.A2(n_956),
.B1(n_1032),
.B2(n_903),
.Y(n_1192)
);

AO22x2_ASAP7_75t_L g1193 ( 
.A1(n_1166),
.A2(n_1179),
.B1(n_988),
.B2(n_1043),
.Y(n_1193)
);

OAI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1176),
.A2(n_1130),
.B1(n_888),
.B2(n_936),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1173),
.A2(n_1129),
.B1(n_828),
.B2(n_1001),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1169),
.A2(n_1064),
.B1(n_1102),
.B2(n_1040),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1160),
.B(n_1042),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1159),
.B(n_993),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1174),
.A2(n_812),
.B1(n_816),
.B2(n_813),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1157),
.B(n_1071),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1175),
.A2(n_818),
.B1(n_821),
.B2(n_817),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1161),
.A2(n_836),
.B1(n_837),
.B2(n_835),
.Y(n_1202)
);

OAI22xp33_ASAP7_75t_R g1203 ( 
.A1(n_1154),
.A2(n_831),
.B1(n_832),
.B2(n_825),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1163),
.A2(n_840),
.B1(n_843),
.B2(n_839),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1178),
.B(n_1137),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1178),
.B(n_1137),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1151),
.B(n_1039),
.Y(n_1207)
);

AO22x2_ASAP7_75t_L g1208 ( 
.A1(n_1179),
.A2(n_1088),
.B1(n_924),
.B2(n_851),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1168),
.A2(n_855),
.B1(n_858),
.B2(n_847),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1156),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1156),
.Y(n_1211)
);

AO22x2_ASAP7_75t_L g1212 ( 
.A1(n_1162),
.A2(n_853),
.B1(n_860),
.B2(n_849),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1165),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_SL g1214 ( 
.A(n_1158),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1184),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1210),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1189),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1211),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1213),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1197),
.B(n_1091),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1186),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1205),
.A2(n_1170),
.B(n_867),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1185),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1191),
.B(n_1177),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1200),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1198),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1207),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_1206),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1212),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1212),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1183),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1183),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1193),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1204),
.B(n_1181),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1193),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1208),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1208),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1214),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1188),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1209),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1199),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1203),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1187),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1196),
.B(n_1177),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1201),
.B(n_1165),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1202),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1195),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1192),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1194),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1182),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1190),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1210),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1197),
.B(n_872),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1210),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1197),
.B(n_1132),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1210),
.Y(n_1256)
);

XOR2xp5_ASAP7_75t_L g1257 ( 
.A(n_1190),
.B(n_810),
.Y(n_1257)
);

NOR2xp67_ASAP7_75t_L g1258 ( 
.A(n_1196),
.B(n_815),
.Y(n_1258)
);

XOR2xp5_ASAP7_75t_L g1259 ( 
.A(n_1190),
.B(n_819),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1197),
.B(n_1115),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1210),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1210),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1254),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1215),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1225),
.B(n_1221),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1222),
.A2(n_875),
.B(n_861),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1255),
.B(n_880),
.Y(n_1267)
);

AND2x2_ASAP7_75t_SL g1268 ( 
.A(n_1253),
.B(n_955),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1260),
.B(n_883),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1215),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1224),
.B(n_1227),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1228),
.B(n_1009),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1216),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1220),
.B(n_859),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1216),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1226),
.B(n_886),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1254),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1244),
.B(n_1009),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1218),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1217),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1254),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1251),
.B(n_873),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1257),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1229),
.B(n_891),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1234),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1240),
.B(n_1241),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1246),
.B(n_897),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1234),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1258),
.B(n_820),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1219),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1252),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1245),
.B(n_1233),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1249),
.B(n_1053),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1256),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1250),
.B(n_1248),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1259),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1235),
.B(n_1053),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1242),
.B(n_893),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1231),
.B(n_899),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1261),
.Y(n_1300)
);

XNOR2xp5_ASAP7_75t_L g1301 ( 
.A(n_1239),
.B(n_930),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1262),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1223),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1247),
.B(n_945),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1232),
.B(n_902),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1230),
.B(n_913),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1236),
.B(n_918),
.Y(n_1307)
);

AND2x2_ASAP7_75t_SL g1308 ( 
.A(n_1243),
.B(n_1237),
.Y(n_1308)
);

INVxp67_ASAP7_75t_L g1309 ( 
.A(n_1238),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1224),
.B(n_869),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1255),
.B(n_827),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1224),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1255),
.B(n_938),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1225),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1215),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1215),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1255),
.B(n_941),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1215),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1217),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1225),
.B(n_957),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_R g1321 ( 
.A(n_1217),
.B(n_838),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1255),
.B(n_954),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1215),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1255),
.B(n_862),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1225),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1215),
.Y(n_1326)
);

CKINVDCx8_ASAP7_75t_R g1327 ( 
.A(n_1217),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1224),
.B(n_967),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1225),
.Y(n_1329)
);

AND2x2_ASAP7_75t_SL g1330 ( 
.A(n_1253),
.B(n_955),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1224),
.B(n_970),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1224),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1222),
.A2(n_1007),
.B(n_995),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1225),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1224),
.B(n_1010),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1225),
.B(n_964),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1215),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1254),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1215),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1224),
.B(n_1047),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1255),
.B(n_1049),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1215),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1225),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1225),
.Y(n_1344)
);

INVx4_ASAP7_75t_L g1345 ( 
.A(n_1224),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1215),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1215),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1255),
.A2(n_846),
.B1(n_848),
.B2(n_841),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1225),
.B(n_981),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1225),
.B(n_1019),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1215),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1254),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1215),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1225),
.B(n_1046),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1215),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1224),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1225),
.B(n_1077),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1215),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1255),
.B(n_1060),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1215),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1255),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1225),
.B(n_1082),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1217),
.Y(n_1363)
);

AND2x6_ASAP7_75t_L g1364 ( 
.A(n_1231),
.B(n_1067),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1215),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1225),
.B(n_1092),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1225),
.B(n_1093),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1277),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1315),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1326),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1277),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1314),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_1325),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1334),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1361),
.B(n_866),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1338),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1337),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1324),
.B(n_1080),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1329),
.B(n_1144),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1339),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1274),
.B(n_1094),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1338),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1284),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1312),
.B(n_877),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1332),
.B(n_1271),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1267),
.B(n_1098),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1345),
.B(n_850),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1343),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1356),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1342),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1347),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1351),
.Y(n_1392)
);

NAND2x1p5_ASAP7_75t_L g1393 ( 
.A(n_1265),
.B(n_850),
.Y(n_1393)
);

OR2x6_ASAP7_75t_L g1394 ( 
.A(n_1288),
.B(n_1285),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1264),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1271),
.B(n_882),
.Y(n_1396)
);

NAND2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1263),
.B(n_850),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1310),
.B(n_1284),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1353),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1278),
.B(n_868),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1320),
.B(n_1147),
.Y(n_1401)
);

AND2x6_ASAP7_75t_L g1402 ( 
.A(n_1295),
.B(n_889),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1344),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1352),
.B(n_1281),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1336),
.B(n_1128),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1269),
.B(n_1117),
.Y(n_1406)
);

BUFx4f_ASAP7_75t_L g1407 ( 
.A(n_1364),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1270),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1305),
.B(n_896),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1313),
.B(n_1122),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1316),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1360),
.Y(n_1412)
);

NAND2x1p5_ASAP7_75t_L g1413 ( 
.A(n_1318),
.B(n_989),
.Y(n_1413)
);

AND2x2_ASAP7_75t_SL g1414 ( 
.A(n_1268),
.B(n_977),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1305),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1330),
.B(n_1282),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1303),
.B(n_908),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1317),
.B(n_1322),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1293),
.B(n_1272),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1323),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1341),
.B(n_1143),
.Y(n_1421)
);

NAND2x1_ASAP7_75t_SL g1422 ( 
.A(n_1349),
.B(n_911),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1350),
.B(n_881),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1346),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1354),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1357),
.Y(n_1426)
);

AND2x6_ASAP7_75t_L g1427 ( 
.A(n_1297),
.B(n_912),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1280),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1319),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1286),
.B(n_1127),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1363),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1365),
.Y(n_1432)
);

AND2x2_ASAP7_75t_SL g1433 ( 
.A(n_1367),
.B(n_977),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_L g1434 ( 
.A(n_1292),
.B(n_987),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1366),
.B(n_885),
.Y(n_1435)
);

AND2x2_ASAP7_75t_SL g1436 ( 
.A(n_1362),
.B(n_977),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1328),
.B(n_940),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1364),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1328),
.B(n_1331),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1359),
.B(n_854),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1266),
.B(n_857),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1304),
.B(n_887),
.Y(n_1442)
);

CKINVDCx6p67_ASAP7_75t_R g1443 ( 
.A(n_1308),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1333),
.B(n_865),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1355),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1358),
.B(n_870),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1273),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1298),
.B(n_894),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1296),
.B(n_895),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1331),
.B(n_898),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1287),
.B(n_876),
.Y(n_1451)
);

AND2x6_ASAP7_75t_L g1452 ( 
.A(n_1307),
.B(n_949),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1275),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1335),
.B(n_950),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1335),
.B(n_958),
.Y(n_1455)
);

BUFx8_ASAP7_75t_L g1456 ( 
.A(n_1307),
.Y(n_1456)
);

INVxp67_ASAP7_75t_SL g1457 ( 
.A(n_1279),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1311),
.B(n_890),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1291),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1348),
.B(n_901),
.Y(n_1460)
);

INVx5_ASAP7_75t_L g1461 ( 
.A(n_1364),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1294),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_SL g1463 ( 
.A(n_1327),
.B(n_892),
.Y(n_1463)
);

BUFx4f_ASAP7_75t_L g1464 ( 
.A(n_1340),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1309),
.B(n_965),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1340),
.B(n_904),
.Y(n_1466)
);

NAND2x1_ASAP7_75t_SL g1467 ( 
.A(n_1290),
.B(n_976),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1300),
.Y(n_1468)
);

INVx6_ASAP7_75t_L g1469 ( 
.A(n_1321),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1302),
.B(n_996),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1276),
.B(n_909),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1299),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1306),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1289),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1283),
.B(n_999),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1301),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1301),
.Y(n_1477)
);

OR2x2_ASAP7_75t_SL g1478 ( 
.A(n_1314),
.B(n_826),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1264),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1314),
.Y(n_1480)
);

NAND2x1p5_ASAP7_75t_L g1481 ( 
.A(n_1312),
.B(n_989),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1361),
.B(n_905),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1314),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1264),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1315),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1361),
.B(n_906),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1315),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1361),
.B(n_907),
.Y(n_1488)
);

AND2x6_ASAP7_75t_L g1489 ( 
.A(n_1278),
.B(n_1015),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1361),
.B(n_915),
.Y(n_1490)
);

NOR2xp67_ASAP7_75t_L g1491 ( 
.A(n_1280),
.B(n_914),
.Y(n_1491)
);

NAND2x1_ASAP7_75t_SL g1492 ( 
.A(n_1278),
.B(n_1016),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1312),
.B(n_1017),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1361),
.B(n_920),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1361),
.B(n_919),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1315),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1361),
.B(n_921),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1264),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1277),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1361),
.B(n_923),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1277),
.Y(n_1501)
);

BUFx4f_ASAP7_75t_L g1502 ( 
.A(n_1364),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1315),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1280),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1361),
.B(n_927),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1264),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_1329),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1361),
.B(n_925),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1264),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1361),
.B(n_926),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1288),
.B(n_1020),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1312),
.B(n_1022),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1361),
.B(n_928),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1329),
.Y(n_1514)
);

AND2x2_ASAP7_75t_SL g1515 ( 
.A(n_1268),
.B(n_1085),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1312),
.B(n_1033),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1264),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1329),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_SL g1519 ( 
.A(n_1327),
.B(n_939),
.Y(n_1519)
);

AND2x6_ASAP7_75t_L g1520 ( 
.A(n_1278),
.B(n_1034),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1312),
.B(n_1041),
.Y(n_1521)
);

CKINVDCx6p67_ASAP7_75t_R g1522 ( 
.A(n_1431),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

BUFx12f_ASAP7_75t_L g1524 ( 
.A(n_1456),
.Y(n_1524)
);

BUFx2_ASAP7_75t_SL g1525 ( 
.A(n_1429),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1419),
.B(n_929),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1453),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1395),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1408),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1472),
.B(n_951),
.Y(n_1530)
);

INVx8_ASAP7_75t_L g1531 ( 
.A(n_1371),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1428),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1469),
.Y(n_1533)
);

INVx5_ASAP7_75t_L g1534 ( 
.A(n_1504),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1403),
.Y(n_1535)
);

BUFx5_ASAP7_75t_L g1536 ( 
.A(n_1411),
.Y(n_1536)
);

INVx4_ASAP7_75t_L g1537 ( 
.A(n_1371),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1376),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1514),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1420),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1424),
.Y(n_1541)
);

INVx5_ASAP7_75t_L g1542 ( 
.A(n_1402),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1376),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1382),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1430),
.B(n_935),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1374),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1372),
.B(n_960),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1445),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_943),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1388),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1479),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1484),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1443),
.Y(n_1553)
);

INVx5_ASAP7_75t_SL g1554 ( 
.A(n_1511),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1498),
.Y(n_1555)
);

BUFx12f_ASAP7_75t_L g1556 ( 
.A(n_1478),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1418),
.B(n_961),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1369),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1382),
.Y(n_1559)
);

BUFx8_ASAP7_75t_L g1560 ( 
.A(n_1475),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_1425),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1394),
.B(n_1439),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1521),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1506),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1499),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1509),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1499),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1501),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1501),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1415),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1517),
.Y(n_1571)
);

BUFx4_ASAP7_75t_SL g1572 ( 
.A(n_1465),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1384),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1415),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1373),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1370),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_SL g1577 ( 
.A(n_1416),
.B(n_973),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1468),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1480),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1377),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1473),
.B(n_975),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1380),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1375),
.B(n_946),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1389),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1398),
.B(n_1056),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1483),
.B(n_948),
.Y(n_1586)
);

BUFx12f_ASAP7_75t_L g1587 ( 
.A(n_1426),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1493),
.Y(n_1588)
);

INVx8_ASAP7_75t_L g1589 ( 
.A(n_1452),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1379),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1449),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1422),
.Y(n_1592)
);

INVx6_ASAP7_75t_SL g1593 ( 
.A(n_1512),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1476),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1492),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1383),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1477),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1390),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1516),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1396),
.Y(n_1600)
);

BUFx10_ASAP7_75t_L g1601 ( 
.A(n_1486),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1385),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1368),
.Y(n_1603)
);

BUFx12f_ASAP7_75t_L g1604 ( 
.A(n_1409),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1495),
.Y(n_1605)
);

INVx3_ASAP7_75t_SL g1606 ( 
.A(n_1417),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1383),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1467),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1470),
.Y(n_1609)
);

INVx3_ASAP7_75t_SL g1610 ( 
.A(n_1437),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1454),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1402),
.Y(n_1612)
);

CKINVDCx16_ASAP7_75t_R g1613 ( 
.A(n_1463),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1391),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1392),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1455),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1399),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1412),
.Y(n_1618)
);

NAND2x1_ASAP7_75t_L g1619 ( 
.A(n_1432),
.B(n_989),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1490),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1472),
.B(n_978),
.Y(n_1621)
);

INVx8_ASAP7_75t_L g1622 ( 
.A(n_1452),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1464),
.Y(n_1623)
);

INVx5_ASAP7_75t_L g1624 ( 
.A(n_1427),
.Y(n_1624)
);

BUFx2_ASAP7_75t_R g1625 ( 
.A(n_1438),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1427),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1404),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1447),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1460),
.A2(n_1138),
.B1(n_1139),
.B2(n_1135),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1485),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1487),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1407),
.Y(n_1632)
);

NAND2x1p5_ASAP7_75t_L g1633 ( 
.A(n_1461),
.B(n_1085),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1459),
.B(n_1068),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1401),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1457),
.Y(n_1636)
);

CKINVDCx6p67_ASAP7_75t_R g1637 ( 
.A(n_1461),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1489),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1502),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1545),
.A2(n_1414),
.B1(n_1515),
.B2(n_1378),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1578),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1635),
.A2(n_1433),
.B1(n_1436),
.B2(n_1381),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1528),
.Y(n_1643)
);

INVx6_ASAP7_75t_L g1644 ( 
.A(n_1534),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1539),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1529),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1523),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1561),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1613),
.A2(n_1520),
.B1(n_1489),
.B2(n_1435),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1540),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1541),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1550),
.Y(n_1652)
);

BUFx2_ASAP7_75t_SL g1653 ( 
.A(n_1534),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1577),
.A2(n_1520),
.B1(n_1519),
.B2(n_1494),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1548),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1533),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1551),
.Y(n_1657)
);

BUFx8_ASAP7_75t_L g1658 ( 
.A(n_1524),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1605),
.A2(n_1508),
.B1(n_1510),
.B2(n_1448),
.Y(n_1659)
);

INVx5_ASAP7_75t_L g1660 ( 
.A(n_1531),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1552),
.Y(n_1661)
);

BUFx12f_ASAP7_75t_L g1662 ( 
.A(n_1560),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1555),
.Y(n_1663)
);

BUFx4f_ASAP7_75t_SL g1664 ( 
.A(n_1587),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_SL g1665 ( 
.A1(n_1601),
.A2(n_1442),
.B1(n_1400),
.B2(n_1482),
.Y(n_1665)
);

CKINVDCx6p67_ASAP7_75t_R g1666 ( 
.A(n_1624),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_SL g1667 ( 
.A1(n_1591),
.A2(n_1488),
.B1(n_1500),
.B2(n_1497),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1620),
.A2(n_1441),
.B1(n_1444),
.B2(n_1450),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1564),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1583),
.A2(n_1466),
.B1(n_1434),
.B2(n_1474),
.Y(n_1670)
);

CKINVDCx11_ASAP7_75t_R g1671 ( 
.A(n_1522),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1566),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1595),
.A2(n_1526),
.B1(n_1592),
.B2(n_1629),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1571),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1636),
.A2(n_1505),
.B1(n_1440),
.B2(n_1451),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1590),
.A2(n_1423),
.B1(n_1405),
.B2(n_1513),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1544),
.Y(n_1677)
);

CKINVDCx6p67_ASAP7_75t_R g1678 ( 
.A(n_1624),
.Y(n_1678)
);

NAND2x1p5_ASAP7_75t_L g1679 ( 
.A(n_1535),
.B(n_1496),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1634),
.A2(n_1462),
.B1(n_1503),
.B2(n_1406),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1623),
.Y(n_1681)
);

CKINVDCx11_ASAP7_75t_R g1682 ( 
.A(n_1610),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1544),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1575),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1549),
.B(n_1491),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1557),
.A2(n_1471),
.B1(n_1458),
.B2(n_1446),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1527),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1558),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_SL g1689 ( 
.A1(n_1599),
.A2(n_1393),
.B(n_1410),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1594),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1576),
.Y(n_1691)
);

NAND2x1p5_ASAP7_75t_L g1692 ( 
.A(n_1584),
.B(n_1386),
.Y(n_1692)
);

INVx6_ASAP7_75t_L g1693 ( 
.A(n_1565),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1580),
.Y(n_1694)
);

INVx6_ASAP7_75t_L g1695 ( 
.A(n_1565),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1598),
.A2(n_1421),
.B1(n_1387),
.B2(n_1481),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1614),
.Y(n_1697)
);

INVx8_ASAP7_75t_L g1698 ( 
.A(n_1589),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1579),
.Y(n_1699)
);

CKINVDCx11_ASAP7_75t_R g1700 ( 
.A(n_1604),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1538),
.Y(n_1701)
);

CKINVDCx11_ASAP7_75t_R g1702 ( 
.A(n_1606),
.Y(n_1702)
);

BUFx4f_ASAP7_75t_SL g1703 ( 
.A(n_1593),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1615),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1617),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1628),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1608),
.A2(n_1413),
.B1(n_1397),
.B2(n_1145),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1630),
.A2(n_1076),
.B(n_1072),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1582),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1556),
.A2(n_1581),
.B1(n_1597),
.B2(n_1586),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1618),
.A2(n_994),
.B1(n_997),
.B2(n_990),
.Y(n_1711)
);

CKINVDCx20_ASAP7_75t_R g1712 ( 
.A(n_1525),
.Y(n_1712)
);

BUFx2_ASAP7_75t_SL g1713 ( 
.A(n_1537),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1631),
.A2(n_1546),
.B1(n_1621),
.B2(n_1627),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1602),
.A2(n_1004),
.B1(n_1005),
.B2(n_998),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1585),
.A2(n_1131),
.B1(n_1133),
.B2(n_1125),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1543),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_1532),
.Y(n_1718)
);

CKINVDCx11_ASAP7_75t_R g1719 ( 
.A(n_1632),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1553),
.Y(n_1720)
);

OAI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1542),
.A2(n_959),
.B1(n_962),
.B2(n_952),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1563),
.A2(n_1140),
.B1(n_1146),
.B2(n_1136),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1536),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1536),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1637),
.Y(n_1725)
);

BUFx2_ASAP7_75t_SL g1726 ( 
.A(n_1568),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1536),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1572),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1619),
.Y(n_1729)
);

AO22x1_ASAP7_75t_L g1730 ( 
.A1(n_1542),
.A2(n_968),
.B1(n_969),
.B2(n_963),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1607),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1569),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1570),
.Y(n_1733)
);

CKINVDCx20_ASAP7_75t_R g1734 ( 
.A(n_1638),
.Y(n_1734)
);

INVx4_ASAP7_75t_L g1735 ( 
.A(n_1570),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1603),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_SL g1737 ( 
.A1(n_1609),
.A2(n_980),
.B1(n_983),
.B2(n_974),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1562),
.A2(n_1530),
.B1(n_1625),
.B2(n_1547),
.Y(n_1738)
);

INVx4_ASAP7_75t_L g1739 ( 
.A(n_1574),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1611),
.A2(n_1086),
.B1(n_1087),
.B2(n_1081),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1559),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1616),
.A2(n_1095),
.B1(n_1099),
.B2(n_1089),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1567),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1574),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1632),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1639),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1573),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1588),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1626),
.A2(n_1112),
.B(n_1111),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1612),
.A2(n_1021),
.B1(n_1029),
.B2(n_1018),
.Y(n_1750)
);

BUFx8_ASAP7_75t_L g1751 ( 
.A(n_1639),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1554),
.A2(n_986),
.B1(n_991),
.B2(n_984),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1600),
.A2(n_1036),
.B1(n_1037),
.B2(n_1035),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1633),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1596),
.A2(n_1048),
.B1(n_1050),
.B2(n_1044),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1622),
.A2(n_1124),
.B1(n_1126),
.B2(n_1121),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1590),
.B(n_992),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1578),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1578),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_SL g1760 ( 
.A1(n_1545),
.A2(n_1002),
.B1(n_1003),
.B2(n_1000),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1545),
.A2(n_1052),
.B1(n_1061),
.B2(n_1051),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1531),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1544),
.Y(n_1763)
);

BUFx12f_ASAP7_75t_L g1764 ( 
.A(n_1524),
.Y(n_1764)
);

BUFx3_ASAP7_75t_L g1765 ( 
.A(n_1531),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1578),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1646),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1685),
.A2(n_1008),
.B1(n_1011),
.B2(n_1006),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1640),
.A2(n_1013),
.B1(n_1024),
.B2(n_1012),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1651),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1659),
.A2(n_1038),
.B1(n_1045),
.B2(n_1025),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1642),
.A2(n_1059),
.B1(n_1062),
.B2(n_1055),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1654),
.A2(n_1649),
.B(n_1665),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1661),
.Y(n_1774)
);

OAI21xp33_ASAP7_75t_L g1775 ( 
.A1(n_1760),
.A2(n_1069),
.B(n_1065),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1684),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1667),
.A2(n_1066),
.B1(n_1074),
.B2(n_1063),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1645),
.B(n_1078),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1676),
.A2(n_1085),
.B1(n_1090),
.B2(n_1075),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1673),
.A2(n_1101),
.B1(n_1103),
.B2(n_1096),
.Y(n_1780)
);

OAI21xp33_ASAP7_75t_L g1781 ( 
.A1(n_1668),
.A2(n_1106),
.B(n_1105),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1761),
.A2(n_1118),
.B1(n_1119),
.B2(n_1116),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1670),
.A2(n_1123),
.B1(n_1120),
.B2(n_874),
.Y(n_1783)
);

OAI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1689),
.A2(n_878),
.B1(n_932),
.B2(n_833),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1686),
.A2(n_944),
.B1(n_966),
.B2(n_937),
.Y(n_1785)
);

OAI21xp33_ASAP7_75t_L g1786 ( 
.A1(n_1740),
.A2(n_1142),
.B(n_1134),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1699),
.B(n_1079),
.Y(n_1787)
);

OAI21xp33_ASAP7_75t_L g1788 ( 
.A1(n_1742),
.A2(n_1023),
.B(n_1014),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_SL g1789 ( 
.A1(n_1738),
.A2(n_1031),
.B1(n_1054),
.B2(n_1028),
.Y(n_1789)
);

BUFx4f_ASAP7_75t_SL g1790 ( 
.A(n_1764),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1744),
.B(n_606),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1660),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1712),
.A2(n_1070),
.B1(n_1058),
.B2(n_1084),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1672),
.B(n_1097),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1647),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1710),
.A2(n_1107),
.B1(n_1108),
.B2(n_1104),
.Y(n_1796)
);

INVxp67_ASAP7_75t_SL g1797 ( 
.A(n_1758),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1675),
.A2(n_1110),
.B1(n_1113),
.B2(n_1109),
.Y(n_1798)
);

AOI222xp33_ASAP7_75t_L g1799 ( 
.A1(n_1722),
.A2(n_1114),
.B1(n_16),
.B2(n_18),
.C1(n_19),
.C2(n_15),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_SL g1800 ( 
.A1(n_1653),
.A2(n_22),
.B1(n_30),
.B2(n_14),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1648),
.B(n_607),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_SL g1802 ( 
.A1(n_1690),
.A2(n_1714),
.B1(n_1734),
.B2(n_1720),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1680),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1752),
.A2(n_19),
.B(n_18),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1759),
.Y(n_1805)
);

OAI21xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1737),
.A2(n_21),
.B(n_20),
.Y(n_1806)
);

CKINVDCx20_ASAP7_75t_R g1807 ( 
.A(n_1671),
.Y(n_1807)
);

OAI222xp33_ASAP7_75t_L g1808 ( 
.A1(n_1757),
.A2(n_21),
.B1(n_23),
.B2(n_17),
.C1(n_20),
.C2(n_22),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1687),
.B(n_23),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1721),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1749),
.A2(n_1730),
.B(n_1708),
.C(n_1715),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1641),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_1656),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1652),
.A2(n_28),
.B1(n_24),
.B2(n_27),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_SL g1815 ( 
.A1(n_1644),
.A2(n_35),
.B1(n_44),
.B2(n_27),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1688),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1643),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1691),
.B(n_28),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1679),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1650),
.B(n_29),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1753),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1701),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1696),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1711),
.A2(n_1709),
.B1(n_1692),
.B2(n_1697),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1655),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1694),
.A2(n_1705),
.B1(n_1706),
.B2(n_1704),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1731),
.B(n_34),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1644),
.A2(n_46),
.B1(n_54),
.B2(n_37),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1657),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1663),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_SL g1831 ( 
.A1(n_1664),
.A2(n_47),
.B1(n_55),
.B2(n_37),
.Y(n_1831)
);

CKINVDCx11_ASAP7_75t_R g1832 ( 
.A(n_1662),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1669),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1660),
.Y(n_1834)
);

OAI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1716),
.A2(n_38),
.B(n_39),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1677),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1693),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1674),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1750),
.A2(n_1766),
.B1(n_1755),
.B2(n_1743),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1681),
.B(n_38),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_SL g1841 ( 
.A1(n_1756),
.A2(n_41),
.B(n_40),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1747),
.A2(n_1748),
.B1(n_1741),
.B2(n_1723),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1724),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1717),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1727),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1718),
.B(n_42),
.Y(n_1846)
);

OAI222xp33_ASAP7_75t_L g1847 ( 
.A1(n_1754),
.A2(n_45),
.B1(n_48),
.B2(n_42),
.C1(n_44),
.C2(n_47),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1729),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1707),
.A2(n_49),
.B(n_48),
.Y(n_1849)
);

OAI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1736),
.A2(n_45),
.B(n_49),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1666),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1733),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1678),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1732),
.A2(n_57),
.B(n_55),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1733),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_SL g1856 ( 
.A1(n_1703),
.A2(n_65),
.B1(n_74),
.B2(n_54),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1726),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1799),
.A2(n_1702),
.B1(n_1682),
.B2(n_1700),
.Y(n_1858)
);

OAI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1841),
.A2(n_1745),
.B1(n_1728),
.B2(n_1746),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1850),
.A2(n_1658),
.B1(n_1713),
.B2(n_1725),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1797),
.B(n_1735),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_L g1862 ( 
.A(n_1811),
.B(n_1751),
.C(n_1739),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1767),
.B(n_1677),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_SL g1864 ( 
.A1(n_1802),
.A2(n_1698),
.B1(n_1765),
.B2(n_1762),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1835),
.A2(n_1719),
.B1(n_1698),
.B2(n_1683),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1773),
.A2(n_1695),
.B1(n_1763),
.B2(n_1683),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_L g1867 ( 
.A(n_1798),
.B(n_60),
.C(n_61),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1821),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1810),
.A2(n_66),
.B1(n_62),
.B2(n_63),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1779),
.A2(n_69),
.B1(n_66),
.B2(n_67),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1775),
.A2(n_71),
.B1(n_67),
.B2(n_70),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1851),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1823),
.A2(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1789),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1793),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1780),
.A2(n_81),
.B1(n_78),
.B2(n_80),
.Y(n_1876)
);

OAI222xp33_ASAP7_75t_L g1877 ( 
.A1(n_1800),
.A2(n_82),
.B1(n_84),
.B2(n_80),
.C1(n_81),
.C2(n_83),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1803),
.A2(n_85),
.B1(n_82),
.B2(n_83),
.Y(n_1878)
);

OAI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1804),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.C(n_89),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1796),
.A2(n_1768),
.B1(n_1783),
.B2(n_1824),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1781),
.A2(n_1857),
.B1(n_1771),
.B2(n_1814),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_SL g1882 ( 
.A1(n_1819),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1812),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_SL g1884 ( 
.A1(n_1769),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1770),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1853),
.A2(n_93),
.B1(n_90),
.B2(n_92),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1839),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1795),
.B(n_94),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1815),
.A2(n_98),
.B1(n_95),
.B2(n_97),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1828),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1856),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1777),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1817),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1825),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_SL g1895 ( 
.A1(n_1843),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1826),
.A2(n_107),
.B1(n_103),
.B2(n_106),
.Y(n_1896)
);

AOI22xp33_ASAP7_75t_L g1897 ( 
.A1(n_1785),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_1897)
);

NAND3xp33_ASAP7_75t_L g1898 ( 
.A(n_1806),
.B(n_110),
.C(n_111),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1831),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1784),
.A2(n_116),
.B1(n_113),
.B2(n_115),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1854),
.A2(n_116),
.B(n_117),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1842),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1902)
);

AOI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1808),
.A2(n_1772),
.B1(n_1847),
.B2(n_1849),
.C(n_1782),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1776),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1786),
.A2(n_1788),
.B1(n_1801),
.B2(n_1778),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1791),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1829),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1774),
.B(n_123),
.Y(n_1908)
);

OAI221xp5_ASAP7_75t_SL g1909 ( 
.A1(n_1846),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.C(n_126),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1805),
.B(n_124),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1791),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1840),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1827),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1822),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1844),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1809),
.A2(n_1818),
.B1(n_1787),
.B2(n_1848),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1820),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_1917)
);

OAI222xp33_ASAP7_75t_L g1918 ( 
.A1(n_1833),
.A2(n_138),
.B1(n_140),
.B2(n_136),
.C1(n_137),
.C2(n_139),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1816),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_L g1920 ( 
.A(n_1794),
.B(n_140),
.C(n_141),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1830),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1838),
.B(n_142),
.Y(n_1922)
);

OAI221xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1834),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1792),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1790),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1845),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1852),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1836),
.B(n_608),
.Y(n_1928)
);

AOI22xp33_ASAP7_75t_L g1929 ( 
.A1(n_1855),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1836),
.B(n_1837),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1807),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_1931)
);

AOI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1832),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1836),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1813),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_SL g1935 ( 
.A1(n_1880),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_L g1936 ( 
.A(n_1867),
.B(n_161),
.C(n_162),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1858),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1907),
.B(n_163),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1885),
.B(n_164),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1920),
.B(n_165),
.C(n_166),
.Y(n_1940)
);

NAND4xp25_ASAP7_75t_L g1941 ( 
.A(n_1909),
.B(n_168),
.C(n_166),
.D(n_167),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1881),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1883),
.B(n_169),
.Y(n_1943)
);

NAND3xp33_ASAP7_75t_L g1944 ( 
.A(n_1898),
.B(n_170),
.C(n_171),
.Y(n_1944)
);

NAND3xp33_ASAP7_75t_L g1945 ( 
.A(n_1923),
.B(n_171),
.C(n_172),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1893),
.B(n_1894),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1863),
.B(n_172),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1861),
.B(n_173),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1916),
.B(n_174),
.Y(n_1949)
);

NAND3xp33_ASAP7_75t_L g1950 ( 
.A(n_1884),
.B(n_174),
.C(n_175),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1922),
.B(n_1927),
.Y(n_1951)
);

OAI21xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1901),
.A2(n_177),
.B(n_176),
.Y(n_1952)
);

OAI221xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1879),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.C(n_178),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1930),
.B(n_179),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1864),
.B(n_180),
.Y(n_1955)
);

OAI21xp5_ASAP7_75t_SL g1956 ( 
.A1(n_1860),
.A2(n_182),
.B(n_181),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1903),
.A2(n_615),
.B(n_611),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1908),
.B(n_180),
.Y(n_1958)
);

OA211x2_ASAP7_75t_L g1959 ( 
.A1(n_1862),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_1959)
);

NOR2xp67_ASAP7_75t_L g1960 ( 
.A(n_1910),
.B(n_183),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1888),
.B(n_184),
.Y(n_1961)
);

OAI221xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1932),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.C(n_188),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1866),
.B(n_185),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1887),
.B(n_188),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1859),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_1965)
);

OA21x2_ASAP7_75t_L g1966 ( 
.A1(n_1918),
.A2(n_190),
.B(n_191),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1865),
.B(n_1905),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1906),
.B(n_1911),
.Y(n_1968)
);

NAND4xp25_ASAP7_75t_L g1969 ( 
.A(n_1931),
.B(n_196),
.C(n_194),
.D(n_195),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1917),
.B(n_1913),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1877),
.A2(n_198),
.B(n_197),
.Y(n_1971)
);

NAND3xp33_ASAP7_75t_L g1972 ( 
.A(n_1892),
.B(n_196),
.C(n_197),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1912),
.B(n_198),
.Y(n_1973)
);

NAND3xp33_ASAP7_75t_L g1974 ( 
.A(n_1872),
.B(n_1871),
.C(n_1875),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1904),
.B(n_1921),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1919),
.B(n_199),
.Y(n_1976)
);

OAI221xp5_ASAP7_75t_L g1977 ( 
.A1(n_1899),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.C(n_202),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1933),
.B(n_200),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1926),
.B(n_201),
.Y(n_1979)
);

OA21x2_ASAP7_75t_L g1980 ( 
.A1(n_1918),
.A2(n_203),
.B(n_204),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1882),
.B(n_203),
.Y(n_1981)
);

NAND3xp33_ASAP7_75t_L g1982 ( 
.A(n_1876),
.B(n_204),
.C(n_205),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_SL g1983 ( 
.A1(n_1928),
.A2(n_617),
.B(n_616),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_SL g1984 ( 
.A1(n_1902),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_1984)
);

INVxp67_ASAP7_75t_SL g1985 ( 
.A(n_1896),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1929),
.B(n_206),
.Y(n_1986)
);

OA21x2_ASAP7_75t_L g1987 ( 
.A1(n_1877),
.A2(n_207),
.B(n_208),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1895),
.B(n_620),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1924),
.B(n_209),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1934),
.B(n_209),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1874),
.B(n_622),
.Y(n_1991)
);

OAI221xp5_ASAP7_75t_SL g1992 ( 
.A1(n_1891),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.C(n_214),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_L g1993 ( 
.A(n_1868),
.B(n_210),
.C(n_211),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1869),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_1994)
);

NAND3xp33_ASAP7_75t_L g1995 ( 
.A(n_1870),
.B(n_215),
.C(n_216),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1925),
.B(n_217),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1889),
.B(n_218),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1914),
.B(n_220),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1890),
.B(n_221),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1915),
.B(n_221),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1873),
.B(n_222),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1886),
.B(n_223),
.Y(n_2002)
);

NAND3xp33_ASAP7_75t_L g2003 ( 
.A(n_1900),
.B(n_224),
.C(n_225),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1897),
.B(n_224),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1878),
.B(n_225),
.Y(n_2005)
);

OAI21xp33_ASAP7_75t_SL g2006 ( 
.A1(n_1887),
.A2(n_226),
.B(n_227),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1907),
.B(n_226),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1907),
.B(n_227),
.Y(n_2008)
);

AOI21xp5_ASAP7_75t_SL g2009 ( 
.A1(n_1880),
.A2(n_624),
.B(n_623),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1858),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1907),
.B(n_228),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1907),
.B(n_229),
.Y(n_2012)
);

OAI21xp5_ASAP7_75t_SL g2013 ( 
.A1(n_1901),
.A2(n_232),
.B(n_231),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1907),
.B(n_230),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1907),
.B(n_231),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1907),
.B(n_232),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1907),
.B(n_233),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1907),
.B(n_234),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1907),
.B(n_234),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1907),
.B(n_235),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1903),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_2021)
);

AOI22xp33_ASAP7_75t_L g2022 ( 
.A1(n_1903),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_2022)
);

NAND3xp33_ASAP7_75t_L g2023 ( 
.A(n_1867),
.B(n_238),
.C(n_239),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1907),
.B(n_239),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1859),
.B(n_625),
.Y(n_2025)
);

OAI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1858),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.C(n_243),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1946),
.B(n_241),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1951),
.B(n_242),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1948),
.B(n_244),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1943),
.Y(n_2030)
);

NAND4xp75_ASAP7_75t_L g2031 ( 
.A(n_1959),
.B(n_246),
.C(n_244),
.D(n_245),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_2011),
.B(n_245),
.Y(n_2032)
);

AO21x2_ASAP7_75t_L g2033 ( 
.A1(n_1957),
.A2(n_247),
.B(n_248),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_2012),
.B(n_248),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1961),
.B(n_249),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1958),
.B(n_249),
.Y(n_2036)
);

HB1xp67_ASAP7_75t_L g2037 ( 
.A(n_2015),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1939),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1954),
.B(n_250),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1938),
.B(n_250),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1974),
.A2(n_254),
.B1(n_251),
.B2(n_252),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2007),
.B(n_251),
.Y(n_2042)
);

NAND3xp33_ASAP7_75t_L g2043 ( 
.A(n_1940),
.B(n_252),
.C(n_254),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_2008),
.B(n_256),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_1941),
.A2(n_259),
.B1(n_256),
.B2(n_258),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2014),
.B(n_259),
.Y(n_2046)
);

NAND4xp75_ASAP7_75t_L g2047 ( 
.A(n_1987),
.B(n_1966),
.C(n_1980),
.D(n_2025),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2016),
.B(n_260),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1945),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2020),
.B(n_261),
.Y(n_2050)
);

NAND3xp33_ASAP7_75t_SL g2051 ( 
.A(n_1971),
.B(n_262),
.C(n_263),
.Y(n_2051)
);

AO21x2_ASAP7_75t_L g2052 ( 
.A1(n_1949),
.A2(n_264),
.B(n_265),
.Y(n_2052)
);

NOR3xp33_ASAP7_75t_L g2053 ( 
.A(n_1953),
.B(n_264),
.C(n_265),
.Y(n_2053)
);

NOR2x1_ASAP7_75t_L g2054 ( 
.A(n_2017),
.B(n_266),
.Y(n_2054)
);

NAND4xp75_ASAP7_75t_L g2055 ( 
.A(n_1987),
.B(n_268),
.C(n_266),
.D(n_267),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_1952),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_L g2057 ( 
.A(n_1935),
.B(n_270),
.C(n_271),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_1936),
.B(n_271),
.C(n_272),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2018),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2019),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_2024),
.Y(n_2061)
);

NAND2x1p5_ASAP7_75t_L g2062 ( 
.A(n_1966),
.B(n_626),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1937),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_2063)
);

OAI211xp5_ASAP7_75t_SL g2064 ( 
.A1(n_1990),
.A2(n_276),
.B(n_273),
.C(n_274),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_2026),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1947),
.B(n_277),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1963),
.Y(n_2067)
);

OAI211xp5_ASAP7_75t_L g2068 ( 
.A1(n_2013),
.A2(n_288),
.B(n_296),
.C(n_278),
.Y(n_2068)
);

OAI21xp33_ASAP7_75t_L g2069 ( 
.A1(n_1969),
.A2(n_280),
.B(n_281),
.Y(n_2069)
);

NOR2x1_ASAP7_75t_L g2070 ( 
.A(n_2009),
.B(n_280),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_1972),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_2071)
);

AO21x2_ASAP7_75t_L g2072 ( 
.A1(n_1944),
.A2(n_2023),
.B(n_1982),
.Y(n_2072)
);

NAND3xp33_ASAP7_75t_L g2073 ( 
.A(n_1950),
.B(n_282),
.C(n_283),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1967),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1960),
.B(n_284),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1955),
.B(n_284),
.Y(n_2076)
);

AOI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_1993),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.Y(n_2077)
);

NOR3xp33_ASAP7_75t_L g2078 ( 
.A(n_1962),
.B(n_287),
.C(n_289),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_1985),
.B(n_289),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_1970),
.B(n_290),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_1975),
.B(n_290),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_1956),
.B(n_291),
.Y(n_2082)
);

AOI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_1992),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.C(n_294),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1981),
.B(n_295),
.Y(n_2084)
);

AO21x2_ASAP7_75t_L g2085 ( 
.A1(n_1976),
.A2(n_295),
.B(n_296),
.Y(n_2085)
);

INVx3_ASAP7_75t_L g2086 ( 
.A(n_1980),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1998),
.B(n_297),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2000),
.B(n_297),
.Y(n_2088)
);

AO21x2_ASAP7_75t_L g2089 ( 
.A1(n_1973),
.A2(n_1999),
.B(n_1997),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1968),
.B(n_1978),
.Y(n_2090)
);

NOR2x1_ASAP7_75t_L g2091 ( 
.A(n_1983),
.B(n_298),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1979),
.B(n_1942),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1964),
.Y(n_2093)
);

NAND3xp33_ASAP7_75t_L g2094 ( 
.A(n_2021),
.B(n_299),
.C(n_300),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1986),
.B(n_299),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1988),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_2010),
.B(n_301),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_1996),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1989),
.B(n_303),
.Y(n_2099)
);

INVxp67_ASAP7_75t_L g2100 ( 
.A(n_2004),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1965),
.B(n_304),
.Y(n_2101)
);

NOR2x1_ASAP7_75t_L g2102 ( 
.A(n_2003),
.B(n_304),
.Y(n_2102)
);

NOR3xp33_ASAP7_75t_L g2103 ( 
.A(n_1977),
.B(n_306),
.C(n_308),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2002),
.B(n_306),
.Y(n_2104)
);

NAND4xp75_ASAP7_75t_L g2105 ( 
.A(n_2006),
.B(n_310),
.C(n_308),
.D(n_309),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_2001),
.Y(n_2106)
);

AOI22xp33_ASAP7_75t_L g2107 ( 
.A1(n_2022),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_2005),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1995),
.Y(n_2109)
);

OAI211xp5_ASAP7_75t_SL g2110 ( 
.A1(n_1984),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1991),
.B(n_312),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1994),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1946),
.B(n_313),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1946),
.B(n_314),
.Y(n_2114)
);

NAND3xp33_ASAP7_75t_SL g2115 ( 
.A(n_1971),
.B(n_315),
.C(n_316),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1954),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1946),
.Y(n_2117)
);

NOR3xp33_ASAP7_75t_L g2118 ( 
.A(n_1953),
.B(n_315),
.C(n_317),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1946),
.Y(n_2119)
);

INVx2_ASAP7_75t_SL g2120 ( 
.A(n_1938),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1951),
.B(n_317),
.Y(n_2121)
);

AO21x2_ASAP7_75t_L g2122 ( 
.A1(n_1957),
.A2(n_318),
.B(n_319),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1946),
.B(n_318),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1946),
.B(n_319),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2117),
.Y(n_2125)
);

HB1xp67_ASAP7_75t_L g2126 ( 
.A(n_2119),
.Y(n_2126)
);

XNOR2xp5_ASAP7_75t_L g2127 ( 
.A(n_2116),
.B(n_320),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_2037),
.B(n_320),
.Y(n_2128)
);

NAND3xp33_ASAP7_75t_SL g2129 ( 
.A(n_2053),
.B(n_324),
.C(n_323),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2074),
.B(n_321),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2086),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2086),
.Y(n_2132)
);

INVx1_ASAP7_75t_SL g2133 ( 
.A(n_2059),
.Y(n_2133)
);

NOR3xp33_ASAP7_75t_SL g2134 ( 
.A(n_2051),
.B(n_323),
.C(n_324),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2061),
.B(n_325),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_2060),
.Y(n_2136)
);

NAND4xp75_ASAP7_75t_SL g2137 ( 
.A(n_2082),
.B(n_2097),
.C(n_2111),
.D(n_2101),
.Y(n_2137)
);

INVxp33_ASAP7_75t_SL g2138 ( 
.A(n_2029),
.Y(n_2138)
);

XOR2xp5_ASAP7_75t_L g2139 ( 
.A(n_2080),
.B(n_628),
.Y(n_2139)
);

OAI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_2056),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2038),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2067),
.B(n_327),
.Y(n_2142)
);

BUFx4f_ASAP7_75t_L g2143 ( 
.A(n_2066),
.Y(n_2143)
);

BUFx2_ASAP7_75t_L g2144 ( 
.A(n_2038),
.Y(n_2144)
);

INVxp67_ASAP7_75t_SL g2145 ( 
.A(n_2030),
.Y(n_2145)
);

NAND3xp33_ASAP7_75t_SL g2146 ( 
.A(n_2118),
.B(n_2078),
.C(n_2103),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2100),
.B(n_328),
.Y(n_2147)
);

NAND4xp75_ASAP7_75t_SL g2148 ( 
.A(n_2036),
.B(n_333),
.C(n_329),
.D(n_332),
.Y(n_2148)
);

INVx2_ASAP7_75t_SL g2149 ( 
.A(n_2028),
.Y(n_2149)
);

XNOR2xp5_ASAP7_75t_L g2150 ( 
.A(n_2098),
.B(n_333),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2108),
.B(n_334),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2030),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2093),
.Y(n_2153)
);

NOR2x1_ASAP7_75t_R g2154 ( 
.A(n_2095),
.B(n_336),
.Y(n_2154)
);

INVxp67_ASAP7_75t_L g2155 ( 
.A(n_2054),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2106),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2093),
.Y(n_2157)
);

NAND2xp33_ASAP7_75t_R g2158 ( 
.A(n_2081),
.B(n_2075),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2089),
.B(n_336),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2027),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2113),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_2039),
.Y(n_2162)
);

XOR2x2_ASAP7_75t_L g2163 ( 
.A(n_2115),
.B(n_337),
.Y(n_2163)
);

NAND4xp75_ASAP7_75t_SL g2164 ( 
.A(n_2104),
.B(n_2035),
.C(n_2099),
.D(n_2070),
.Y(n_2164)
);

BUFx2_ASAP7_75t_SL g2165 ( 
.A(n_2114),
.Y(n_2165)
);

NAND4xp75_ASAP7_75t_L g2166 ( 
.A(n_2091),
.B(n_339),
.C(n_337),
.D(n_338),
.Y(n_2166)
);

NAND4xp75_ASAP7_75t_SL g2167 ( 
.A(n_2088),
.B(n_340),
.C(n_338),
.D(n_339),
.Y(n_2167)
);

XOR2x2_ASAP7_75t_L g2168 ( 
.A(n_2076),
.B(n_340),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2123),
.Y(n_2169)
);

XOR2x2_ASAP7_75t_L g2170 ( 
.A(n_2084),
.B(n_341),
.Y(n_2170)
);

INVxp67_ASAP7_75t_L g2171 ( 
.A(n_2048),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2124),
.B(n_341),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2121),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2109),
.B(n_342),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2032),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2079),
.Y(n_2176)
);

INVx2_ASAP7_75t_SL g2177 ( 
.A(n_2034),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2052),
.Y(n_2178)
);

INVxp67_ASAP7_75t_L g2179 ( 
.A(n_2040),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2087),
.B(n_342),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2085),
.B(n_343),
.Y(n_2181)
);

INVxp67_ASAP7_75t_SL g2182 ( 
.A(n_2062),
.Y(n_2182)
);

BUFx2_ASAP7_75t_L g2183 ( 
.A(n_2095),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2047),
.Y(n_2184)
);

XOR2x2_ASAP7_75t_L g2185 ( 
.A(n_2042),
.B(n_2044),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2046),
.B(n_343),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2092),
.B(n_344),
.Y(n_2187)
);

INVx5_ASAP7_75t_L g2188 ( 
.A(n_2050),
.Y(n_2188)
);

HB1xp67_ASAP7_75t_L g2189 ( 
.A(n_2072),
.Y(n_2189)
);

BUFx2_ASAP7_75t_L g2190 ( 
.A(n_2033),
.Y(n_2190)
);

OAI31xp33_ASAP7_75t_L g2191 ( 
.A1(n_2068),
.A2(n_346),
.A3(n_344),
.B(n_345),
.Y(n_2191)
);

NAND4xp75_ASAP7_75t_SL g2192 ( 
.A(n_2055),
.B(n_348),
.C(n_346),
.D(n_347),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2122),
.Y(n_2193)
);

OAI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_2063),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_2194)
);

NAND4xp75_ASAP7_75t_L g2195 ( 
.A(n_2102),
.B(n_351),
.C(n_349),
.D(n_350),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2058),
.Y(n_2196)
);

INVx3_ASAP7_75t_L g2197 ( 
.A(n_2112),
.Y(n_2197)
);

INVx6_ASAP7_75t_L g2198 ( 
.A(n_2031),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2043),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2069),
.B(n_351),
.Y(n_2200)
);

BUFx2_ASAP7_75t_L g2201 ( 
.A(n_2073),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2041),
.B(n_352),
.Y(n_2202)
);

OAI31xp33_ASAP7_75t_L g2203 ( 
.A1(n_2064),
.A2(n_354),
.A3(n_352),
.B(n_353),
.Y(n_2203)
);

NOR2xp33_ASAP7_75t_L g2204 ( 
.A(n_2057),
.B(n_353),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_2105),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_2083),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2071),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2049),
.B(n_354),
.Y(n_2208)
);

NAND3xp33_ASAP7_75t_L g2209 ( 
.A(n_2077),
.B(n_355),
.C(n_356),
.Y(n_2209)
);

INVx1_ASAP7_75t_SL g2210 ( 
.A(n_2094),
.Y(n_2210)
);

NOR4xp25_ASAP7_75t_L g2211 ( 
.A(n_2110),
.B(n_357),
.C(n_355),
.D(n_356),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2045),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_2096),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2065),
.B(n_358),
.Y(n_2214)
);

NAND4xp75_ASAP7_75t_L g2215 ( 
.A(n_2107),
.B(n_360),
.C(n_358),
.D(n_359),
.Y(n_2215)
);

XNOR2xp5_ASAP7_75t_L g2216 ( 
.A(n_2116),
.B(n_360),
.Y(n_2216)
);

XOR2x2_ASAP7_75t_L g2217 ( 
.A(n_2090),
.B(n_361),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_L g2218 ( 
.A(n_2074),
.B(n_361),
.Y(n_2218)
);

HB1xp67_ASAP7_75t_L g2219 ( 
.A(n_2117),
.Y(n_2219)
);

XNOR2xp5_ASAP7_75t_L g2220 ( 
.A(n_2116),
.B(n_362),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2117),
.Y(n_2221)
);

AOI211xp5_ASAP7_75t_SL g2222 ( 
.A1(n_2068),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2117),
.Y(n_2223)
);

INVx2_ASAP7_75t_SL g2224 ( 
.A(n_2120),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2037),
.B(n_363),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2119),
.B(n_364),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2117),
.Y(n_2227)
);

INVx4_ASAP7_75t_L g2228 ( 
.A(n_2052),
.Y(n_2228)
);

INVx2_ASAP7_75t_SL g2229 ( 
.A(n_2120),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_R g2230 ( 
.A(n_2116),
.B(n_365),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2037),
.B(n_366),
.Y(n_2231)
);

AOI22x1_ASAP7_75t_SL g2232 ( 
.A1(n_2184),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_2232)
);

XNOR2x1_ASAP7_75t_L g2233 ( 
.A(n_2217),
.B(n_368),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2131),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2145),
.Y(n_2235)
);

XNOR2xp5_ASAP7_75t_L g2236 ( 
.A(n_2168),
.B(n_367),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2126),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2197),
.B(n_369),
.Y(n_2238)
);

INVx5_ASAP7_75t_L g2239 ( 
.A(n_2228),
.Y(n_2239)
);

XOR2x2_ASAP7_75t_L g2240 ( 
.A(n_2170),
.B(n_370),
.Y(n_2240)
);

INVx4_ASAP7_75t_L g2241 ( 
.A(n_2188),
.Y(n_2241)
);

INVx2_ASAP7_75t_SL g2242 ( 
.A(n_2188),
.Y(n_2242)
);

INVx4_ASAP7_75t_L g2243 ( 
.A(n_2188),
.Y(n_2243)
);

AOI22x1_ASAP7_75t_SL g2244 ( 
.A1(n_2210),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2153),
.Y(n_2245)
);

INVxp67_ASAP7_75t_L g2246 ( 
.A(n_2189),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_L g2247 ( 
.A(n_2173),
.B(n_372),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2157),
.Y(n_2248)
);

XOR2x2_ASAP7_75t_L g2249 ( 
.A(n_2185),
.B(n_373),
.Y(n_2249)
);

OA22x2_ASAP7_75t_L g2250 ( 
.A1(n_2155),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_SL g2251 ( 
.A1(n_2201),
.A2(n_376),
.B1(n_377),
.B2(n_375),
.Y(n_2251)
);

XOR2xp5_ASAP7_75t_L g2252 ( 
.A(n_2127),
.B(n_374),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2132),
.Y(n_2253)
);

XOR2x2_ASAP7_75t_L g2254 ( 
.A(n_2216),
.B(n_378),
.Y(n_2254)
);

XOR2x2_ASAP7_75t_L g2255 ( 
.A(n_2220),
.B(n_2164),
.Y(n_2255)
);

XOR2x2_ASAP7_75t_L g2256 ( 
.A(n_2137),
.B(n_379),
.Y(n_2256)
);

XOR2x2_ASAP7_75t_L g2257 ( 
.A(n_2150),
.B(n_379),
.Y(n_2257)
);

INVxp33_ASAP7_75t_SL g2258 ( 
.A(n_2230),
.Y(n_2258)
);

INVx2_ASAP7_75t_SL g2259 ( 
.A(n_2183),
.Y(n_2259)
);

XOR2x2_ASAP7_75t_L g2260 ( 
.A(n_2138),
.B(n_380),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2175),
.B(n_381),
.Y(n_2261)
);

XOR2xp5_ASAP7_75t_L g2262 ( 
.A(n_2139),
.B(n_382),
.Y(n_2262)
);

XOR2x2_ASAP7_75t_L g2263 ( 
.A(n_2163),
.B(n_2146),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2141),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2152),
.Y(n_2265)
);

XOR2x2_ASAP7_75t_L g2266 ( 
.A(n_2206),
.B(n_383),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2144),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2133),
.B(n_383),
.Y(n_2268)
);

XNOR2xp5_ASAP7_75t_L g2269 ( 
.A(n_2213),
.B(n_384),
.Y(n_2269)
);

INVxp67_ASAP7_75t_SL g2270 ( 
.A(n_2159),
.Y(n_2270)
);

AO22x1_ASAP7_75t_L g2271 ( 
.A1(n_2228),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_2271)
);

XOR2x2_ASAP7_75t_L g2272 ( 
.A(n_2192),
.B(n_385),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2156),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2136),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2125),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2219),
.Y(n_2276)
);

XNOR2x1_ASAP7_75t_L g2277 ( 
.A(n_2162),
.B(n_388),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2223),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2221),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2178),
.B(n_387),
.Y(n_2280)
);

XOR2x2_ASAP7_75t_L g2281 ( 
.A(n_2148),
.B(n_389),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2227),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2171),
.B(n_2174),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2224),
.B(n_390),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2149),
.B(n_390),
.Y(n_2285)
);

XNOR2x1_ASAP7_75t_L g2286 ( 
.A(n_2186),
.B(n_392),
.Y(n_2286)
);

INVx1_ASAP7_75t_SL g2287 ( 
.A(n_2165),
.Y(n_2287)
);

XNOR2xp5_ASAP7_75t_L g2288 ( 
.A(n_2167),
.B(n_391),
.Y(n_2288)
);

XOR2x2_ASAP7_75t_L g2289 ( 
.A(n_2187),
.B(n_392),
.Y(n_2289)
);

XNOR2xp5_ASAP7_75t_L g2290 ( 
.A(n_2172),
.B(n_393),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2229),
.B(n_393),
.Y(n_2291)
);

INVx1_ASAP7_75t_SL g2292 ( 
.A(n_2128),
.Y(n_2292)
);

INVx1_ASAP7_75t_SL g2293 ( 
.A(n_2151),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_2177),
.B(n_394),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2176),
.Y(n_2295)
);

XNOR2x1_ASAP7_75t_L g2296 ( 
.A(n_2180),
.B(n_2161),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_2158),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2193),
.Y(n_2298)
);

XOR2x2_ASAP7_75t_L g2299 ( 
.A(n_2166),
.B(n_394),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_2169),
.Y(n_2300)
);

INVxp67_ASAP7_75t_L g2301 ( 
.A(n_2154),
.Y(n_2301)
);

XOR2x2_ASAP7_75t_L g2302 ( 
.A(n_2195),
.B(n_396),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2190),
.Y(n_2303)
);

XOR2x2_ASAP7_75t_L g2304 ( 
.A(n_2129),
.B(n_396),
.Y(n_2304)
);

INVxp67_ASAP7_75t_L g2305 ( 
.A(n_2181),
.Y(n_2305)
);

NOR2x1_ASAP7_75t_R g2306 ( 
.A(n_2198),
.B(n_397),
.Y(n_2306)
);

XOR2x2_ASAP7_75t_L g2307 ( 
.A(n_2222),
.B(n_397),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2160),
.Y(n_2308)
);

HB1xp67_ASAP7_75t_L g2309 ( 
.A(n_2179),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2182),
.B(n_398),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2226),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_2143),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2135),
.Y(n_2313)
);

AND2x4_ASAP7_75t_L g2314 ( 
.A(n_2225),
.B(n_398),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2147),
.Y(n_2315)
);

XNOR2xp5_ASAP7_75t_L g2316 ( 
.A(n_2205),
.B(n_399),
.Y(n_2316)
);

XNOR2x1_ASAP7_75t_L g2317 ( 
.A(n_2231),
.B(n_400),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2196),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2142),
.Y(n_2319)
);

XNOR2x1_ASAP7_75t_L g2320 ( 
.A(n_2130),
.B(n_400),
.Y(n_2320)
);

INVx1_ASAP7_75t_SL g2321 ( 
.A(n_2198),
.Y(n_2321)
);

INVxp33_ASAP7_75t_L g2322 ( 
.A(n_2218),
.Y(n_2322)
);

XNOR2xp5_ASAP7_75t_L g2323 ( 
.A(n_2212),
.B(n_399),
.Y(n_2323)
);

XNOR2xp5_ASAP7_75t_L g2324 ( 
.A(n_2207),
.B(n_401),
.Y(n_2324)
);

CKINVDCx16_ASAP7_75t_R g2325 ( 
.A(n_2204),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2199),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2200),
.Y(n_2327)
);

XNOR2x2_ASAP7_75t_L g2328 ( 
.A(n_2215),
.B(n_402),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2208),
.Y(n_2329)
);

XOR2xp5_ASAP7_75t_L g2330 ( 
.A(n_2209),
.B(n_402),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2202),
.Y(n_2331)
);

XOR2x2_ASAP7_75t_L g2332 ( 
.A(n_2214),
.B(n_403),
.Y(n_2332)
);

XOR2x2_ASAP7_75t_L g2333 ( 
.A(n_2194),
.B(n_403),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2203),
.Y(n_2334)
);

XOR2x2_ASAP7_75t_L g2335 ( 
.A(n_2191),
.B(n_404),
.Y(n_2335)
);

INVx1_ASAP7_75t_SL g2336 ( 
.A(n_2134),
.Y(n_2336)
);

XNOR2xp5_ASAP7_75t_L g2337 ( 
.A(n_2140),
.B(n_405),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2211),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2131),
.Y(n_2339)
);

NOR2x1_ASAP7_75t_L g2340 ( 
.A(n_2228),
.B(n_405),
.Y(n_2340)
);

INVxp67_ASAP7_75t_SL g2341 ( 
.A(n_2189),
.Y(n_2341)
);

INVx1_ASAP7_75t_SL g2342 ( 
.A(n_2230),
.Y(n_2342)
);

OA22x2_ASAP7_75t_L g2343 ( 
.A1(n_2155),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2189),
.B(n_408),
.Y(n_2344)
);

XOR2x2_ASAP7_75t_L g2345 ( 
.A(n_2217),
.B(n_409),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2264),
.Y(n_2346)
);

INVx1_ASAP7_75t_SL g2347 ( 
.A(n_2342),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2241),
.Y(n_2348)
);

OA22x2_ASAP7_75t_L g2349 ( 
.A1(n_2297),
.A2(n_2338),
.B1(n_2334),
.B2(n_2321),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2273),
.Y(n_2350)
);

OA22x2_ASAP7_75t_L g2351 ( 
.A1(n_2287),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_2351)
);

OA22x2_ASAP7_75t_L g2352 ( 
.A1(n_2316),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_2352)
);

AO22x2_ASAP7_75t_L g2353 ( 
.A1(n_2243),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2295),
.Y(n_2354)
);

AOI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_2263),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_2355)
);

OA22x2_ASAP7_75t_L g2356 ( 
.A1(n_2330),
.A2(n_418),
.B1(n_415),
.B2(n_416),
.Y(n_2356)
);

INVxp67_ASAP7_75t_L g2357 ( 
.A(n_2306),
.Y(n_2357)
);

OA22x2_ASAP7_75t_L g2358 ( 
.A1(n_2324),
.A2(n_420),
.B1(n_416),
.B2(n_418),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2325),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_2359)
);

INVxp67_ASAP7_75t_SL g2360 ( 
.A(n_2340),
.Y(n_2360)
);

AO22x1_ASAP7_75t_L g2361 ( 
.A1(n_2239),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2279),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_SL g2363 ( 
.A1(n_2258),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_2363)
);

OA22x2_ASAP7_75t_L g2364 ( 
.A1(n_2336),
.A2(n_427),
.B1(n_424),
.B2(n_426),
.Y(n_2364)
);

INVx3_ASAP7_75t_L g2365 ( 
.A(n_2312),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2282),
.Y(n_2366)
);

AOI22x1_ASAP7_75t_L g2367 ( 
.A1(n_2251),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_2367)
);

INVx2_ASAP7_75t_SL g2368 ( 
.A(n_2242),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2309),
.Y(n_2369)
);

INVxp33_ASAP7_75t_L g2370 ( 
.A(n_2283),
.Y(n_2370)
);

AO22x1_ASAP7_75t_L g2371 ( 
.A1(n_2239),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_2371)
);

AOI22x1_ASAP7_75t_L g2372 ( 
.A1(n_2236),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_2372)
);

AOI22x1_ASAP7_75t_L g2373 ( 
.A1(n_2337),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_2373)
);

OA22x2_ASAP7_75t_L g2374 ( 
.A1(n_2323),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_2374)
);

AOI22x1_ASAP7_75t_L g2375 ( 
.A1(n_2269),
.A2(n_438),
.B1(n_435),
.B2(n_437),
.Y(n_2375)
);

OAI22xp5_ASAP7_75t_SL g2376 ( 
.A1(n_2301),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2318),
.Y(n_2377)
);

XNOR2x1_ASAP7_75t_L g2378 ( 
.A(n_2249),
.B(n_440),
.Y(n_2378)
);

XOR2x2_ASAP7_75t_L g2379 ( 
.A(n_2255),
.B(n_440),
.Y(n_2379)
);

OA22x2_ASAP7_75t_L g2380 ( 
.A1(n_2326),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_2235),
.Y(n_2381)
);

XNOR2xp5_ASAP7_75t_L g2382 ( 
.A(n_2345),
.B(n_442),
.Y(n_2382)
);

AO22x1_ASAP7_75t_L g2383 ( 
.A1(n_2239),
.A2(n_2270),
.B1(n_2322),
.B2(n_2344),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2237),
.Y(n_2384)
);

OA22x2_ASAP7_75t_L g2385 ( 
.A1(n_2259),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_2385)
);

INVx2_ASAP7_75t_SL g2386 ( 
.A(n_2274),
.Y(n_2386)
);

INVx2_ASAP7_75t_SL g2387 ( 
.A(n_2319),
.Y(n_2387)
);

INVx2_ASAP7_75t_SL g2388 ( 
.A(n_2300),
.Y(n_2388)
);

AO22x1_ASAP7_75t_L g2389 ( 
.A1(n_2247),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_2389)
);

AOI22x1_ASAP7_75t_L g2390 ( 
.A1(n_2252),
.A2(n_450),
.B1(n_447),
.B2(n_448),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2308),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2245),
.Y(n_2392)
);

AOI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_2335),
.A2(n_451),
.B1(n_447),
.B2(n_450),
.Y(n_2393)
);

AO22x1_ASAP7_75t_L g2394 ( 
.A1(n_2310),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_2394)
);

INVxp67_ASAP7_75t_SL g2395 ( 
.A(n_2296),
.Y(n_2395)
);

OA22x2_ASAP7_75t_L g2396 ( 
.A1(n_2305),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2248),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_2314),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2298),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_2315),
.B(n_454),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2234),
.Y(n_2401)
);

AO22x2_ASAP7_75t_L g2402 ( 
.A1(n_2303),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_2402)
);

BUFx3_ASAP7_75t_L g2403 ( 
.A(n_2284),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2265),
.Y(n_2404)
);

AOI22x1_ASAP7_75t_L g2405 ( 
.A1(n_2288),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2275),
.Y(n_2406)
);

OAI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2233),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_2407)
);

OA22x2_ASAP7_75t_L g2408 ( 
.A1(n_2293),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_2408)
);

AO22x2_ASAP7_75t_L g2409 ( 
.A1(n_2232),
.A2(n_464),
.B1(n_462),
.B2(n_463),
.Y(n_2409)
);

OAI22x1_ASAP7_75t_L g2410 ( 
.A1(n_2292),
.A2(n_466),
.B1(n_462),
.B2(n_463),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2253),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2256),
.A2(n_469),
.B1(n_467),
.B2(n_468),
.Y(n_2412)
);

XNOR2xp5_ASAP7_75t_L g2413 ( 
.A(n_2240),
.B(n_468),
.Y(n_2413)
);

OA22x2_ASAP7_75t_L g2414 ( 
.A1(n_2290),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_2414)
);

XOR2x2_ASAP7_75t_L g2415 ( 
.A(n_2266),
.B(n_470),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2276),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2267),
.Y(n_2417)
);

AO22x1_ASAP7_75t_L g2418 ( 
.A1(n_2341),
.A2(n_474),
.B1(n_471),
.B2(n_472),
.Y(n_2418)
);

AO22x1_ASAP7_75t_L g2419 ( 
.A1(n_2238),
.A2(n_475),
.B1(n_472),
.B2(n_474),
.Y(n_2419)
);

BUFx2_ASAP7_75t_L g2420 ( 
.A(n_2327),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2339),
.Y(n_2421)
);

XNOR2xp5_ASAP7_75t_L g2422 ( 
.A(n_2254),
.B(n_475),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_2246),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2278),
.Y(n_2424)
);

AOI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2307),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2280),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2250),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_2427)
);

OA22x2_ASAP7_75t_L g2428 ( 
.A1(n_2329),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_2428)
);

OA22x2_ASAP7_75t_L g2429 ( 
.A1(n_2331),
.A2(n_482),
.B1(n_479),
.B2(n_480),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_2311),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2313),
.Y(n_2431)
);

OR2x2_ASAP7_75t_L g2432 ( 
.A(n_2268),
.B(n_2285),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2291),
.Y(n_2433)
);

AOI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2304),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2261),
.Y(n_2435)
);

AOI22x1_ASAP7_75t_L g2436 ( 
.A1(n_2262),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_2294),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_2277),
.Y(n_2438)
);

INVxp67_ASAP7_75t_L g2439 ( 
.A(n_2244),
.Y(n_2439)
);

XNOR2x2_ASAP7_75t_L g2440 ( 
.A(n_2328),
.B(n_487),
.Y(n_2440)
);

OA22x2_ASAP7_75t_L g2441 ( 
.A1(n_2343),
.A2(n_490),
.B1(n_487),
.B2(n_489),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2271),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2289),
.Y(n_2443)
);

OA22x2_ASAP7_75t_L g2444 ( 
.A1(n_2260),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_2444)
);

CKINVDCx14_ASAP7_75t_R g2445 ( 
.A(n_2332),
.Y(n_2445)
);

BUFx3_ASAP7_75t_L g2446 ( 
.A(n_2320),
.Y(n_2446)
);

AOI22xp5_ASAP7_75t_L g2447 ( 
.A1(n_2333),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_2447)
);

XOR2x2_ASAP7_75t_L g2448 ( 
.A(n_2257),
.B(n_493),
.Y(n_2448)
);

INVx2_ASAP7_75t_SL g2449 ( 
.A(n_2317),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2302),
.Y(n_2450)
);

OA22x2_ASAP7_75t_L g2451 ( 
.A1(n_2299),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2286),
.Y(n_2452)
);

OA22x2_ASAP7_75t_L g2453 ( 
.A1(n_2281),
.A2(n_498),
.B1(n_494),
.B2(n_497),
.Y(n_2453)
);

OA22x2_ASAP7_75t_L g2454 ( 
.A1(n_2272),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_2454)
);

INVx1_ASAP7_75t_SL g2455 ( 
.A(n_2342),
.Y(n_2455)
);

INVx2_ASAP7_75t_SL g2456 ( 
.A(n_2241),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2242),
.Y(n_2457)
);

AO22x2_ASAP7_75t_L g2458 ( 
.A1(n_2241),
.A2(n_503),
.B1(n_501),
.B2(n_502),
.Y(n_2458)
);

OA22x2_ASAP7_75t_L g2459 ( 
.A1(n_2297),
.A2(n_503),
.B1(n_501),
.B2(n_502),
.Y(n_2459)
);

OAI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2297),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_2460)
);

XNOR2x1_ASAP7_75t_L g2461 ( 
.A(n_2249),
.B(n_505),
.Y(n_2461)
);

AOI22x1_ASAP7_75t_L g2462 ( 
.A1(n_2297),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2264),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2264),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2242),
.Y(n_2465)
);

OA22x2_ASAP7_75t_L g2466 ( 
.A1(n_2297),
.A2(n_510),
.B1(n_508),
.B2(n_509),
.Y(n_2466)
);

AO22x2_ASAP7_75t_L g2467 ( 
.A1(n_2241),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.Y(n_2467)
);

OA22x2_ASAP7_75t_L g2468 ( 
.A1(n_2297),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_2468)
);

INVx2_ASAP7_75t_SL g2469 ( 
.A(n_2241),
.Y(n_2469)
);

OA22x2_ASAP7_75t_L g2470 ( 
.A1(n_2297),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.Y(n_2470)
);

AOI22xp5_ASAP7_75t_L g2471 ( 
.A1(n_2334),
.A2(n_516),
.B1(n_514),
.B2(n_515),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2270),
.B(n_515),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2264),
.Y(n_2473)
);

HB1xp67_ASAP7_75t_L g2474 ( 
.A(n_2235),
.Y(n_2474)
);

OA22x2_ASAP7_75t_L g2475 ( 
.A1(n_2297),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2264),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2242),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2264),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2264),
.Y(n_2479)
);

INVx2_ASAP7_75t_SL g2480 ( 
.A(n_2241),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_SL g2481 ( 
.A1(n_2297),
.A2(n_520),
.B1(n_517),
.B2(n_519),
.Y(n_2481)
);

OAI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2297),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.Y(n_2482)
);

OA22x2_ASAP7_75t_L g2483 ( 
.A1(n_2297),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2264),
.Y(n_2484)
);

OA22x2_ASAP7_75t_L g2485 ( 
.A1(n_2297),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_2485)
);

AO22x1_ASAP7_75t_L g2486 ( 
.A1(n_2297),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2242),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2264),
.Y(n_2488)
);

OA22x2_ASAP7_75t_L g2489 ( 
.A1(n_2297),
.A2(n_529),
.B1(n_527),
.B2(n_528),
.Y(n_2489)
);

XOR2x2_ASAP7_75t_L g2490 ( 
.A(n_2255),
.B(n_527),
.Y(n_2490)
);

AOI22x1_ASAP7_75t_L g2491 ( 
.A1(n_2297),
.A2(n_530),
.B1(n_528),
.B2(n_529),
.Y(n_2491)
);

XOR2xp5_ASAP7_75t_L g2492 ( 
.A(n_2236),
.B(n_531),
.Y(n_2492)
);

XOR2x2_ASAP7_75t_L g2493 ( 
.A(n_2255),
.B(n_531),
.Y(n_2493)
);

AO22x2_ASAP7_75t_L g2494 ( 
.A1(n_2241),
.A2(n_535),
.B1(n_532),
.B2(n_534),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2242),
.Y(n_2495)
);

OA22x2_ASAP7_75t_L g2496 ( 
.A1(n_2297),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_2496)
);

OA22x2_ASAP7_75t_L g2497 ( 
.A1(n_2297),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_2497)
);

OA22x2_ASAP7_75t_L g2498 ( 
.A1(n_2297),
.A2(n_542),
.B1(n_539),
.B2(n_540),
.Y(n_2498)
);

OA22x2_ASAP7_75t_L g2499 ( 
.A1(n_2297),
.A2(n_542),
.B1(n_539),
.B2(n_540),
.Y(n_2499)
);

AOI22x1_ASAP7_75t_L g2500 ( 
.A1(n_2297),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_2500)
);

OAI22x1_ASAP7_75t_SL g2501 ( 
.A1(n_2258),
.A2(n_546),
.B1(n_543),
.B2(n_545),
.Y(n_2501)
);

OAI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2297),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.Y(n_2502)
);

OA22x2_ASAP7_75t_L g2503 ( 
.A1(n_2297),
.A2(n_550),
.B1(n_547),
.B2(n_549),
.Y(n_2503)
);

OA22x2_ASAP7_75t_L g2504 ( 
.A1(n_2297),
.A2(n_552),
.B1(n_550),
.B2(n_551),
.Y(n_2504)
);

HB1xp67_ASAP7_75t_L g2505 ( 
.A(n_2235),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2264),
.Y(n_2506)
);

HB1xp67_ASAP7_75t_L g2507 ( 
.A(n_2235),
.Y(n_2507)
);

OA22x2_ASAP7_75t_L g2508 ( 
.A1(n_2297),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.Y(n_2508)
);

AO22x1_ASAP7_75t_L g2509 ( 
.A1(n_2297),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2242),
.Y(n_2510)
);

OA22x2_ASAP7_75t_L g2511 ( 
.A1(n_2297),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.Y(n_2511)
);

OAI22x1_ASAP7_75t_L g2512 ( 
.A1(n_2297),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2346),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2463),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2464),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2473),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2360),
.B(n_557),
.Y(n_2517)
);

AOI322xp5_ASAP7_75t_L g2518 ( 
.A1(n_2395),
.A2(n_559),
.A3(n_560),
.B1(n_561),
.B2(n_562),
.C1(n_563),
.C2(n_564),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2476),
.Y(n_2519)
);

AOI22xp5_ASAP7_75t_SL g2520 ( 
.A1(n_2442),
.A2(n_2445),
.B1(n_2439),
.B2(n_2459),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2478),
.Y(n_2521)
);

AOI322xp5_ASAP7_75t_L g2522 ( 
.A1(n_2393),
.A2(n_559),
.A3(n_560),
.B1(n_561),
.B2(n_563),
.C1(n_564),
.C2(n_565),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2479),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2484),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2488),
.Y(n_2525)
);

INVxp67_ASAP7_75t_SL g2526 ( 
.A(n_2437),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2506),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2348),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2362),
.Y(n_2529)
);

INVxp67_ASAP7_75t_SL g2530 ( 
.A(n_2440),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2366),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2391),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2354),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2381),
.Y(n_2534)
);

OA22x2_ASAP7_75t_L g2535 ( 
.A1(n_2355),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_2535)
);

AOI322xp5_ASAP7_75t_L g2536 ( 
.A1(n_2450),
.A2(n_567),
.A3(n_568),
.B1(n_570),
.B2(n_571),
.C1(n_572),
.C2(n_573),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2474),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2505),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2507),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2350),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2456),
.Y(n_2541)
);

OAI322xp33_ASAP7_75t_L g2542 ( 
.A1(n_2451),
.A2(n_570),
.A3(n_571),
.B1(n_572),
.B2(n_573),
.C1(n_574),
.C2(n_575),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_2469),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2480),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2377),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2365),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2431),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2423),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2392),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2397),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2404),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2406),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2368),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2347),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2430),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2416),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2457),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2384),
.Y(n_2558)
);

OAI322xp33_ASAP7_75t_L g2559 ( 
.A1(n_2434),
.A2(n_576),
.A3(n_577),
.B1(n_578),
.B2(n_579),
.C1(n_580),
.C2(n_581),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2369),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2420),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2417),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2465),
.Y(n_2563)
);

BUFx2_ASAP7_75t_L g2564 ( 
.A(n_2477),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2424),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2426),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2401),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2411),
.Y(n_2568)
);

INVxp67_ASAP7_75t_SL g2569 ( 
.A(n_2349),
.Y(n_2569)
);

INVx5_ASAP7_75t_SL g2570 ( 
.A(n_2400),
.Y(n_2570)
);

INVxp67_ASAP7_75t_SL g2571 ( 
.A(n_2357),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2421),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2387),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2435),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2472),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2399),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2433),
.Y(n_2577)
);

HB1xp67_ASAP7_75t_L g2578 ( 
.A(n_2386),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2487),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2495),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2510),
.Y(n_2581)
);

OAI322xp33_ASAP7_75t_L g2582 ( 
.A1(n_2454),
.A2(n_577),
.A3(n_578),
.B1(n_580),
.B2(n_581),
.C1(n_582),
.C2(n_583),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2402),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2432),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2455),
.Y(n_2585)
);

INVx2_ASAP7_75t_SL g2586 ( 
.A(n_2398),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2403),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2388),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2438),
.Y(n_2589)
);

BUFx2_ASAP7_75t_L g2590 ( 
.A(n_2383),
.Y(n_2590)
);

XNOR2x2_ASAP7_75t_L g2591 ( 
.A(n_2409),
.B(n_582),
.Y(n_2591)
);

CKINVDCx20_ASAP7_75t_R g2592 ( 
.A(n_2446),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2353),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2353),
.Y(n_2594)
);

BUFx2_ASAP7_75t_L g2595 ( 
.A(n_2458),
.Y(n_2595)
);

BUFx2_ASAP7_75t_L g2596 ( 
.A(n_2467),
.Y(n_2596)
);

INVx1_ASAP7_75t_SL g2597 ( 
.A(n_2501),
.Y(n_2597)
);

OAI322xp33_ASAP7_75t_L g2598 ( 
.A1(n_2453),
.A2(n_584),
.A3(n_585),
.B1(n_586),
.B2(n_587),
.C1(n_588),
.C2(n_589),
.Y(n_2598)
);

OAI322xp33_ASAP7_75t_L g2599 ( 
.A1(n_2441),
.A2(n_584),
.A3(n_585),
.B1(n_586),
.B2(n_587),
.C1(n_588),
.C2(n_589),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2408),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2380),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2351),
.Y(n_2602)
);

INVx5_ASAP7_75t_L g2603 ( 
.A(n_2379),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2418),
.Y(n_2604)
);

OAI322xp33_ASAP7_75t_L g2605 ( 
.A1(n_2425),
.A2(n_590),
.A3(n_591),
.B1(n_592),
.B2(n_593),
.C1(n_594),
.C2(n_595),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2409),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2385),
.Y(n_2607)
);

INVxp67_ASAP7_75t_SL g2608 ( 
.A(n_2370),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2410),
.Y(n_2609)
);

INVxp67_ASAP7_75t_L g2610 ( 
.A(n_2494),
.Y(n_2610)
);

INVx2_ASAP7_75t_SL g2611 ( 
.A(n_2364),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2428),
.Y(n_2612)
);

OAI322xp33_ASAP7_75t_L g2613 ( 
.A1(n_2396),
.A2(n_590),
.A3(n_591),
.B1(n_592),
.B2(n_593),
.C1(n_594),
.C2(n_595),
.Y(n_2613)
);

INVx3_ASAP7_75t_L g2614 ( 
.A(n_2443),
.Y(n_2614)
);

INVx1_ASAP7_75t_SL g2615 ( 
.A(n_2490),
.Y(n_2615)
);

INVxp67_ASAP7_75t_L g2616 ( 
.A(n_2449),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2452),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2429),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2361),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2493),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2371),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2419),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2466),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2468),
.Y(n_2624)
);

INVx2_ASAP7_75t_SL g2625 ( 
.A(n_2444),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2470),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2475),
.Y(n_2627)
);

XNOR2x1_ASAP7_75t_L g2628 ( 
.A(n_2415),
.B(n_596),
.Y(n_2628)
);

INVx1_ASAP7_75t_SL g2629 ( 
.A(n_2512),
.Y(n_2629)
);

INVxp67_ASAP7_75t_SL g2630 ( 
.A(n_2483),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2485),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2489),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2496),
.Y(n_2633)
);

OAI322xp33_ASAP7_75t_L g2634 ( 
.A1(n_2447),
.A2(n_596),
.A3(n_597),
.B1(n_598),
.B2(n_599),
.C1(n_600),
.C2(n_601),
.Y(n_2634)
);

INVxp67_ASAP7_75t_SL g2635 ( 
.A(n_2497),
.Y(n_2635)
);

INVxp67_ASAP7_75t_L g2636 ( 
.A(n_2604),
.Y(n_2636)
);

AOI22xp5_ASAP7_75t_L g2637 ( 
.A1(n_2530),
.A2(n_2606),
.B1(n_2595),
.B2(n_2596),
.Y(n_2637)
);

NOR4xp25_ASAP7_75t_L g2638 ( 
.A(n_2582),
.B(n_2407),
.C(n_2412),
.D(n_2427),
.Y(n_2638)
);

AOI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2630),
.A2(n_2511),
.B1(n_2499),
.B2(n_2503),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2548),
.Y(n_2640)
);

AOI22x1_ASAP7_75t_L g2641 ( 
.A1(n_2590),
.A2(n_2382),
.B1(n_2413),
.B2(n_2422),
.Y(n_2641)
);

AOI22xp5_ASAP7_75t_L g2642 ( 
.A1(n_2635),
.A2(n_2504),
.B1(n_2508),
.B2(n_2498),
.Y(n_2642)
);

AO22x2_ASAP7_75t_L g2643 ( 
.A1(n_2526),
.A2(n_2461),
.B1(n_2378),
.B2(n_2460),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2513),
.Y(n_2644)
);

AOI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2610),
.A2(n_2376),
.B1(n_2363),
.B2(n_2374),
.Y(n_2645)
);

OAI322xp33_ASAP7_75t_L g2646 ( 
.A1(n_2591),
.A2(n_2356),
.A3(n_2414),
.B1(n_2352),
.B2(n_2358),
.C1(n_2471),
.C2(n_2359),
.Y(n_2646)
);

AOI221xp5_ASAP7_75t_L g2647 ( 
.A1(n_2569),
.A2(n_2502),
.B1(n_2482),
.B2(n_2509),
.C(n_2486),
.Y(n_2647)
);

OAI322xp33_ASAP7_75t_L g2648 ( 
.A1(n_2520),
.A2(n_2367),
.A3(n_2372),
.B1(n_2373),
.B2(n_2375),
.C1(n_2390),
.C2(n_2405),
.Y(n_2648)
);

AOI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2633),
.A2(n_2481),
.B1(n_2389),
.B2(n_2448),
.Y(n_2649)
);

AOI31xp33_ASAP7_75t_L g2650 ( 
.A1(n_2619),
.A2(n_2492),
.A3(n_2491),
.B(n_2462),
.Y(n_2650)
);

AOI221xp5_ASAP7_75t_L g2651 ( 
.A1(n_2593),
.A2(n_2394),
.B1(n_2500),
.B2(n_2436),
.C(n_600),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2514),
.Y(n_2652)
);

OAI22x1_ASAP7_75t_SL g2653 ( 
.A1(n_2603),
.A2(n_601),
.B1(n_597),
.B2(n_599),
.Y(n_2653)
);

AOI22x1_ASAP7_75t_L g2654 ( 
.A1(n_2597),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2515),
.Y(n_2655)
);

AO22x2_ASAP7_75t_L g2656 ( 
.A1(n_2594),
.A2(n_2583),
.B1(n_2629),
.B2(n_2608),
.Y(n_2656)
);

INVx2_ASAP7_75t_SL g2657 ( 
.A(n_2578),
.Y(n_2657)
);

AOI22xp5_ASAP7_75t_SL g2658 ( 
.A1(n_2621),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_2658)
);

OAI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2603),
.A2(n_632),
.B1(n_629),
.B2(n_630),
.Y(n_2659)
);

AOI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2622),
.A2(n_636),
.B1(n_634),
.B2(n_635),
.Y(n_2660)
);

INVxp67_ASAP7_75t_L g2661 ( 
.A(n_2555),
.Y(n_2661)
);

HB1xp67_ASAP7_75t_L g2662 ( 
.A(n_2616),
.Y(n_2662)
);

AOI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2571),
.A2(n_639),
.B1(n_637),
.B2(n_638),
.Y(n_2663)
);

AOI221xp5_ASAP7_75t_L g2664 ( 
.A1(n_2598),
.A2(n_643),
.B1(n_640),
.B2(n_642),
.C(n_644),
.Y(n_2664)
);

OAI22xp5_ASAP7_75t_SL g2665 ( 
.A1(n_2603),
.A2(n_648),
.B1(n_645),
.B2(n_646),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2516),
.Y(n_2666)
);

AO22x2_ASAP7_75t_L g2667 ( 
.A1(n_2587),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2519),
.Y(n_2668)
);

AOI221xp5_ASAP7_75t_L g2669 ( 
.A1(n_2542),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.C(n_656),
.Y(n_2669)
);

BUFx4_ASAP7_75t_R g2670 ( 
.A(n_2589),
.Y(n_2670)
);

BUFx2_ASAP7_75t_L g2671 ( 
.A(n_2543),
.Y(n_2671)
);

NAND4xp75_ASAP7_75t_L g2672 ( 
.A(n_2611),
.B(n_659),
.C(n_657),
.D(n_658),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2586),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2521),
.Y(n_2674)
);

AO22x2_ASAP7_75t_L g2675 ( 
.A1(n_2585),
.A2(n_663),
.B1(n_660),
.B2(n_661),
.Y(n_2675)
);

OAI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2625),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.Y(n_2676)
);

NAND4xp25_ASAP7_75t_L g2677 ( 
.A(n_2518),
.B(n_669),
.C(n_667),
.D(n_668),
.Y(n_2677)
);

AOI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2614),
.A2(n_673),
.B1(n_670),
.B2(n_671),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2523),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2524),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2525),
.Y(n_2681)
);

INVx2_ASAP7_75t_SL g2682 ( 
.A(n_2564),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2527),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2529),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2531),
.Y(n_2685)
);

OAI322xp33_ASAP7_75t_L g2686 ( 
.A1(n_2601),
.A2(n_674),
.A3(n_677),
.B1(n_678),
.B2(n_679),
.C1(n_680),
.C2(n_681),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2554),
.A2(n_2624),
.B1(n_2627),
.B2(n_2626),
.Y(n_2687)
);

AOI22xp5_ASAP7_75t_L g2688 ( 
.A1(n_2632),
.A2(n_686),
.B1(n_683),
.B2(n_685),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2592),
.Y(n_2689)
);

AND4x1_ASAP7_75t_L g2690 ( 
.A(n_2600),
.B(n_689),
.C(n_687),
.D(n_688),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2532),
.Y(n_2691)
);

AO22x1_ASAP7_75t_L g2692 ( 
.A1(n_2609),
.A2(n_809),
.B1(n_697),
.B2(n_690),
.Y(n_2692)
);

AOI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2528),
.A2(n_700),
.B1(n_695),
.B2(n_698),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2662),
.Y(n_2694)
);

AOI221xp5_ASAP7_75t_L g2695 ( 
.A1(n_2656),
.A2(n_2599),
.B1(n_2613),
.B2(n_2634),
.C(n_2605),
.Y(n_2695)
);

INVxp67_ASAP7_75t_SL g2696 ( 
.A(n_2653),
.Y(n_2696)
);

NOR2x1_ASAP7_75t_L g2697 ( 
.A(n_2671),
.B(n_2628),
.Y(n_2697)
);

AOI22xp33_ASAP7_75t_L g2698 ( 
.A1(n_2643),
.A2(n_2584),
.B1(n_2617),
.B2(n_2546),
.Y(n_2698)
);

OAI221xp5_ASAP7_75t_L g2699 ( 
.A1(n_2637),
.A2(n_2620),
.B1(n_2615),
.B2(n_2561),
.C(n_2623),
.Y(n_2699)
);

INVxp67_ASAP7_75t_L g2700 ( 
.A(n_2689),
.Y(n_2700)
);

OAI22xp5_ASAP7_75t_L g2701 ( 
.A1(n_2639),
.A2(n_2631),
.B1(n_2607),
.B2(n_2602),
.Y(n_2701)
);

O2A1O1Ixp33_ASAP7_75t_L g2702 ( 
.A1(n_2650),
.A2(n_2517),
.B(n_2559),
.C(n_2618),
.Y(n_2702)
);

AOI22x1_ASAP7_75t_L g2703 ( 
.A1(n_2643),
.A2(n_2544),
.B1(n_2541),
.B2(n_2537),
.Y(n_2703)
);

A2O1A1Ixp33_ASAP7_75t_SL g2704 ( 
.A1(n_2636),
.A2(n_2538),
.B(n_2539),
.C(n_2534),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2640),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2656),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2642),
.A2(n_2612),
.B1(n_2535),
.B2(n_2553),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2661),
.Y(n_2708)
);

AOI22xp5_ASAP7_75t_L g2709 ( 
.A1(n_2647),
.A2(n_2588),
.B1(n_2573),
.B2(n_2563),
.Y(n_2709)
);

AOI221xp5_ASAP7_75t_L g2710 ( 
.A1(n_2638),
.A2(n_2560),
.B1(n_2579),
.B2(n_2581),
.C(n_2580),
.Y(n_2710)
);

OAI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2645),
.A2(n_2570),
.B1(n_2557),
.B2(n_2575),
.Y(n_2711)
);

AOI221xp5_ASAP7_75t_L g2712 ( 
.A1(n_2648),
.A2(n_2566),
.B1(n_2558),
.B2(n_2556),
.C(n_2552),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2644),
.Y(n_2713)
);

AOI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2651),
.A2(n_2577),
.B1(n_2574),
.B2(n_2567),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2652),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_2682),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2670),
.Y(n_2717)
);

AOI211xp5_ASAP7_75t_SL g2718 ( 
.A1(n_2646),
.A2(n_2576),
.B(n_2565),
.C(n_2572),
.Y(n_2718)
);

AND4x1_ASAP7_75t_L g2719 ( 
.A(n_2664),
.B(n_2568),
.C(n_2562),
.D(n_2547),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2655),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2666),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2668),
.Y(n_2722)
);

AOI31xp33_ASAP7_75t_L g2723 ( 
.A1(n_2658),
.A2(n_2533),
.A3(n_2545),
.B(n_2540),
.Y(n_2723)
);

NAND4xp25_ASAP7_75t_L g2724 ( 
.A(n_2687),
.B(n_2522),
.C(n_2536),
.D(n_2549),
.Y(n_2724)
);

OAI221xp5_ASAP7_75t_L g2725 ( 
.A1(n_2649),
.A2(n_2551),
.B1(n_2550),
.B2(n_2570),
.C(n_703),
.Y(n_2725)
);

NOR4xp25_ASAP7_75t_L g2726 ( 
.A(n_2699),
.B(n_2657),
.C(n_2673),
.D(n_2674),
.Y(n_2726)
);

NOR2x1_ASAP7_75t_L g2727 ( 
.A(n_2697),
.B(n_2706),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2694),
.Y(n_2728)
);

AO22x2_ASAP7_75t_L g2729 ( 
.A1(n_2707),
.A2(n_2679),
.B1(n_2681),
.B2(n_2680),
.Y(n_2729)
);

AOI22xp5_ASAP7_75t_L g2730 ( 
.A1(n_2696),
.A2(n_2665),
.B1(n_2677),
.B2(n_2669),
.Y(n_2730)
);

AOI22xp5_ASAP7_75t_L g2731 ( 
.A1(n_2695),
.A2(n_2659),
.B1(n_2660),
.B2(n_2688),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2708),
.Y(n_2732)
);

HB1xp67_ASAP7_75t_L g2733 ( 
.A(n_2717),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2705),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2700),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2716),
.B(n_2641),
.Y(n_2736)
);

INVxp67_ASAP7_75t_L g2737 ( 
.A(n_2723),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2713),
.Y(n_2738)
);

AOI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2724),
.A2(n_2676),
.B1(n_2672),
.B2(n_2663),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2703),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2715),
.Y(n_2741)
);

AO22x2_ASAP7_75t_L g2742 ( 
.A1(n_2701),
.A2(n_2683),
.B1(n_2685),
.B2(n_2684),
.Y(n_2742)
);

NOR2x1_ASAP7_75t_L g2743 ( 
.A(n_2725),
.B(n_2691),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2720),
.Y(n_2744)
);

OAI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2737),
.A2(n_2714),
.B1(n_2698),
.B2(n_2709),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2733),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2735),
.Y(n_2747)
);

AOI22xp5_ASAP7_75t_L g2748 ( 
.A1(n_2740),
.A2(n_2711),
.B1(n_2710),
.B2(n_2712),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2726),
.B(n_2718),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2727),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_SL g2751 ( 
.A(n_2730),
.B(n_2719),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2728),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2732),
.Y(n_2753)
);

INVxp67_ASAP7_75t_L g2754 ( 
.A(n_2742),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_2750),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2745),
.B(n_2736),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2749),
.A2(n_2729),
.B1(n_2731),
.B2(n_2739),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2746),
.B(n_2702),
.Y(n_2758)
);

OAI22xp5_ASAP7_75t_SL g2759 ( 
.A1(n_2748),
.A2(n_2743),
.B1(n_2734),
.B2(n_2741),
.Y(n_2759)
);

NOR4xp25_ASAP7_75t_L g2760 ( 
.A(n_2754),
.B(n_2744),
.C(n_2738),
.D(n_2721),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2747),
.Y(n_2761)
);

INVx2_ASAP7_75t_SL g2762 ( 
.A(n_2752),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2753),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2755),
.Y(n_2764)
);

HB1xp67_ASAP7_75t_L g2765 ( 
.A(n_2762),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2758),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2761),
.Y(n_2767)
);

HB1xp67_ASAP7_75t_L g2768 ( 
.A(n_2759),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2763),
.Y(n_2769)
);

NAND4xp25_ASAP7_75t_L g2770 ( 
.A(n_2766),
.B(n_2757),
.C(n_2756),
.D(n_2751),
.Y(n_2770)
);

AOI22xp5_ASAP7_75t_L g2771 ( 
.A1(n_2768),
.A2(n_2722),
.B1(n_2760),
.B2(n_2692),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2765),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2772),
.Y(n_2773)
);

AOI22xp33_ASAP7_75t_SL g2774 ( 
.A1(n_2773),
.A2(n_2764),
.B1(n_2654),
.B2(n_2767),
.Y(n_2774)
);

INVxp67_ASAP7_75t_SL g2775 ( 
.A(n_2774),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2775),
.A2(n_2771),
.B1(n_2770),
.B2(n_2769),
.Y(n_2776)
);

INVxp67_ASAP7_75t_L g2777 ( 
.A(n_2776),
.Y(n_2777)
);

AOI221xp5_ASAP7_75t_L g2778 ( 
.A1(n_2777),
.A2(n_2704),
.B1(n_2667),
.B2(n_2675),
.C(n_2686),
.Y(n_2778)
);

AOI211xp5_ASAP7_75t_L g2779 ( 
.A1(n_2778),
.A2(n_2678),
.B(n_2693),
.C(n_2690),
.Y(n_2779)
);


endmodule