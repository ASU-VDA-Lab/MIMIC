module fake_ariane_2121_n_7880 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_702, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_7880);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_702;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_7880;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_7832;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_7805;
wire n_2790;
wire n_7542;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6358;
wire n_6293;
wire n_2482;
wire n_1682;
wire n_7001;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_4260;
wire n_903;
wire n_7626;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_7368;
wire n_1690;
wire n_2807;
wire n_6664;
wire n_7562;
wire n_7534;
wire n_1018;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_4132;
wire n_1364;
wire n_7373;
wire n_2390;
wire n_6891;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_6539;
wire n_4824;
wire n_7467;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_7526;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_786;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_7200;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_5691;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_863;
wire n_6992;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_899;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_6681;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_5092;
wire n_2456;
wire n_1924;
wire n_6542;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_7507;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_1213;
wire n_2382;
wire n_7379;
wire n_7441;
wire n_780;
wire n_5292;
wire n_1918;
wire n_7438;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_5843;
wire n_7874;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_7695;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_6872;
wire n_6644;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_7607;
wire n_7642;
wire n_1386;
wire n_6236;
wire n_7104;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_7259;
wire n_7838;
wire n_5984;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_7840;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_6624;
wire n_1357;
wire n_6710;
wire n_6883;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_4033;
wire n_2659;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_6261;
wire n_6659;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_7583;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_2954;
wire n_4438;
wire n_6538;
wire n_974;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7599;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_5708;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_3147;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_1247;
wire n_6860;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_6382;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_6615;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_720;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_5985;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_7868;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_7176;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_7547;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_7527;
wire n_4856;
wire n_2618;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_6482;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_3070;
wire n_1005;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_7869;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_6631;
wire n_5889;
wire n_7151;
wire n_3944;
wire n_7762;
wire n_5632;
wire n_4729;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_7611;
wire n_7796;
wire n_6508;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_2211;
wire n_951;
wire n_7546;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_722;
wire n_7407;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_2958;
wire n_7481;
wire n_1044;
wire n_4429;
wire n_6484;
wire n_5435;
wire n_1714;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_5476;
wire n_5483;
wire n_7605;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_6639;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_7736;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_811;
wire n_6600;
wire n_7010;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_7346;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_5077;
wire n_6102;
wire n_1874;
wire n_3780;
wire n_1657;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_1330;
wire n_906;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_7148;
wire n_3142;
wire n_7169;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_7600;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_6946;
wire n_5931;
wire n_1829;
wire n_4635;
wire n_7847;
wire n_1450;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_7660;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6442;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_6840;
wire n_6645;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_7831;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_7455;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_7509;
wire n_6205;
wire n_2506;
wire n_4825;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_7497;
wire n_7315;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_6706;
wire n_7431;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_7521;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_1291;
wire n_7253;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_7569;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_7505;
wire n_3921;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_7573;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_7498;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_3822;
wire n_889;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_6141;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_7240;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_1056;
wire n_5584;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6248;
wire n_6541;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_4733;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_6351;
wire n_4509;
wire n_4935;
wire n_2073;
wire n_7382;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_7510;
wire n_3786;
wire n_875;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_7691;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_6744;
wire n_3645;
wire n_793;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_6116;
wire n_3550;
wire n_5510;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_3610;
wire n_2443;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_7671;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_7528;
wire n_6209;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_7413;
wire n_7821;
wire n_7620;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_1775;
wire n_908;
wire n_1036;
wire n_7109;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_6716;
wire n_3565;
wire n_6905;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_7817;
wire n_6413;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_1261;
wire n_7249;
wire n_5763;
wire n_3633;
wire n_857;
wire n_6061;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_7297;
wire n_7730;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_2324;
wire n_840;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_7140;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_3303;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_7741;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_6668;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_7698;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_4266;
wire n_6336;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_5399;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_7747;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_7650;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_708;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_4548;
wire n_7819;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_774;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_7794;
wire n_1705;
wire n_768;
wire n_3707;
wire n_3895;
wire n_1091;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_7630;
wire n_4161;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_1581;
wire n_946;
wire n_3058;
wire n_5355;
wire n_757;
wire n_2047;
wire n_1655;
wire n_3398;
wire n_1146;
wire n_3709;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_5915;
wire n_7276;
wire n_6379;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_7753;
wire n_6834;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_719;
wire n_7541;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7841;
wire n_7160;
wire n_7324;
wire n_6046;
wire n_7054;
wire n_1233;
wire n_4493;
wire n_6055;
wire n_7161;
wire n_1808;
wire n_6364;
wire n_6091;
wire n_6348;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_886;
wire n_7837;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_7676;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_7644;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_7879;
wire n_6607;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_829;
wire n_4814;
wire n_6178;
wire n_6677;
wire n_2221;
wire n_7875;
wire n_5502;
wire n_1283;
wire n_7550;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_7238;
wire n_6862;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_7804;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_1276;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_7826;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_3999;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_4576;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_6935;
wire n_2899;
wire n_1560;
wire n_6984;
wire n_6778;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_6386;
wire n_2722;
wire n_3728;
wire n_6596;
wire n_5107;
wire n_7165;
wire n_4680;
wire n_5067;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_772;
wire n_6741;
wire n_1245;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_2969;
wire n_3429;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_6947;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_912;
wire n_6375;
wire n_7781;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_2855;
wire n_794;
wire n_2848;
wire n_7675;
wire n_6775;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_7774;
wire n_6970;
wire n_1026;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_7873;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_1399;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_2224;
wire n_1226;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_6390;
wire n_7640;
wire n_2302;
wire n_6799;
wire n_3014;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_5661;
wire n_3760;
wire n_7641;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_7764;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_7520;
wire n_5314;
wire n_7616;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_7235;
wire n_2511;
wire n_6572;
wire n_3981;
wire n_7271;
wire n_2681;
wire n_7222;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_6387;
wire n_4201;
wire n_6470;
wire n_7206;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_7854;
wire n_926;
wire n_2296;
wire n_5735;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_7533;
wire n_3377;
wire n_6722;
wire n_1518;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_1287;
wire n_1611;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_7436;
wire n_7020;
wire n_5935;
wire n_6696;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_5488;
wire n_1105;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1614;
wire n_1377;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_7465;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_729;
wire n_6222;
wire n_2218;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_6969;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_6587;
wire n_6688;
wire n_6505;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_3908;
wire n_6453;
wire n_6308;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_7449;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_3216;
wire n_3568;
wire n_2555;
wire n_2708;
wire n_6187;
wire n_735;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_7479;
wire n_1649;
wire n_2470;
wire n_7517;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_6547;
wire n_7177;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_6478;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_6906;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3669;
wire n_3367;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_7818;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_7862;
wire n_3735;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_7721;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_6999;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_6440;
wire n_4977;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_5936;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_7348;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_6464;
wire n_5129;
wire n_806;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_6850;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_7743;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_6550;
wire n_6656;
wire n_6972;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_3317;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_7035;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_7442;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_6258;
wire n_1288;
wire n_7715;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_7699;
wire n_1153;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_5911;
wire n_7340;
wire n_3600;
wire n_7303;
wire n_1023;
wire n_914;
wire n_7870;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_7207;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_7618;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_7633;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_2592;
wire n_3490;
wire n_7280;
wire n_962;
wire n_5043;
wire n_7339;
wire n_7597;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_5645;
wire n_5020;
wire n_6455;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6183;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_4256;
wire n_2560;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_7612;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_2150;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_6695;
wire n_7529;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_3807;
wire n_2951;
wire n_4048;
wire n_6213;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_7101;
wire n_1204;
wire n_7843;
wire n_994;
wire n_2428;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_7578;
wire n_3410;
wire n_5415;
wire n_856;
wire n_7261;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_6993;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_6755;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7310;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_7514;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_6105;
wire n_826;
wire n_5512;
wire n_7738;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_7609;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_7282;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_6331;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_6023;
wire n_7820;
wire n_816;
wire n_7833;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_7750;
wire n_5057;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_7697;
wire n_5887;
wire n_7808;
wire n_3068;
wire n_1629;
wire n_7603;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_6450;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_1236;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_2048;
wire n_7723;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_838;
wire n_1941;
wire n_7045;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_7777;
wire n_4258;
wire n_5756;
wire n_7693;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_7682;
wire n_7300;
wire n_1410;
wire n_939;
wire n_6861;
wire n_2297;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_7798;
wire n_4767;
wire n_4569;
wire n_948;
wire n_6528;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_7672;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_6885;
wire n_7681;
wire n_5039;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_4265;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_7491;
wire n_1583;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_7150;
wire n_1264;
wire n_6602;
wire n_6530;
wire n_4958;
wire n_1827;
wire n_4149;
wire n_6135;
wire n_2361;
wire n_1752;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_7336;
wire n_5932;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_7493;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_5823;
wire n_2423;
wire n_2208;
wire n_1421;
wire n_5422;
wire n_5944;
wire n_6989;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_1069;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_7273;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_6758;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_7601;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_5294;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1187;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_7138;
wire n_766;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_7617;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_7700;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_6654;
wire n_7661;
wire n_4968;
wire n_7801;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_5316;
wire n_7876;
wire n_2735;
wire n_953;
wire n_4214;
wire n_5290;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_7323;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_795;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_4176;
wire n_7556;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_6691;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_6771;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_5718;
wire n_1461;
wire n_7208;
wire n_7718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_5658;
wire n_1112;
wire n_4174;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_5610;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1468;
wire n_1253;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_7289;
wire n_7538;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_6533;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_7483;
wire n_5710;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_3510;
wire n_7046;
wire n_7834;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_6357;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_7811;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_6713;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_6108;
wire n_7664;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_5862;
wire n_7477;
wire n_1914;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_7714;
wire n_6415;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_7858;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6513;
wire n_6392;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_7680;
wire n_5630;
wire n_6666;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_7710;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_7061;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_7783;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_4728;
wire n_7171;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_3968;
wire n_1365;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_7501;
wire n_6432;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_7589;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_3983;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_7511;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_6957;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_6694;
wire n_3260;
wire n_2496;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_3139;
wire n_5681;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_7621;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_7572;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_6662;
wire n_7494;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_6433;
wire n_1763;
wire n_6200;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_2660;
wire n_3426;
wire n_1859;
wire n_6902;
wire n_4615;
wire n_3492;
wire n_3044;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_5657;
wire n_3579;
wire n_2379;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_6956;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_5420;
wire n_6497;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_4387;
wire n_1711;
wire n_2508;
wire n_3186;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_7032;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_7752;
wire n_5081;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_6362;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_7126;
wire n_5867;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_7518;
wire n_4385;
wire n_7779;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_1786;
wire n_6309;
wire n_3732;
wire n_1804;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_1318;
wire n_1769;
wire n_1632;
wire n_7349;
wire n_1929;
wire n_4319;
wire n_6585;
wire n_7786;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_7579;
wire n_7122;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_7624;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_7828;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_7543;
wire n_5475;
wire n_7727;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_7019;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_7702;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_6685;
wire n_756;
wire n_3390;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_4666;
wire n_3140;
wire n_2320;
wire n_4082;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_7347;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_1659;
wire n_3955;
wire n_885;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_3336;
wire n_7739;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_6549;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7610;
wire n_7107;
wire n_4561;
wire n_3291;
wire n_1541;
wire n_7456;
wire n_7369;
wire n_1472;
wire n_1050;
wire n_7548;
wire n_2578;
wire n_1201;
wire n_7598;
wire n_2475;
wire n_1185;
wire n_7250;
wire n_7823;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_1090;
wire n_4536;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_7525;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_6923;
wire n_7649;
wire n_843;
wire n_3358;
wire n_6704;
wire n_7634;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_4682;
wire n_1128;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_7844;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_7009;
wire n_3376;
wire n_7371;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_7463;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5755;
wire n_5700;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_4711;
wire n_2553;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_6184;
wire n_1767;
wire n_4138;
wire n_3131;
wire n_1040;
wire n_7083;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_6312;
wire n_7683;
wire n_2154;
wire n_7669;
wire n_1986;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_7330;
wire n_6007;
wire n_6734;
wire n_6535;
wire n_1772;
wire n_6879;
wire n_1311;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_6457;
wire n_4924;
wire n_4044;
wire n_6270;
wire n_2305;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7082;
wire n_7237;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_7042;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_3178;
wire n_7023;
wire n_2251;
wire n_5842;
wire n_5758;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_7787;
wire n_7836;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_6764;
wire n_7871;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_6955;
wire n_7563;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_6569;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_3897;
wire n_7103;
wire n_6605;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_6832;
wire n_5980;
wire n_956;
wire n_4092;
wire n_765;
wire n_4875;
wire n_7771;
wire n_4255;
wire n_2758;
wire n_6544;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_7133;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_6289;
wire n_6651;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_7706;
wire n_7813;
wire n_2420;
wire n_7643;
wire n_6836;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_835;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_7628;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_839;
wire n_1754;
wire n_7236;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_6786;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7519;
wire n_7802;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_2933;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_6214;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_6945;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_977;
wire n_2339;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_7674;
wire n_6175;
wire n_6445;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_6499;
wire n_1982;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_7361;
wire n_1114;
wire n_4679;
wire n_1742;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_3504;
wire n_2587;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_6732;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_7646;
wire n_3779;
wire n_6982;
wire n_1063;
wire n_7291;
wire n_991;
wire n_2275;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_7017;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_7861;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_7554;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_7648;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_7653;
wire n_6400;
wire n_1644;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_7551;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_6621;
wire n_6851;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_7606;
wire n_7420;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_7319;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_7516;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_7244;
wire n_1463;
wire n_4626;
wire n_7625;
wire n_4997;
wire n_5065;
wire n_6806;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_7857;
wire n_2461;
wire n_1706;
wire n_3719;
wire n_7154;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_7068;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_7864;
wire n_3451;
wire n_4734;
wire n_6675;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_7384;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_7761;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_1544;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_7859;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_7523;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_7559;
wire n_7576;
wire n_6988;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_7081;
wire n_7742;
wire n_5253;
wire n_3588;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_4775;
wire n_1442;
wire n_6256;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_7264;
wire n_7842;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_7492;
wire n_804;
wire n_6649;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_955;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_6431;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_824;
wire n_5659;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_7793;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_7746;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_7570;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_6473;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_6857;
wire n_1455;
wire n_2287;
wire n_3415;
wire n_836;
wire n_6975;
wire n_7763;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_7703;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_6622;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_7665;
wire n_5262;
wire n_7677;
wire n_3262;
wire n_5319;
wire n_927;
wire n_7469;
wire n_3699;
wire n_6118;
wire n_2120;
wire n_706;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_4725;
wire n_2168;
wire n_2757;
wire n_2404;
wire n_2312;
wire n_7203;
wire n_7797;
wire n_1826;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_7111;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_6617;
wire n_7725;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2027;
wire n_2932;
wire n_6217;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3922;
wire n_3039;
wire n_2195;
wire n_5455;
wire n_6777;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_4889;
wire n_2159;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_7365;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_5022;
wire n_6370;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_3009;
wire n_777;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_6712;
wire n_7530;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_7471;
wire n_6465;
wire n_5673;
wire n_861;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_3326;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_7581;
wire n_1222;
wire n_7139;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_4463;
wire n_5357;
wire n_7173;
wire n_3648;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_6667;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_6305;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7751;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_7591;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_7444;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_2071;
wire n_7426;
wire n_3953;
wire n_4400;
wire n_7502;
wire n_2414;
wire n_5434;
wire n_2959;
wire n_2082;
wire n_1532;
wire n_6855;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_7252;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_7065;
wire n_1466;
wire n_6177;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_7367;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_4035;
wire n_6952;
wire n_1480;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_7685;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_7619;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_5577;
wire n_876;
wire n_5872;
wire n_6692;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_3694;
wire n_6854;
wire n_771;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_7537;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_819;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_3543;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_6377;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_7765;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_7815;
wire n_1052;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_7785;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_7728;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_7181;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_928;
wire n_3769;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_748;
wire n_7089;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_5868;
wire n_6417;
wire n_7145;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_7803;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_7622;
wire n_7839;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_1356;
wire n_6831;
wire n_1773;
wire n_4544;
wire n_3175;
wire n_2666;
wire n_5578;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_7564;
wire n_5863;
wire n_6633;
wire n_3790;
wire n_7775;
wire n_907;
wire n_7118;
wire n_6152;
wire n_5734;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_7636;
wire n_4341;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_6428;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_7666;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_5977;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_7262;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_3310;
wire n_4423;
wire n_2642;
wire n_3689;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_763;
wire n_6301;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_6282;
wire n_4934;
wire n_7686;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_6737;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_6448;
wire n_5186;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_7077;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_7663;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_7214;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_3989;
wire n_7652;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_7566;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_6816;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_7553;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_7086;
wire n_5689;
wire n_7732;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_1922;
wire n_940;
wire n_4877;
wire n_1537;
wire n_2065;
wire n_7038;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_7593;
wire n_898;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_5343;
wire n_6672;
wire n_7757;
wire n_1093;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_6242;
wire n_6601;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_1003;
wire n_7758;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_7439;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_7744;
wire n_3898;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_4749;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_7684;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_4238;
wire n_6371;
wire n_904;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_6264;
wire n_5782;
wire n_4168;
wire n_1369;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_7480;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_7380;
wire n_2839;
wire n_3237;
wire n_7708;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_6277;
wire n_5115;
wire n_7376;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_6409;
wire n_4095;
wire n_1310;
wire n_5927;
wire n_4485;
wire n_7657;
wire n_6388;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_6679;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_937;
wire n_1631;
wire n_7602;
wire n_6566;
wire n_1794;
wire n_5696;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_7627;
wire n_6436;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_7450;
wire n_3217;
wire n_6081;
wire n_1249;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_7582;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_7555;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_841;
wire n_3204;
wire n_7451;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_563),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_404),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_395),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_434),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_686),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_440),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_638),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_432),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_70),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_465),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_58),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_454),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_703),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_494),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_172),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_515),
.Y(n_721)
);

BUFx8_ASAP7_75t_SL g722 ( 
.A(n_517),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_25),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_230),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_590),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_3),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_336),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_275),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_650),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_184),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_341),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_262),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_105),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_419),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_652),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_426),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_258),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_618),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_566),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_458),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_138),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_196),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_34),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_68),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_443),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_550),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_691),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_311),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_632),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_272),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_139),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_576),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_308),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_481),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_0),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_609),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_217),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_478),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_242),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_631),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_655),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_230),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_315),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_284),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_115),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_344),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_519),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_578),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_605),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_680),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_342),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_691),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_268),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_639),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_281),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_624),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_18),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_565),
.Y(n_778)
);

INVxp33_ASAP7_75t_R g779 ( 
.A(n_606),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_576),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_528),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_303),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_81),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_704),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_613),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_538),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_306),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_296),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_356),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_488),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_50),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_305),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_375),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_173),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_656),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_261),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_58),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_608),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_511),
.Y(n_799)
);

CKINVDCx16_ASAP7_75t_R g800 ( 
.A(n_140),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_231),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_308),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_255),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_638),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_242),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_371),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_562),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_71),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_573),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_381),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_555),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_132),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_136),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_82),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_675),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_364),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_302),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_194),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_620),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_8),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_678),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_530),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_601),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_385),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_159),
.Y(n_825)
);

BUFx8_ASAP7_75t_SL g826 ( 
.A(n_509),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_514),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_305),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_553),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_273),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_60),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_562),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_86),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_551),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_687),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_383),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_60),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_320),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_580),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_525),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_437),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_678),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_372),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_393),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_186),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_461),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_500),
.Y(n_847)
);

HB1xp67_ASAP7_75t_SL g848 ( 
.A(n_348),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_379),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_224),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_27),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_215),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_468),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_275),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_616),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_98),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_630),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_239),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_15),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_1),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_341),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_436),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_35),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_91),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_229),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_279),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_589),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_253),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_625),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_699),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_266),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_444),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_392),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_269),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_87),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_383),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_660),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_122),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_442),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_438),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_637),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_151),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_286),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_382),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_407),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_82),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_620),
.Y(n_887)
);

BUFx2_ASAP7_75t_SL g888 ( 
.A(n_453),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_86),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_696),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_192),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_428),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_395),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_244),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_11),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_73),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_28),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_52),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_46),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_397),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_68),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_332),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_217),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_298),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_594),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_621),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_14),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_604),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_76),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_348),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_322),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_150),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_664),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_607),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_146),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_500),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_522),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_437),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_20),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_520),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_215),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_51),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_220),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_534),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_570),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_531),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_584),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_226),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_611),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_651),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_525),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_493),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_618),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_504),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_583),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_302),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_91),
.Y(n_937)
);

INVx4_ASAP7_75t_R g938 ( 
.A(n_685),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_306),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_97),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_542),
.Y(n_941)
);

CKINVDCx14_ASAP7_75t_R g942 ( 
.A(n_374),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_697),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_684),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_600),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_577),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_438),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_522),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_624),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_699),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_145),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_56),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_172),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_44),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_301),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_2),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_693),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_492),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_402),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_586),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_40),
.Y(n_961)
);

BUFx5_ASAP7_75t_L g962 ( 
.A(n_159),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_55),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_343),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_568),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_665),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_176),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_547),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_220),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_546),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_235),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_325),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_197),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_523),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_476),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_88),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_227),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_578),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_539),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_75),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_649),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_227),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_95),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_277),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_137),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_43),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_377),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_389),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_573),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_593),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_418),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_572),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_257),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_74),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_425),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_656),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_364),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_145),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_300),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_561),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_224),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_70),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_496),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_290),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_433),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_346),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_517),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_464),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_394),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_537),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_290),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_473),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_195),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_221),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_90),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_246),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_219),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_440),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_45),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_591),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_111),
.Y(n_1021)
);

CKINVDCx16_ASAP7_75t_R g1022 ( 
.A(n_102),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_553),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_535),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_463),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_148),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_84),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_704),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_6),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_622),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_219),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_568),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_28),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_642),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_502),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_245),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_29),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_418),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_608),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_304),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_488),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_468),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_249),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_546),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_448),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_477),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_48),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_112),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_486),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_483),
.Y(n_1050)
);

INVxp33_ASAP7_75t_SL g1051 ( 
.A(n_478),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_550),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_338),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_98),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_0),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_330),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_118),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_337),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_212),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_303),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_426),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_628),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_52),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_264),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_435),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_664),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_229),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_516),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_59),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_334),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_0),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_327),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_350),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_449),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_44),
.Y(n_1075)
);

BUFx10_ASAP7_75t_L g1076 ( 
.A(n_538),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_572),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_199),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_18),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_115),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_320),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_535),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_417),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_299),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_416),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_390),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_108),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_294),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_183),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_539),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_343),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_643),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_26),
.Y(n_1093)
);

BUFx10_ASAP7_75t_L g1094 ( 
.A(n_674),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_405),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_157),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_261),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_269),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_436),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_27),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_105),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_434),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_196),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_677),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_226),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_483),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_580),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_406),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_471),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_26),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_666),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_241),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_644),
.Y(n_1113)
);

BUFx10_ASAP7_75t_L g1114 ( 
.A(n_499),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_111),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_543),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_481),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_248),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_376),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_233),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_346),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_153),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_272),
.Y(n_1123)
);

BUFx10_ASAP7_75t_L g1124 ( 
.A(n_127),
.Y(n_1124)
);

CKINVDCx14_ASAP7_75t_R g1125 ( 
.A(n_180),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_422),
.Y(n_1126)
);

CKINVDCx16_ASAP7_75t_R g1127 ( 
.A(n_570),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_267),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_512),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_646),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_477),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_595),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_513),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_85),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_406),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_250),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_259),
.Y(n_1137)
);

BUFx5_ASAP7_75t_L g1138 ( 
.A(n_281),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_66),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_496),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_158),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_255),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_212),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_122),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_558),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_25),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_126),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_137),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_148),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_450),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_240),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_268),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_559),
.Y(n_1153)
);

CKINVDCx16_ASAP7_75t_R g1154 ( 
.A(n_444),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_71),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_287),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_112),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_315),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_651),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_324),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_83),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_581),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_501),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_103),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_179),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_690),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_162),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_286),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_563),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_322),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_14),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_198),
.Y(n_1172)
);

CKINVDCx14_ASAP7_75t_R g1173 ( 
.A(n_639),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_509),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_9),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_54),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_181),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_551),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_170),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_448),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_12),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_697),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_567),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_630),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_530),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_127),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_24),
.Y(n_1187)
);

BUFx2_ASAP7_75t_R g1188 ( 
.A(n_311),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_447),
.Y(n_1189)
);

BUFx10_ASAP7_75t_L g1190 ( 
.A(n_523),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_601),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_648),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_454),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_424),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_669),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_282),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_299),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_174),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_533),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_405),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_54),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_284),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_599),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_619),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_631),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_533),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_39),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_167),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_492),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_424),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_374),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_362),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_139),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_386),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_684),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_309),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_587),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_452),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_192),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_657),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_35),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_681),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_78),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_88),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_487),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_330),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_644),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_680),
.Y(n_1228)
);

CKINVDCx16_ASAP7_75t_R g1229 ( 
.A(n_80),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_606),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_695),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_511),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_247),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_534),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_602),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_50),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_18),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_411),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_435),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_382),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_513),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_625),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_675),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_187),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_294),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_564),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_526),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_271),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_962),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_746),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_962),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_962),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_962),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_962),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_962),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_962),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_962),
.Y(n_1257)
);

CKINVDCx14_ASAP7_75t_R g1258 ( 
.A(n_942),
.Y(n_1258)
);

CKINVDCx16_ASAP7_75t_R g1259 ( 
.A(n_942),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1125),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_863),
.Y(n_1261)
);

INVxp67_ASAP7_75t_SL g1262 ( 
.A(n_863),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_863),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_707),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_746),
.B(n_1),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_707),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1125),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_707),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_746),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1247),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_787),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_787),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_962),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_787),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1175),
.Y(n_1275)
);

INVxp67_ASAP7_75t_SL g1276 ( 
.A(n_1171),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_802),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1175),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1247),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_802),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_802),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_714),
.Y(n_1282)
);

INVxp33_ASAP7_75t_L g1283 ( 
.A(n_791),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_815),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_962),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_1171),
.Y(n_1286)
);

INVxp33_ASAP7_75t_SL g1287 ( 
.A(n_791),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_815),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_757),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_815),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_714),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_962),
.Y(n_1292)
);

INVxp67_ASAP7_75t_SL g1293 ( 
.A(n_1171),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_757),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1173),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1173),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_854),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_854),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_854),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_722),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_716),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_862),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_862),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_862),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_886),
.Y(n_1305)
);

INVxp33_ASAP7_75t_SL g1306 ( 
.A(n_831),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_886),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_886),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1138),
.Y(n_1309)
);

INVxp33_ASAP7_75t_SL g1310 ( 
.A(n_831),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_757),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_891),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_891),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_891),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_899),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_722),
.Y(n_1316)
);

INVxp33_ASAP7_75t_SL g1317 ( 
.A(n_858),
.Y(n_1317)
);

CKINVDCx16_ASAP7_75t_R g1318 ( 
.A(n_800),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1247),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_1171),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_899),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_716),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1171),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1138),
.Y(n_1324)
);

CKINVDCx14_ASAP7_75t_R g1325 ( 
.A(n_1221),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_899),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_733),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1138),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_936),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1221),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_1171),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1138),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1138),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1138),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1138),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1138),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1138),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_733),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1247),
.Y(n_1339)
);

NOR2xp67_ASAP7_75t_L g1340 ( 
.A(n_897),
.B(n_1),
.Y(n_1340)
);

INVxp33_ASAP7_75t_SL g1341 ( 
.A(n_858),
.Y(n_1341)
);

XNOR2xp5_ASAP7_75t_L g1342 ( 
.A(n_735),
.B(n_2),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_826),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1138),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_936),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1138),
.Y(n_1346)
);

CKINVDCx14_ASAP7_75t_R g1347 ( 
.A(n_1221),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1171),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_737),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_737),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_783),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_737),
.Y(n_1352)
);

INVxp33_ASAP7_75t_SL g1353 ( 
.A(n_879),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_897),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_897),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_764),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_764),
.Y(n_1357)
);

CKINVDCx14_ASAP7_75t_R g1358 ( 
.A(n_1221),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_764),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1247),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_803),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_803),
.Y(n_1362)
);

INVxp33_ASAP7_75t_L g1363 ( 
.A(n_879),
.Y(n_1363)
);

INVxp33_ASAP7_75t_L g1364 ( 
.A(n_884),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_803),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_813),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_813),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_782),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_813),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_828),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_828),
.Y(n_1371)
);

CKINVDCx16_ASAP7_75t_R g1372 ( 
.A(n_800),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_826),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_828),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_878),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_878),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_878),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_900),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_755),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_900),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_848),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_783),
.Y(n_1382)
);

INVxp33_ASAP7_75t_SL g1383 ( 
.A(n_884),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_900),
.Y(n_1384)
);

INVxp67_ASAP7_75t_SL g1385 ( 
.A(n_755),
.Y(n_1385)
);

INVxp67_ASAP7_75t_SL g1386 ( 
.A(n_1055),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_782),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_848),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_936),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_929),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_929),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_735),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_929),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_931),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_782),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_931),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_931),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_782),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_783),
.B(n_2),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_982),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1188),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_982),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_982),
.Y(n_1403)
);

BUFx8_ASAP7_75t_SL g1404 ( 
.A(n_829),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1022),
.Y(n_1405)
);

BUFx5_ASAP7_75t_L g1406 ( 
.A(n_996),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_996),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_756),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_996),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1001),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_782),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1001),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_756),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1022),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1188),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1001),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1009),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1009),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1009),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1135),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_829),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_860),
.Y(n_1422)
);

INVxp33_ASAP7_75t_L g1423 ( 
.A(n_920),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1135),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1135),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1145),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1145),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1055),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1127),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_829),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1145),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1215),
.Y(n_1432)
);

INVxp33_ASAP7_75t_L g1433 ( 
.A(n_920),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1215),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_782),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_782),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1215),
.Y(n_1437)
);

INVxp33_ASAP7_75t_SL g1438 ( 
.A(n_1011),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_1110),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1127),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_832),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1154),
.Y(n_1442)
);

INVxp33_ASAP7_75t_SL g1443 ( 
.A(n_1011),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_773),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_923),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_773),
.Y(n_1446)
);

CKINVDCx14_ASAP7_75t_R g1447 ( 
.A(n_1221),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1154),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_832),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_832),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1200),
.Y(n_1451)
);

CKINVDCx14_ASAP7_75t_R g1452 ( 
.A(n_712),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_873),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_873),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_835),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_873),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1200),
.Y(n_1457)
);

CKINVDCx16_ASAP7_75t_R g1458 ( 
.A(n_1229),
.Y(n_1458)
);

XOR2xp5_ASAP7_75t_L g1459 ( 
.A(n_835),
.B(n_3),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_875),
.Y(n_1460)
);

CKINVDCx16_ASAP7_75t_R g1461 ( 
.A(n_1229),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_708),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_923),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_875),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_875),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_916),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_916),
.Y(n_1467)
);

CKINVDCx16_ASAP7_75t_R g1468 ( 
.A(n_712),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_916),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1014),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1014),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_945),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_923),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_709),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1014),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_710),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1110),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_923),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1119),
.Y(n_1479)
);

INVxp67_ASAP7_75t_SL g1480 ( 
.A(n_1207),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1119),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1119),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1172),
.Y(n_1483)
);

INVxp33_ASAP7_75t_SL g1484 ( 
.A(n_1038),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1172),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1172),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_745),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_745),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1038),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_745),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_748),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_923),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_923),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_748),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_1207),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_748),
.Y(n_1496)
);

CKINVDCx16_ASAP7_75t_R g1497 ( 
.A(n_712),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_752),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_752),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_752),
.Y(n_1500)
);

INVxp33_ASAP7_75t_SL g1501 ( 
.A(n_1081),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1081),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_867),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_867),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_923),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_867),
.Y(n_1506)
);

CKINVDCx16_ASAP7_75t_R g1507 ( 
.A(n_712),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_988),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_988),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_988),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_991),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_711),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_991),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_991),
.Y(n_1514)
);

INVxp67_ASAP7_75t_SL g1515 ( 
.A(n_1237),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1080),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1080),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1080),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1176),
.Y(n_1519)
);

INVxp33_ASAP7_75t_L g1520 ( 
.A(n_1176),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1189),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1189),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1237),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_860),
.Y(n_1524)
);

CKINVDCx16_ASAP7_75t_R g1525 ( 
.A(n_712),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_812),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_986),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_945),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_945),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_839),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_977),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_977),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_977),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_984),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_839),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_984),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_984),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1000),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_713),
.Y(n_1539)
);

INVxp33_ASAP7_75t_L g1540 ( 
.A(n_724),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1000),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_888),
.Y(n_1542)
);

INVxp33_ASAP7_75t_L g1543 ( 
.A(n_724),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1000),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1070),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1070),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1070),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_715),
.Y(n_1548)
);

INVxp33_ASAP7_75t_SL g1549 ( 
.A(n_820),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1117),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1117),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1117),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1126),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1126),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1126),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1158),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1158),
.Y(n_1557)
);

INVxp33_ASAP7_75t_L g1558 ( 
.A(n_725),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1158),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1186),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1186),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1186),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1194),
.Y(n_1563)
);

INVxp33_ASAP7_75t_SL g1564 ( 
.A(n_820),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1003),
.Y(n_1565)
);

INVxp33_ASAP7_75t_L g1566 ( 
.A(n_725),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1194),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1194),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_727),
.Y(n_1569)
);

CKINVDCx16_ASAP7_75t_R g1570 ( 
.A(n_812),
.Y(n_1570)
);

INVxp33_ASAP7_75t_SL g1571 ( 
.A(n_723),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_726),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_727),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_729),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_845),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_729),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_717),
.Y(n_1577)
);

CKINVDCx16_ASAP7_75t_R g1578 ( 
.A(n_812),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_736),
.Y(n_1579)
);

INVxp67_ASAP7_75t_SL g1580 ( 
.A(n_1003),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_718),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_845),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_736),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_738),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_738),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_740),
.Y(n_1586)
);

INVx4_ASAP7_75t_R g1587 ( 
.A(n_986),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_740),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_742),
.Y(n_1589)
);

INVxp33_ASAP7_75t_L g1590 ( 
.A(n_742),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_719),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_749),
.Y(n_1592)
);

INVxp33_ASAP7_75t_SL g1593 ( 
.A(n_743),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_749),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1003),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_750),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_750),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1003),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_754),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_720),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_754),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_758),
.Y(n_1602)
);

INVxp33_ASAP7_75t_SL g1603 ( 
.A(n_777),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_758),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_721),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_760),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1003),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_760),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_762),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_762),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_763),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_763),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_768),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_768),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1003),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_728),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_770),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1003),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_770),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_771),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_771),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_887),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_772),
.Y(n_1623)
);

INVxp67_ASAP7_75t_SL g1624 ( 
.A(n_1060),
.Y(n_1624)
);

INVxp33_ASAP7_75t_SL g1625 ( 
.A(n_851),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_772),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1060),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_775),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_775),
.Y(n_1629)
);

INVxp33_ASAP7_75t_SL g1630 ( 
.A(n_859),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_776),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_776),
.Y(n_1632)
);

CKINVDCx14_ASAP7_75t_R g1633 ( 
.A(n_812),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1060),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_781),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_887),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_781),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_786),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_786),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_792),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1060),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_730),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_792),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_888),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_805),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1060),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_805),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_806),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_806),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_808),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_731),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_808),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_809),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_809),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1060),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1060),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_811),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_811),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_814),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_814),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1051),
.B(n_3),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_818),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_818),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_819),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_819),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_822),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_822),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_823),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_823),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_841),
.Y(n_1670)
);

CKINVDCx16_ASAP7_75t_R g1671 ( 
.A(n_812),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_732),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_841),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1089),
.Y(n_1674)
);

INVxp33_ASAP7_75t_L g1675 ( 
.A(n_856),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1089),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1089),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_734),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1076),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_739),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_741),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1089),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1089),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_856),
.B(n_4),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_747),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1089),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1089),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_903),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1129),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1129),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1129),
.Y(n_1691)
);

CKINVDCx20_ASAP7_75t_R g1692 ( 
.A(n_903),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_908),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1129),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1129),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1285),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1627),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1550),
.Y(n_1698)
);

INVx5_ASAP7_75t_L g1699 ( 
.A(n_1270),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1422),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1627),
.Y(n_1701)
);

AOI22x1_ASAP7_75t_SL g1702 ( 
.A1(n_1275),
.A2(n_933),
.B1(n_935),
.B2(n_908),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1270),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1282),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1381),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1270),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1389),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1330),
.B(n_1129),
.Y(n_1708)
);

AOI22x1_ASAP7_75t_SL g1709 ( 
.A1(n_1275),
.A2(n_935),
.B1(n_966),
.B2(n_933),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1259),
.B(n_1246),
.Y(n_1710)
);

INVx5_ASAP7_75t_L g1711 ( 
.A(n_1270),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1260),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_1282),
.Y(n_1713)
);

INVx5_ASAP7_75t_L g1714 ( 
.A(n_1270),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1279),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1389),
.B(n_857),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1330),
.B(n_1129),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1285),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1354),
.B(n_1203),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1381),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1260),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1355),
.B(n_1203),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1324),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1524),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1627),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1388),
.Y(n_1726)
);

BUFx12f_ASAP7_75t_L g1727 ( 
.A(n_1300),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1689),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1526),
.B(n_1203),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1689),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1279),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1410),
.B(n_857),
.Y(n_1732)
);

BUFx12f_ASAP7_75t_L g1733 ( 
.A(n_1300),
.Y(n_1733)
);

NOR2x1_ASAP7_75t_L g1734 ( 
.A(n_1410),
.B(n_861),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1279),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1526),
.B(n_1203),
.Y(n_1736)
);

INVx5_ASAP7_75t_L g1737 ( 
.A(n_1279),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1324),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1463),
.Y(n_1739)
);

OA21x2_ASAP7_75t_L g1740 ( 
.A1(n_1348),
.A2(n_866),
.B(n_861),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1287),
.A2(n_990),
.B1(n_1004),
.B2(n_966),
.Y(n_1741)
);

INVx5_ASAP7_75t_L g1742 ( 
.A(n_1279),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1487),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1325),
.B(n_1076),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1488),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1388),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1689),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1490),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1319),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1347),
.B(n_1203),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1267),
.B(n_1051),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1491),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1360),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1527),
.Y(n_1754)
);

BUFx6f_ASAP7_75t_L g1755 ( 
.A(n_1319),
.Y(n_1755)
);

CKINVDCx6p67_ASAP7_75t_R g1756 ( 
.A(n_1468),
.Y(n_1756)
);

INVx5_ASAP7_75t_L g1757 ( 
.A(n_1319),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_SL g1758 ( 
.A(n_1497),
.B(n_1076),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1358),
.B(n_1076),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1494),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1496),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1319),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1498),
.Y(n_1763)
);

INVx5_ASAP7_75t_L g1764 ( 
.A(n_1319),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1499),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1500),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1318),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1503),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1287),
.A2(n_1004),
.B1(n_1006),
.B2(n_990),
.Y(n_1769)
);

NOR2x1_ASAP7_75t_L g1770 ( 
.A(n_1345),
.B(n_866),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1267),
.B(n_1295),
.Y(n_1771)
);

BUFx12f_ASAP7_75t_L g1772 ( 
.A(n_1316),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1360),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1447),
.B(n_1203),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1504),
.Y(n_1775)
);

AND2x2_ASAP7_75t_SL g1776 ( 
.A(n_1265),
.B(n_868),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1506),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1339),
.Y(n_1778)
);

BUFx12f_ASAP7_75t_L g1779 ( 
.A(n_1316),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1372),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1295),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1339),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1339),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_L g1784 ( 
.A(n_1345),
.B(n_1508),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1368),
.Y(n_1785)
);

OAI22x1_ASAP7_75t_R g1786 ( 
.A1(n_1278),
.A2(n_1017),
.B1(n_1020),
.B2(n_1006),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1339),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1458),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1461),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1452),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1679),
.B(n_1203),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1368),
.Y(n_1792)
);

INVxp67_ASAP7_75t_L g1793 ( 
.A(n_1572),
.Y(n_1793)
);

INVx5_ASAP7_75t_L g1794 ( 
.A(n_1339),
.Y(n_1794)
);

OA21x2_ASAP7_75t_L g1795 ( 
.A1(n_1348),
.A2(n_870),
.B(n_868),
.Y(n_1795)
);

BUFx12f_ASAP7_75t_L g1796 ( 
.A(n_1343),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1509),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1255),
.A2(n_872),
.B(n_870),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1463),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1387),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1493),
.Y(n_1801)
);

BUFx12f_ASAP7_75t_L g1802 ( 
.A(n_1343),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1510),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_1406),
.Y(n_1804)
);

OAI22x1_ASAP7_75t_SL g1805 ( 
.A1(n_1278),
.A2(n_1020),
.B1(n_1023),
.B2(n_1017),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1679),
.B(n_1247),
.Y(n_1806)
);

BUFx6f_ASAP7_75t_L g1807 ( 
.A(n_1387),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1405),
.Y(n_1808)
);

INVx5_ASAP7_75t_L g1809 ( 
.A(n_1387),
.Y(n_1809)
);

BUFx8_ASAP7_75t_L g1810 ( 
.A(n_1294),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1511),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1513),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1395),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1387),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1387),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1405),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1395),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1262),
.B(n_1247),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1411),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1306),
.A2(n_907),
.B1(n_919),
.B2(n_895),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1414),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1514),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1516),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1414),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1345),
.B(n_872),
.Y(n_1825)
);

BUFx8_ASAP7_75t_L g1826 ( 
.A(n_1294),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1517),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1429),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1493),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1411),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1518),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1435),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1398),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1429),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1261),
.B(n_1263),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1264),
.Y(n_1836)
);

INVx5_ASAP7_75t_L g1837 ( 
.A(n_1398),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1565),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1398),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1435),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1436),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1436),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1565),
.Y(n_1843)
);

INVx4_ASAP7_75t_L g1844 ( 
.A(n_1398),
.Y(n_1844)
);

INVx5_ASAP7_75t_L g1845 ( 
.A(n_1398),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1406),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1266),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1633),
.B(n_956),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1406),
.B(n_961),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1473),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1406),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1404),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1268),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1379),
.B(n_874),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1271),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1272),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1473),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1445),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1473),
.Y(n_1859)
);

OAI22x1_ASAP7_75t_SL g1860 ( 
.A1(n_1291),
.A2(n_1322),
.B1(n_1327),
.B2(n_1301),
.Y(n_1860)
);

BUFx8_ASAP7_75t_SL g1861 ( 
.A(n_1291),
.Y(n_1861)
);

CKINVDCx16_ASAP7_75t_R g1862 ( 
.A(n_1507),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1540),
.B(n_1076),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1641),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1440),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1543),
.B(n_1094),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1641),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1406),
.B(n_1029),
.Y(n_1868)
);

INVx5_ASAP7_75t_L g1869 ( 
.A(n_1473),
.Y(n_1869)
);

INVx6_ASAP7_75t_L g1870 ( 
.A(n_1406),
.Y(n_1870)
);

OAI22x1_ASAP7_75t_R g1871 ( 
.A1(n_1301),
.A2(n_1039),
.B1(n_1049),
.B2(n_1023),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1445),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1274),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1473),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1478),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1277),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1492),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1478),
.Y(n_1878)
);

BUFx8_ASAP7_75t_SL g1879 ( 
.A(n_1322),
.Y(n_1879)
);

AND2x6_ASAP7_75t_L g1880 ( 
.A(n_1492),
.B(n_874),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1280),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1558),
.B(n_1566),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1505),
.Y(n_1883)
);

INVx5_ASAP7_75t_L g1884 ( 
.A(n_1478),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1505),
.Y(n_1885)
);

BUFx12f_ASAP7_75t_L g1886 ( 
.A(n_1373),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1276),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1655),
.Y(n_1888)
);

BUFx6f_ASAP7_75t_L g1889 ( 
.A(n_1478),
.Y(n_1889)
);

BUFx8_ASAP7_75t_L g1890 ( 
.A(n_1311),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1595),
.Y(n_1891)
);

AOI22x1_ASAP7_75t_SL g1892 ( 
.A1(n_1327),
.A2(n_1049),
.B1(n_1072),
.B2(n_1039),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1296),
.B(n_1246),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1281),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1385),
.B(n_876),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1655),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1386),
.B(n_1428),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1440),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1590),
.B(n_1094),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1478),
.Y(n_1900)
);

BUFx3_ASAP7_75t_L g1901 ( 
.A(n_1406),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1442),
.Y(n_1902)
);

INVx6_ASAP7_75t_L g1903 ( 
.A(n_1406),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1595),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1439),
.B(n_876),
.Y(n_1905)
);

BUFx6f_ASAP7_75t_L g1906 ( 
.A(n_1656),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1615),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1284),
.Y(n_1908)
);

CKINVDCx16_ASAP7_75t_R g1909 ( 
.A(n_1525),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_1373),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1288),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1306),
.A2(n_1073),
.B1(n_1095),
.B2(n_1072),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1290),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1656),
.Y(n_1914)
);

BUFx8_ASAP7_75t_SL g1915 ( 
.A(n_1338),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1615),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1297),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1258),
.B(n_1033),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1298),
.Y(n_1919)
);

INVx6_ASAP7_75t_L g1920 ( 
.A(n_1684),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1634),
.Y(n_1921)
);

BUFx2_ASAP7_75t_L g1922 ( 
.A(n_1442),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1448),
.Y(n_1923)
);

BUFx12f_ASAP7_75t_L g1924 ( 
.A(n_1296),
.Y(n_1924)
);

BUFx12f_ASAP7_75t_L g1925 ( 
.A(n_1448),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1675),
.B(n_1094),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1634),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1646),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1299),
.Y(n_1929)
);

BUFx8_ASAP7_75t_SL g1930 ( 
.A(n_1338),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1477),
.B(n_880),
.Y(n_1931)
);

OAI21x1_ASAP7_75t_L g1932 ( 
.A1(n_1255),
.A2(n_1292),
.B(n_1273),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1302),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_1646),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1392),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1683),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1683),
.Y(n_1937)
);

NOR2x1_ASAP7_75t_L g1938 ( 
.A(n_1569),
.B(n_880),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1303),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1674),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1674),
.Y(n_1941)
);

OA21x2_ASAP7_75t_L g1942 ( 
.A1(n_1676),
.A2(n_883),
.B(n_882),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1676),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1304),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1480),
.B(n_1094),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1495),
.B(n_1515),
.Y(n_1946)
);

BUFx12f_ASAP7_75t_L g1947 ( 
.A(n_1451),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1451),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_1677),
.Y(n_1949)
);

BUFx12f_ASAP7_75t_L g1950 ( 
.A(n_1457),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1305),
.B(n_882),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1462),
.Y(n_1952)
);

OAI21x1_ASAP7_75t_L g1953 ( 
.A1(n_1292),
.A2(n_889),
.B(n_883),
.Y(n_1953)
);

BUFx12f_ASAP7_75t_L g1954 ( 
.A(n_1457),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1307),
.B(n_889),
.Y(n_1955)
);

BUFx3_ASAP7_75t_L g1956 ( 
.A(n_1308),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1312),
.Y(n_1957)
);

AND2x6_ASAP7_75t_L g1958 ( 
.A(n_1309),
.B(n_1328),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1313),
.Y(n_1959)
);

BUFx12f_ASAP7_75t_L g1960 ( 
.A(n_1462),
.Y(n_1960)
);

OAI22x1_ASAP7_75t_SL g1961 ( 
.A1(n_1392),
.A2(n_1095),
.B1(n_1101),
.B2(n_1073),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1314),
.Y(n_1962)
);

AND2x2_ASAP7_75t_SL g1963 ( 
.A(n_1399),
.B(n_894),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1349),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1315),
.B(n_894),
.Y(n_1965)
);

BUFx12f_ASAP7_75t_L g1966 ( 
.A(n_1474),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1677),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1682),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1321),
.B(n_1326),
.Y(n_1969)
);

INVx4_ASAP7_75t_L g1970 ( 
.A(n_1328),
.Y(n_1970)
);

INVx5_ASAP7_75t_L g1971 ( 
.A(n_1570),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1682),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1286),
.B(n_1037),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1329),
.B(n_906),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1686),
.Y(n_1975)
);

INVx5_ASAP7_75t_L g1976 ( 
.A(n_1578),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1659),
.B(n_1094),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1293),
.B(n_1320),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1400),
.B(n_906),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1686),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1687),
.Y(n_1981)
);

INVx4_ASAP7_75t_L g1982 ( 
.A(n_1684),
.Y(n_1982)
);

INVx6_ASAP7_75t_L g1983 ( 
.A(n_1671),
.Y(n_1983)
);

OAI21x1_ASAP7_75t_L g1984 ( 
.A1(n_1249),
.A2(n_914),
.B(n_909),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1571),
.B(n_1114),
.Y(n_1985)
);

INVx5_ASAP7_75t_L g1986 ( 
.A(n_1311),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1323),
.B(n_1071),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1687),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1622),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1691),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1691),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1402),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1502),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1403),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1694),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1407),
.Y(n_1996)
);

AND2x4_ASAP7_75t_L g1997 ( 
.A(n_1409),
.B(n_909),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1694),
.Y(n_1998)
);

CKINVDCx16_ASAP7_75t_R g1999 ( 
.A(n_1408),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1412),
.B(n_914),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1695),
.Y(n_2001)
);

OAI21x1_ASAP7_75t_L g2002 ( 
.A1(n_1249),
.A2(n_918),
.B(n_915),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1416),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1417),
.B(n_915),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1695),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1418),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1571),
.B(n_1114),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1419),
.Y(n_2008)
);

OAI22x1_ASAP7_75t_R g2009 ( 
.A1(n_1408),
.A2(n_1134),
.B1(n_1148),
.B2(n_1101),
.Y(n_2009)
);

CKINVDCx11_ASAP7_75t_R g2010 ( 
.A(n_1413),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1251),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1420),
.B(n_918),
.Y(n_2012)
);

BUFx8_ASAP7_75t_L g2013 ( 
.A(n_1382),
.Y(n_2013)
);

BUFx8_ASAP7_75t_SL g2014 ( 
.A(n_1413),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1251),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1252),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1424),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1425),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1426),
.Y(n_2019)
);

CKINVDCx16_ASAP7_75t_R g2020 ( 
.A(n_1444),
.Y(n_2020)
);

BUFx3_ASAP7_75t_L g2021 ( 
.A(n_1427),
.Y(n_2021)
);

CKINVDCx6p67_ASAP7_75t_R g2022 ( 
.A(n_1382),
.Y(n_2022)
);

AOI22x1_ASAP7_75t_SL g2023 ( 
.A1(n_1444),
.A2(n_1148),
.B1(n_1177),
.B2(n_1134),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1431),
.Y(n_2024)
);

AND2x4_ASAP7_75t_L g2025 ( 
.A(n_1432),
.B(n_922),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1252),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_1474),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1434),
.B(n_922),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1253),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1331),
.B(n_1079),
.Y(n_2030)
);

AND2x6_ASAP7_75t_L g2031 ( 
.A(n_1437),
.B(n_924),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1580),
.B(n_1690),
.Y(n_2032)
);

INVx5_ASAP7_75t_L g2033 ( 
.A(n_1598),
.Y(n_2033)
);

BUFx12f_ASAP7_75t_L g2034 ( 
.A(n_1476),
.Y(n_2034)
);

INVx5_ASAP7_75t_L g2035 ( 
.A(n_1607),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_R g2036 ( 
.A1(n_1310),
.A2(n_779),
.B1(n_1100),
.B2(n_1093),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1573),
.Y(n_2037)
);

INVx3_ASAP7_75t_L g2038 ( 
.A(n_1349),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1253),
.Y(n_2039)
);

AND2x6_ASAP7_75t_L g2040 ( 
.A(n_1523),
.B(n_924),
.Y(n_2040)
);

BUFx8_ASAP7_75t_L g2041 ( 
.A(n_1489),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1254),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1476),
.Y(n_2043)
);

XNOR2x2_ASAP7_75t_L g2044 ( 
.A(n_1342),
.B(n_779),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1254),
.Y(n_2045)
);

BUFx3_ASAP7_75t_L g2046 ( 
.A(n_1256),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1256),
.Y(n_2047)
);

INVx5_ASAP7_75t_L g2048 ( 
.A(n_1618),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1574),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1257),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1512),
.Y(n_2051)
);

CKINVDCx20_ASAP7_75t_R g2052 ( 
.A(n_1446),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1542),
.B(n_928),
.Y(n_2053)
);

INVx4_ASAP7_75t_L g2054 ( 
.A(n_1257),
.Y(n_2054)
);

BUFx8_ASAP7_75t_L g2055 ( 
.A(n_1489),
.Y(n_2055)
);

INVxp33_ASAP7_75t_SL g2056 ( 
.A(n_1512),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1539),
.Y(n_2057)
);

INVxp67_ASAP7_75t_L g2058 ( 
.A(n_1539),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1576),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1798),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_1882),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_1882),
.Y(n_2062)
);

BUFx8_ASAP7_75t_L g2063 ( 
.A(n_1727),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1971),
.B(n_1593),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1982),
.B(n_1441),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1971),
.B(n_1593),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_1982),
.B(n_1449),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1887),
.B(n_1624),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1863),
.B(n_1283),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_L g2070 ( 
.A1(n_1932),
.A2(n_1333),
.B(n_1332),
.Y(n_2070)
);

HB1xp67_ASAP7_75t_L g2071 ( 
.A(n_1700),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1932),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1697),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1798),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1697),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1863),
.B(n_1363),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1953),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1866),
.B(n_1364),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1953),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1718),
.Y(n_2080)
);

BUFx3_ASAP7_75t_L g2081 ( 
.A(n_1718),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1906),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1790),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1701),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1701),
.Y(n_2085)
);

INVx6_ASAP7_75t_L g2086 ( 
.A(n_2033),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_1739),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1725),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1725),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1728),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1887),
.B(n_1644),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1728),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1730),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1730),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1866),
.B(n_1423),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1747),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1747),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_1848),
.B(n_1918),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_1906),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2011),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2011),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1940),
.Y(n_2102)
);

AND2x6_ASAP7_75t_L g2103 ( 
.A(n_1744),
.B(n_1661),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1899),
.B(n_1433),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1940),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2015),
.Y(n_2106)
);

INVx5_ASAP7_75t_L g2107 ( 
.A(n_1870),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1943),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1906),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2015),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1906),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1897),
.B(n_1603),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_1698),
.B(n_1603),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1899),
.B(n_1520),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2026),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1943),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2026),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_1982),
.B(n_1450),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1967),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2029),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1926),
.B(n_1579),
.Y(n_2121)
);

BUFx6f_ASAP7_75t_L g2122 ( 
.A(n_1906),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1967),
.Y(n_2123)
);

BUFx6f_ASAP7_75t_L g2124 ( 
.A(n_1914),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1968),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1968),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1790),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1975),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_2046),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1975),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_2046),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1897),
.B(n_1625),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2029),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1960),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1914),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1981),
.Y(n_2136)
);

INVx3_ASAP7_75t_L g2137 ( 
.A(n_1970),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2050),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1926),
.B(n_1583),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1897),
.B(n_1625),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_1724),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1914),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1981),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_1754),
.Y(n_2144)
);

NAND2xp33_ASAP7_75t_SL g2145 ( 
.A(n_1712),
.B(n_1548),
.Y(n_2145)
);

INVx3_ASAP7_75t_L g2146 ( 
.A(n_1970),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1990),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1744),
.B(n_1453),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2050),
.Y(n_2149)
);

XOR2xp5_ASAP7_75t_L g2150 ( 
.A(n_2044),
.B(n_1860),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1990),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1995),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1995),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1998),
.Y(n_2154)
);

NAND2x1p5_ASAP7_75t_L g2155 ( 
.A(n_1740),
.B(n_1340),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_1759),
.B(n_1584),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1753),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1753),
.Y(n_2158)
);

BUFx6f_ASAP7_75t_L g2159 ( 
.A(n_1914),
.Y(n_2159)
);

CKINVDCx16_ASAP7_75t_R g2160 ( 
.A(n_1862),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1998),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1759),
.B(n_1945),
.Y(n_2162)
);

CKINVDCx20_ASAP7_75t_R g2163 ( 
.A(n_1704),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2005),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1971),
.B(n_1630),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2005),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1942),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1973),
.B(n_1630),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1773),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1942),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_1854),
.B(n_1895),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1942),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1945),
.B(n_1585),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_1914),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1740),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1773),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_2016),
.Y(n_2177)
);

BUFx2_ASAP7_75t_L g2178 ( 
.A(n_2022),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1987),
.B(n_2030),
.Y(n_2179)
);

NOR2xp33_ASAP7_75t_L g2180 ( 
.A(n_1751),
.B(n_1549),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1729),
.B(n_1549),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1740),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1795),
.Y(n_2183)
);

OA21x2_ASAP7_75t_L g2184 ( 
.A1(n_1984),
.A2(n_1333),
.B(n_1332),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1795),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1795),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_1970),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1984),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2002),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1971),
.B(n_1548),
.Y(n_2190)
);

INVx3_ASAP7_75t_L g2191 ( 
.A(n_1696),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_1946),
.B(n_1586),
.Y(n_2192)
);

HB1xp67_ASAP7_75t_L g2193 ( 
.A(n_1989),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2002),
.Y(n_2194)
);

BUFx6f_ASAP7_75t_L g2195 ( 
.A(n_2016),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1785),
.Y(n_2196)
);

CKINVDCx6p67_ASAP7_75t_R g2197 ( 
.A(n_1727),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1785),
.Y(n_2198)
);

BUFx6f_ASAP7_75t_L g2199 ( 
.A(n_2016),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1792),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1792),
.Y(n_2201)
);

INVx2_ASAP7_75t_SL g2202 ( 
.A(n_1986),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1813),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_1854),
.B(n_1454),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1946),
.B(n_1588),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1813),
.Y(n_2206)
);

INVx6_ASAP7_75t_L g2207 ( 
.A(n_2033),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1817),
.Y(n_2208)
);

BUFx8_ASAP7_75t_L g2209 ( 
.A(n_1733),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1817),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1819),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_SL g2212 ( 
.A(n_1758),
.B(n_1564),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1819),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1830),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_1767),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1830),
.Y(n_2216)
);

CKINVDCx16_ASAP7_75t_R g2217 ( 
.A(n_1909),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1832),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1832),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1840),
.Y(n_2220)
);

BUFx6f_ASAP7_75t_L g2221 ( 
.A(n_2016),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1840),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1841),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1841),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_SL g2225 ( 
.A(n_1924),
.B(n_1726),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1978),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1729),
.B(n_1736),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1944),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1776),
.B(n_1589),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_1780),
.Y(n_2230)
);

AND2x6_ASAP7_75t_L g2231 ( 
.A(n_1977),
.B(n_928),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1842),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1842),
.Y(n_2233)
);

INVxp33_ASAP7_75t_L g2234 ( 
.A(n_1871),
.Y(n_2234)
);

BUFx8_ASAP7_75t_L g2235 ( 
.A(n_1733),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1858),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1858),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1872),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1729),
.B(n_1564),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_L g2240 ( 
.A(n_2016),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_1986),
.B(n_1577),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_2039),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_1696),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_1696),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_1788),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1872),
.Y(n_2246)
);

XOR2xp5_ASAP7_75t_L g2247 ( 
.A(n_2044),
.B(n_1446),
.Y(n_2247)
);

BUFx6f_ASAP7_75t_L g2248 ( 
.A(n_2039),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1877),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1877),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1883),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1883),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1776),
.B(n_1963),
.Y(n_2253)
);

INVxp67_ASAP7_75t_L g2254 ( 
.A(n_1816),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_2022),
.Y(n_2255)
);

NAND2x1p5_ASAP7_75t_L g2256 ( 
.A(n_1971),
.B(n_1350),
.Y(n_2256)
);

BUFx2_ASAP7_75t_L g2257 ( 
.A(n_1789),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1885),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1885),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1736),
.B(n_1577),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_1963),
.B(n_1592),
.Y(n_2261)
);

OA21x2_ASAP7_75t_L g2262 ( 
.A1(n_1891),
.A2(n_1335),
.B(n_1334),
.Y(n_2262)
);

NAND2xp33_ASAP7_75t_R g2263 ( 
.A(n_1726),
.B(n_1310),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1891),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1736),
.B(n_1791),
.Y(n_2265)
);

INVx3_ASAP7_75t_L g2266 ( 
.A(n_1723),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1904),
.Y(n_2267)
);

INVx3_ASAP7_75t_L g2268 ( 
.A(n_1723),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_1723),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_1854),
.B(n_1456),
.Y(n_2270)
);

INVxp67_ASAP7_75t_L g2271 ( 
.A(n_1816),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1904),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1907),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1944),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1907),
.Y(n_2275)
);

BUFx3_ASAP7_75t_L g2276 ( 
.A(n_1739),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_1738),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1927),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_1993),
.B(n_1250),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1927),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_1977),
.B(n_1594),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_1738),
.Y(n_2282)
);

INVx3_ASAP7_75t_L g2283 ( 
.A(n_1738),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_SL g2284 ( 
.A1(n_1741),
.A2(n_1459),
.B1(n_1530),
.B2(n_1455),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_2039),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_1824),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1928),
.Y(n_2287)
);

BUFx8_ASAP7_75t_L g2288 ( 
.A(n_1772),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1928),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1937),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1791),
.B(n_1581),
.Y(n_2291)
);

BUFx6f_ASAP7_75t_L g2292 ( 
.A(n_2039),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1937),
.Y(n_2293)
);

BUFx6f_ASAP7_75t_L g2294 ( 
.A(n_2039),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1964),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_1824),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_2042),
.Y(n_2297)
);

OAI21x1_ASAP7_75t_L g2298 ( 
.A1(n_1849),
.A2(n_1335),
.B(n_1334),
.Y(n_2298)
);

BUFx6f_ASAP7_75t_L g2299 ( 
.A(n_2042),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1964),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1964),
.Y(n_2301)
);

CKINVDCx14_ASAP7_75t_R g2302 ( 
.A(n_1756),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2038),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_2042),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_1986),
.B(n_1581),
.Y(n_2305)
);

BUFx8_ASAP7_75t_L g2306 ( 
.A(n_1772),
.Y(n_2306)
);

INVxp67_ASAP7_75t_L g2307 ( 
.A(n_1828),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2042),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_1920),
.B(n_1596),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2038),
.Y(n_2310)
);

INVxp33_ASAP7_75t_SL g2311 ( 
.A(n_1952),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1956),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2042),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_1920),
.B(n_1597),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2038),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1956),
.Y(n_2316)
);

CKINVDCx8_ASAP7_75t_R g2317 ( 
.A(n_1999),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2045),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1992),
.Y(n_2319)
);

NOR2x1_ASAP7_75t_L g2320 ( 
.A(n_1771),
.B(n_1519),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2045),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_1986),
.B(n_1591),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1791),
.B(n_1806),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_1986),
.B(n_1591),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2045),
.Y(n_2325)
);

INVx1_ASAP7_75t_SL g2326 ( 
.A(n_1828),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_SL g2327 ( 
.A(n_1924),
.B(n_1317),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_1895),
.B(n_1460),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1941),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_1920),
.B(n_1599),
.Y(n_2330)
);

HB1xp67_ASAP7_75t_L g2331 ( 
.A(n_1834),
.Y(n_2331)
);

OAI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_1985),
.A2(n_2007),
.B1(n_1920),
.B2(n_1341),
.Y(n_2332)
);

BUFx2_ASAP7_75t_L g2333 ( 
.A(n_1834),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_1898),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_2045),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2045),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1941),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1941),
.Y(n_2338)
);

XNOR2x2_ASAP7_75t_L g2339 ( 
.A(n_1769),
.B(n_1342),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1806),
.B(n_1600),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2047),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1941),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1941),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1949),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1949),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_1949),
.Y(n_2346)
);

NAND2xp33_ASAP7_75t_L g2347 ( 
.A(n_2040),
.B(n_1600),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2047),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1949),
.Y(n_2349)
);

INVx3_ASAP7_75t_L g2350 ( 
.A(n_1844),
.Y(n_2350)
);

BUFx8_ASAP7_75t_L g2351 ( 
.A(n_1779),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_1895),
.B(n_1464),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1949),
.Y(n_2353)
);

BUFx12f_ASAP7_75t_L g2354 ( 
.A(n_1810),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1972),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_1825),
.B(n_1601),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_1820),
.B(n_1898),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1972),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_2047),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2047),
.Y(n_2360)
);

OAI22xp5_ASAP7_75t_SL g2361 ( 
.A1(n_1912),
.A2(n_1459),
.B1(n_1530),
.B2(n_1455),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1972),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1806),
.B(n_1708),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_1905),
.B(n_1465),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_1825),
.B(n_1602),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_1902),
.Y(n_2366)
);

AND2x4_ASAP7_75t_L g2367 ( 
.A(n_1905),
.B(n_1466),
.Y(n_2367)
);

XNOR2x1_ASAP7_75t_L g2368 ( 
.A(n_2036),
.B(n_1401),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2047),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_1972),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_1902),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_1972),
.Y(n_2372)
);

BUFx6f_ASAP7_75t_L g2373 ( 
.A(n_1980),
.Y(n_2373)
);

INVx3_ASAP7_75t_L g2374 ( 
.A(n_1844),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_1922),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1980),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_1905),
.B(n_1469),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1980),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1980),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_1980),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1708),
.B(n_1605),
.Y(n_2381)
);

OAI22xp5_ASAP7_75t_SL g2382 ( 
.A1(n_1704),
.A2(n_1575),
.B1(n_1582),
.B2(n_1535),
.Y(n_2382)
);

BUFx6f_ASAP7_75t_L g2383 ( 
.A(n_1988),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_1988),
.Y(n_2384)
);

NAND2x1_ASAP7_75t_L g2385 ( 
.A(n_2040),
.B(n_938),
.Y(n_2385)
);

BUFx6f_ASAP7_75t_L g2386 ( 
.A(n_1988),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1708),
.B(n_1605),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1988),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_1825),
.B(n_1604),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_1893),
.B(n_1616),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_1844),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_1988),
.Y(n_2392)
);

AND2x4_ASAP7_75t_L g2393 ( 
.A(n_1931),
.B(n_1470),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_1931),
.B(n_1471),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1991),
.Y(n_2395)
);

BUFx6f_ASAP7_75t_L g2396 ( 
.A(n_1991),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_1976),
.B(n_1746),
.Y(n_2397)
);

BUFx2_ASAP7_75t_L g2398 ( 
.A(n_1922),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1991),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_1717),
.B(n_2032),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_1976),
.B(n_1616),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_1991),
.Y(n_2402)
);

OA21x2_ASAP7_75t_L g2403 ( 
.A1(n_1868),
.A2(n_1337),
.B(n_1336),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1991),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_1835),
.B(n_1606),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2001),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2001),
.Y(n_2407)
);

BUFx8_ASAP7_75t_L g2408 ( 
.A(n_1779),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2001),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2001),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2001),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1739),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_1916),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1799),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_SL g2415 ( 
.A(n_1976),
.B(n_1642),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1799),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_1916),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1916),
.Y(n_2418)
);

OAI22xp5_ASAP7_75t_L g2419 ( 
.A1(n_1712),
.A2(n_1341),
.B1(n_1353),
.B2(n_1317),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_1916),
.Y(n_2420)
);

AND2x4_ASAP7_75t_L g2421 ( 
.A(n_1931),
.B(n_1475),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_1799),
.Y(n_2422)
);

HB1xp67_ASAP7_75t_L g2423 ( 
.A(n_1705),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_1721),
.B(n_1642),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_1983),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_1916),
.Y(n_2426)
);

INVx1_ASAP7_75t_SL g2427 ( 
.A(n_1983),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_1801),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1801),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_1801),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_1921),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1829),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1829),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1829),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_1838),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_1838),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_1838),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_1835),
.B(n_2053),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1843),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1843),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1921),
.Y(n_2441)
);

BUFx2_ASAP7_75t_L g2442 ( 
.A(n_1705),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_L g2443 ( 
.A(n_1921),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_SL g2444 ( 
.A(n_1976),
.B(n_1651),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_1843),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_1921),
.Y(n_2446)
);

INVxp67_ASAP7_75t_L g2447 ( 
.A(n_2041),
.Y(n_2447)
);

BUFx6f_ASAP7_75t_L g2448 ( 
.A(n_1921),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_1864),
.Y(n_2449)
);

NAND2xp33_ASAP7_75t_SL g2450 ( 
.A(n_1721),
.B(n_1651),
.Y(n_2450)
);

INVx3_ASAP7_75t_L g2451 ( 
.A(n_2054),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_1781),
.B(n_1672),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_1934),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_1781),
.B(n_1672),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1864),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_1934),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_SL g2457 ( 
.A(n_1976),
.B(n_1746),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2054),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_2053),
.B(n_1479),
.Y(n_2459)
);

AND2x2_ASAP7_75t_L g2460 ( 
.A(n_1835),
.B(n_1608),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_1934),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_1750),
.B(n_1678),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_1934),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_1934),
.Y(n_2464)
);

AND2x2_ASAP7_75t_SL g2465 ( 
.A(n_1720),
.B(n_951),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_1720),
.Y(n_2466)
);

INVx4_ASAP7_75t_L g2467 ( 
.A(n_1870),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_1864),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_1936),
.Y(n_2469)
);

AND2x4_ASAP7_75t_L g2470 ( 
.A(n_2053),
.B(n_1482),
.Y(n_2470)
);

HB1xp67_ASAP7_75t_L g2471 ( 
.A(n_1793),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_1960),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1867),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_1936),
.Y(n_2474)
);

INVx3_ASAP7_75t_L g2475 ( 
.A(n_2054),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_1867),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_1717),
.B(n_1678),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_1936),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_1867),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2056),
.B(n_1680),
.Y(n_2480)
);

INVx3_ASAP7_75t_L g2481 ( 
.A(n_1958),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_1952),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_1969),
.B(n_1951),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_1936),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_1717),
.B(n_1680),
.Y(n_2485)
);

INVx4_ASAP7_75t_L g2486 ( 
.A(n_2467),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2462),
.B(n_1818),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2171),
.B(n_2056),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2295),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2100),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2295),
.Y(n_2491)
);

INVx2_ASAP7_75t_SL g2492 ( 
.A(n_2171),
.Y(n_2492)
);

AO21x2_ASAP7_75t_L g2493 ( 
.A1(n_2298),
.A2(n_1774),
.B(n_1710),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_2171),
.B(n_2465),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2100),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2101),
.Y(n_2496)
);

AND2x2_ASAP7_75t_L g2497 ( 
.A(n_2253),
.B(n_2043),
.Y(n_2497)
);

NAND2xp33_ASAP7_75t_L g2498 ( 
.A(n_2103),
.B(n_2043),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2226),
.B(n_1818),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2300),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2300),
.Y(n_2501)
);

OAI21xp33_ASAP7_75t_SL g2502 ( 
.A1(n_2253),
.A2(n_1938),
.B(n_1770),
.Y(n_2502)
);

INVx2_ASAP7_75t_SL g2503 ( 
.A(n_2144),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_2465),
.B(n_2058),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2301),
.Y(n_2505)
);

INVx2_ASAP7_75t_SL g2506 ( 
.A(n_2425),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2180),
.B(n_2051),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2301),
.Y(n_2508)
);

AO22x2_ASAP7_75t_L g2509 ( 
.A1(n_2368),
.A2(n_1702),
.B1(n_1709),
.B2(n_1892),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2098),
.B(n_1818),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2303),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2303),
.Y(n_2512)
);

OR2x6_ASAP7_75t_L g2513 ( 
.A(n_2354),
.B(n_1966),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2101),
.Y(n_2514)
);

INVx6_ASAP7_75t_L g2515 ( 
.A(n_2081),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2106),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_2229),
.A2(n_2031),
.B1(n_2040),
.B2(n_1353),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2310),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2310),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2106),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_2481),
.Y(n_2521)
);

INVx1_ASAP7_75t_SL g2522 ( 
.A(n_2326),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2110),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2229),
.B(n_2051),
.Y(n_2524)
);

BUFx2_ASAP7_75t_L g2525 ( 
.A(n_2257),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2424),
.B(n_2057),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2315),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2261),
.B(n_2057),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2315),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2261),
.B(n_1969),
.Y(n_2530)
);

INVxp33_ASAP7_75t_L g2531 ( 
.A(n_2193),
.Y(n_2531)
);

NAND3xp33_ASAP7_75t_L g2532 ( 
.A(n_2179),
.B(n_1722),
.C(n_1719),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2110),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2162),
.B(n_2040),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2332),
.B(n_1983),
.Y(n_2535)
);

INVx4_ASAP7_75t_L g2536 ( 
.A(n_2467),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2115),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2438),
.B(n_1969),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2452),
.B(n_2027),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2115),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2102),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2103),
.A2(n_2040),
.B1(n_2031),
.B2(n_1179),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2102),
.Y(n_2543)
);

BUFx3_ASAP7_75t_L g2544 ( 
.A(n_2081),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_2481),
.Y(n_2545)
);

AOI22xp33_ASAP7_75t_L g2546 ( 
.A1(n_2103),
.A2(n_2031),
.B1(n_2040),
.B2(n_1438),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2117),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2117),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2120),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2120),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2162),
.B(n_1707),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2133),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2133),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_2311),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2138),
.Y(n_2555)
);

BUFx6f_ASAP7_75t_L g2556 ( 
.A(n_2177),
.Y(n_2556)
);

BUFx3_ASAP7_75t_L g2557 ( 
.A(n_2080),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_2454),
.B(n_1808),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2168),
.B(n_1983),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2138),
.Y(n_2560)
);

INVxp33_ASAP7_75t_L g2561 ( 
.A(n_2071),
.Y(n_2561)
);

HB1xp67_ASAP7_75t_L g2562 ( 
.A(n_2257),
.Y(n_2562)
);

AND3x1_ASAP7_75t_L g2563 ( 
.A(n_2212),
.B(n_1865),
.C(n_1821),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2149),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2069),
.B(n_1992),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2105),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2149),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2157),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2105),
.Y(n_2569)
);

OAI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_2357),
.A2(n_2034),
.B1(n_1966),
.B2(n_1179),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2156),
.B(n_2033),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2141),
.B(n_1923),
.Y(n_2572)
);

NAND2xp33_ASAP7_75t_L g2573 ( 
.A(n_2103),
.B(n_2031),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2157),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2158),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2158),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2169),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2156),
.B(n_2231),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2169),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2108),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2231),
.B(n_2033),
.Y(n_2581)
);

AOI22xp33_ASAP7_75t_L g2582 ( 
.A1(n_2103),
.A2(n_2031),
.B1(n_1383),
.B2(n_1443),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2176),
.Y(n_2583)
);

INVx2_ASAP7_75t_SL g2584 ( 
.A(n_2427),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2176),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2231),
.B(n_2033),
.Y(n_2586)
);

INVx3_ASAP7_75t_L g2587 ( 
.A(n_2481),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2108),
.Y(n_2588)
);

AOI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2103),
.A2(n_2031),
.B1(n_1383),
.B2(n_1443),
.Y(n_2589)
);

OAI22xp5_ASAP7_75t_L g2590 ( 
.A1(n_2112),
.A2(n_2132),
.B1(n_2140),
.B2(n_2181),
.Y(n_2590)
);

OAI22xp33_ASAP7_75t_L g2591 ( 
.A1(n_2357),
.A2(n_2034),
.B1(n_1213),
.B2(n_1177),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2203),
.Y(n_2592)
);

INVxp67_ASAP7_75t_SL g2593 ( 
.A(n_2129),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2311),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2116),
.Y(n_2595)
);

INVx4_ASAP7_75t_L g2596 ( 
.A(n_2467),
.Y(n_2596)
);

INVx3_ASAP7_75t_L g2597 ( 
.A(n_2191),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2116),
.Y(n_2598)
);

BUFx6f_ASAP7_75t_L g2599 ( 
.A(n_2177),
.Y(n_2599)
);

INVx2_ASAP7_75t_SL g2600 ( 
.A(n_2309),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2203),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2208),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_SL g2603 ( 
.A(n_2241),
.B(n_1948),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2119),
.Y(n_2604)
);

INVx5_ASAP7_75t_L g2605 ( 
.A(n_2107),
.Y(n_2605)
);

BUFx2_ASAP7_75t_L g2606 ( 
.A(n_2333),
.Y(n_2606)
);

BUFx6f_ASAP7_75t_L g2607 ( 
.A(n_2177),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_2305),
.B(n_1925),
.Y(n_2608)
);

AOI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2103),
.A2(n_1484),
.B1(n_1501),
.B2(n_1438),
.Y(n_2609)
);

BUFx6f_ASAP7_75t_L g2610 ( 
.A(n_2177),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2119),
.Y(n_2611)
);

INVx2_ASAP7_75t_SL g2612 ( 
.A(n_2309),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2208),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2322),
.B(n_1925),
.Y(n_2614)
);

BUFx4f_ASAP7_75t_L g2615 ( 
.A(n_2256),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2211),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2123),
.Y(n_2617)
);

INVx4_ASAP7_75t_L g2618 ( 
.A(n_2107),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_SL g2619 ( 
.A(n_2324),
.B(n_1947),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2231),
.B(n_2035),
.Y(n_2620)
);

AND2x6_ASAP7_75t_L g2621 ( 
.A(n_2167),
.B(n_1804),
.Y(n_2621)
);

INVx2_ASAP7_75t_SL g2622 ( 
.A(n_2314),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_L g2623 ( 
.A(n_2254),
.B(n_1756),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2123),
.Y(n_2624)
);

NAND2xp33_ASAP7_75t_L g2625 ( 
.A(n_2451),
.B(n_1910),
.Y(n_2625)
);

INVx2_ASAP7_75t_SL g2626 ( 
.A(n_2314),
.Y(n_2626)
);

AOI22xp33_ASAP7_75t_L g2627 ( 
.A1(n_2231),
.A2(n_2438),
.B1(n_2270),
.B2(n_2328),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2125),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2211),
.Y(n_2629)
);

AOI21x1_ASAP7_75t_L g2630 ( 
.A1(n_2188),
.A2(n_1337),
.B(n_1336),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2213),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2125),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2126),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2213),
.Y(n_2634)
);

NAND2xp33_ASAP7_75t_L g2635 ( 
.A(n_2451),
.B(n_1910),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2214),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_2271),
.B(n_2307),
.Y(n_2637)
);

AND3x1_ASAP7_75t_L g2638 ( 
.A(n_2113),
.B(n_2036),
.C(n_954),
.Y(n_2638)
);

INVx4_ASAP7_75t_L g2639 ( 
.A(n_2107),
.Y(n_2639)
);

INVxp67_ASAP7_75t_L g2640 ( 
.A(n_2333),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_2390),
.B(n_1947),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2214),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2126),
.Y(n_2643)
);

AOI22xp33_ASAP7_75t_L g2644 ( 
.A1(n_2231),
.A2(n_1501),
.B1(n_1484),
.B2(n_1951),
.Y(n_2644)
);

INVx2_ASAP7_75t_SL g2645 ( 
.A(n_2330),
.Y(n_2645)
);

AND2x6_ASAP7_75t_L g2646 ( 
.A(n_2167),
.B(n_1804),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2442),
.B(n_2148),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2069),
.B(n_2017),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2128),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_2134),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2442),
.B(n_1950),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2218),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_L g2653 ( 
.A(n_2371),
.B(n_1950),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2128),
.Y(n_2654)
);

OAI22x1_ASAP7_75t_L g2655 ( 
.A1(n_2247),
.A2(n_1786),
.B1(n_2009),
.B2(n_1415),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2218),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2471),
.B(n_1954),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2231),
.B(n_2035),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2219),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2219),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2130),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_2177),
.Y(n_2662)
);

INVx4_ASAP7_75t_L g2663 ( 
.A(n_2107),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2130),
.Y(n_2664)
);

AND2x4_ASAP7_75t_L g2665 ( 
.A(n_2483),
.B(n_2017),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2136),
.Y(n_2666)
);

NAND2xp33_ASAP7_75t_L g2667 ( 
.A(n_2451),
.B(n_1958),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2121),
.B(n_2035),
.Y(n_2668)
);

INVx3_ASAP7_75t_L g2669 ( 
.A(n_2191),
.Y(n_2669)
);

OR2x2_ASAP7_75t_L g2670 ( 
.A(n_2279),
.B(n_2020),
.Y(n_2670)
);

INVxp33_ASAP7_75t_L g2671 ( 
.A(n_2382),
.Y(n_2671)
);

INVxp67_ASAP7_75t_SL g2672 ( 
.A(n_2129),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2222),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2148),
.B(n_1954),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2222),
.Y(n_2675)
);

AOI21x1_ASAP7_75t_L g2676 ( 
.A1(n_2188),
.A2(n_1346),
.B(n_1344),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2423),
.B(n_1681),
.Y(n_2677)
);

INVx2_ASAP7_75t_SL g2678 ( 
.A(n_2330),
.Y(n_2678)
);

AO21x2_ASAP7_75t_L g2679 ( 
.A1(n_2298),
.A2(n_1847),
.B(n_1836),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2136),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2076),
.B(n_2021),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2223),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2148),
.B(n_1681),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2223),
.Y(n_2684)
);

INVx4_ASAP7_75t_L g2685 ( 
.A(n_2107),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2143),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2076),
.B(n_2078),
.Y(n_2687)
);

AO22x2_ASAP7_75t_L g2688 ( 
.A1(n_2368),
.A2(n_1709),
.B1(n_1702),
.B2(n_1892),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_2239),
.B(n_1685),
.Y(n_2689)
);

BUFx10_ASAP7_75t_L g2690 ( 
.A(n_2065),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2224),
.Y(n_2691)
);

BUFx10_ASAP7_75t_L g2692 ( 
.A(n_2065),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_L g2693 ( 
.A(n_2466),
.B(n_2419),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2224),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2225),
.B(n_1685),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2143),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2121),
.B(n_2035),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2147),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2232),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2147),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2151),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2151),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2232),
.Y(n_2703)
);

OAI22xp5_ASAP7_75t_L g2704 ( 
.A1(n_2260),
.A2(n_904),
.B1(n_1289),
.B2(n_1269),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2139),
.B(n_2035),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2191),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2152),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2078),
.B(n_2021),
.Y(n_2708)
);

NAND2xp33_ASAP7_75t_L g2709 ( 
.A(n_2458),
.B(n_1958),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2152),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2153),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2153),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2237),
.Y(n_2713)
);

AOI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2173),
.A2(n_1213),
.B1(n_1880),
.B2(n_1958),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2154),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2237),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_SL g2717 ( 
.A(n_2065),
.B(n_1951),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2154),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2139),
.B(n_2048),
.Y(n_2719)
);

BUFx10_ASAP7_75t_L g2720 ( 
.A(n_2067),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2258),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2161),
.Y(n_2722)
);

NOR2xp33_ASAP7_75t_L g2723 ( 
.A(n_2480),
.B(n_1351),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2161),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2258),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2164),
.Y(n_2726)
);

AOI22xp33_ASAP7_75t_L g2727 ( 
.A1(n_2204),
.A2(n_1965),
.B1(n_1974),
.B2(n_1955),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2164),
.Y(n_2728)
);

NOR2xp33_ASAP7_75t_L g2729 ( 
.A(n_2061),
.B(n_1421),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2095),
.B(n_1955),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2173),
.B(n_2281),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2166),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2267),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2166),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2085),
.Y(n_2735)
);

AOI21x1_ASAP7_75t_L g2736 ( 
.A1(n_2189),
.A2(n_1346),
.B(n_1344),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2267),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2272),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2134),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2095),
.B(n_1955),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2085),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2088),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2272),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_SL g2744 ( 
.A(n_2067),
.B(n_1965),
.Y(n_2744)
);

BUFx10_ASAP7_75t_L g2745 ( 
.A(n_2067),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2281),
.B(n_2048),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2472),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2118),
.B(n_2320),
.Y(n_2748)
);

INVx2_ASAP7_75t_SL g2749 ( 
.A(n_2087),
.Y(n_2749)
);

AOI22xp33_ASAP7_75t_L g2750 ( 
.A1(n_2204),
.A2(n_1974),
.B1(n_1979),
.B2(n_1965),
.Y(n_2750)
);

AND2x6_ASAP7_75t_L g2751 ( 
.A(n_2170),
.B(n_1846),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2088),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2192),
.B(n_2048),
.Y(n_2753)
);

NOR2xp33_ASAP7_75t_R g2754 ( 
.A(n_2302),
.B(n_2472),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2090),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_SL g2756 ( 
.A(n_2118),
.B(n_2104),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2192),
.B(n_2048),
.Y(n_2757)
);

INVx5_ASAP7_75t_L g2758 ( 
.A(n_2107),
.Y(n_2758)
);

INVx2_ASAP7_75t_SL g2759 ( 
.A(n_2087),
.Y(n_2759)
);

BUFx3_ASAP7_75t_L g2760 ( 
.A(n_2080),
.Y(n_2760)
);

INVx2_ASAP7_75t_SL g2761 ( 
.A(n_2276),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_SL g2762 ( 
.A(n_2118),
.B(n_1974),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2205),
.B(n_2048),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2243),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2104),
.B(n_1979),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2090),
.Y(n_2766)
);

INVx3_ASAP7_75t_L g2767 ( 
.A(n_2243),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2092),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2273),
.Y(n_2769)
);

INVxp33_ASAP7_75t_L g2770 ( 
.A(n_2215),
.Y(n_2770)
);

OR2x6_ASAP7_75t_L g2771 ( 
.A(n_2354),
.B(n_1796),
.Y(n_2771)
);

AOI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2114),
.A2(n_1880),
.B1(n_1958),
.B2(n_1979),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_2114),
.B(n_1997),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2205),
.B(n_1997),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2356),
.B(n_1997),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2273),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2280),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2280),
.Y(n_2778)
);

INVx1_ASAP7_75t_SL g2779 ( 
.A(n_2375),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2092),
.Y(n_2780)
);

INVx3_ASAP7_75t_L g2781 ( 
.A(n_2243),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2483),
.B(n_2000),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2287),
.Y(n_2783)
);

BUFx6f_ASAP7_75t_L g2784 ( 
.A(n_2195),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2458),
.B(n_2024),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2093),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2093),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2096),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2287),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2096),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2196),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2356),
.B(n_2365),
.Y(n_2792)
);

INVx3_ASAP7_75t_L g2793 ( 
.A(n_2244),
.Y(n_2793)
);

NAND3xp33_ASAP7_75t_L g2794 ( 
.A(n_2347),
.B(n_1732),
.C(n_1716),
.Y(n_2794)
);

NOR2x1p5_ASAP7_75t_L g2795 ( 
.A(n_2197),
.B(n_1796),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_SL g2796 ( 
.A(n_2291),
.B(n_2000),
.Y(n_2796)
);

BUFx2_ASAP7_75t_L g2797 ( 
.A(n_2375),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_L g2798 ( 
.A(n_2062),
.B(n_1430),
.Y(n_2798)
);

INVx3_ASAP7_75t_L g2799 ( 
.A(n_2244),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2340),
.B(n_2000),
.Y(n_2800)
);

AOI22xp33_ASAP7_75t_L g2801 ( 
.A1(n_2204),
.A2(n_2012),
.B1(n_2025),
.B2(n_2004),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2293),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2196),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2365),
.B(n_2004),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2198),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2458),
.B(n_1853),
.Y(n_2806)
);

BUFx6f_ASAP7_75t_L g2807 ( 
.A(n_2195),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2475),
.B(n_1855),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2198),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2200),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2293),
.Y(n_2811)
);

INVxp67_ASAP7_75t_SL g2812 ( 
.A(n_2129),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_SL g2813 ( 
.A(n_2270),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2475),
.B(n_2137),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2073),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2200),
.Y(n_2816)
);

INVxp67_ASAP7_75t_SL g2817 ( 
.A(n_2131),
.Y(n_2817)
);

INVx3_ASAP7_75t_L g2818 ( 
.A(n_2244),
.Y(n_2818)
);

OR2x6_ASAP7_75t_L g2819 ( 
.A(n_2178),
.B(n_2255),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2201),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2073),
.Y(n_2821)
);

INVx8_ASAP7_75t_L g2822 ( 
.A(n_2475),
.Y(n_2822)
);

OAI22xp33_ASAP7_75t_L g2823 ( 
.A1(n_2263),
.A2(n_1481),
.B1(n_1467),
.B2(n_804),
.Y(n_2823)
);

AOI21x1_ASAP7_75t_L g2824 ( 
.A1(n_2189),
.A2(n_1784),
.B(n_1856),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2075),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2075),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2381),
.B(n_2004),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_2387),
.B(n_1802),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2201),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2084),
.Y(n_2830)
);

OR2x6_ASAP7_75t_L g2831 ( 
.A(n_2178),
.B(n_1802),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2206),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2206),
.Y(n_2833)
);

INVx2_ASAP7_75t_SL g2834 ( 
.A(n_2276),
.Y(n_2834)
);

NOR2xp33_ASAP7_75t_L g2835 ( 
.A(n_2477),
.B(n_1886),
.Y(n_2835)
);

AOI22xp5_ASAP7_75t_L g2836 ( 
.A1(n_2389),
.A2(n_1880),
.B1(n_1958),
.B2(n_2012),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2084),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2089),
.Y(n_2838)
);

AND2x4_ASAP7_75t_L g2839 ( 
.A(n_2389),
.B(n_2405),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2210),
.Y(n_2840)
);

INVxp67_ASAP7_75t_SL g2841 ( 
.A(n_2131),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2089),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2210),
.Y(n_2843)
);

BUFx4f_ASAP7_75t_L g2844 ( 
.A(n_2256),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2094),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2137),
.B(n_2019),
.Y(n_2846)
);

NAND3xp33_ASAP7_75t_L g2847 ( 
.A(n_2137),
.B(n_1734),
.C(n_1873),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2146),
.B(n_1876),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2094),
.Y(n_2849)
);

AND3x1_ASAP7_75t_L g2850 ( 
.A(n_2327),
.B(n_954),
.C(n_951),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2097),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2266),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2216),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2216),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2220),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2220),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2485),
.B(n_2012),
.Y(n_2857)
);

AND3x2_ASAP7_75t_L g2858 ( 
.A(n_2255),
.B(n_1852),
.C(n_1861),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2097),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2262),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2233),
.Y(n_2861)
);

INVx8_ASAP7_75t_L g2862 ( 
.A(n_2146),
.Y(n_2862)
);

INVx4_ASAP7_75t_L g2863 ( 
.A(n_2131),
.Y(n_2863)
);

INVx5_ASAP7_75t_L g2864 ( 
.A(n_2195),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2233),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2146),
.B(n_2187),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2187),
.B(n_1881),
.Y(n_2867)
);

BUFx4f_ASAP7_75t_L g2868 ( 
.A(n_2256),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2236),
.Y(n_2869)
);

AOI22xp33_ASAP7_75t_L g2870 ( 
.A1(n_2270),
.A2(n_2028),
.B1(n_2025),
.B2(n_1908),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2236),
.Y(n_2871)
);

OAI22xp33_ASAP7_75t_L g2872 ( 
.A1(n_2398),
.A2(n_804),
.B1(n_816),
.B2(n_751),
.Y(n_2872)
);

BUFx6f_ASAP7_75t_L g2873 ( 
.A(n_2195),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2262),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2262),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2262),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2238),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2238),
.Y(n_2878)
);

NOR2xp33_ASAP7_75t_L g2879 ( 
.A(n_2286),
.B(n_1886),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2246),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2187),
.B(n_2008),
.Y(n_2881)
);

BUFx3_ASAP7_75t_L g2882 ( 
.A(n_2080),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2246),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2091),
.B(n_2018),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2249),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2249),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2250),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2250),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2251),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2398),
.B(n_2025),
.Y(n_2890)
);

AND2x2_ASAP7_75t_SL g2891 ( 
.A(n_2170),
.B(n_967),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2296),
.B(n_1810),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2251),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2252),
.Y(n_2894)
);

NOR2xp33_ASAP7_75t_L g2895 ( 
.A(n_2331),
.B(n_1810),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_2063),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2400),
.B(n_1894),
.Y(n_2897)
);

INVx1_ASAP7_75t_SL g2898 ( 
.A(n_2163),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2252),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2334),
.B(n_2366),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2259),
.Y(n_2901)
);

BUFx2_ASAP7_75t_L g2902 ( 
.A(n_2230),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2259),
.Y(n_2903)
);

CKINVDCx6p67_ASAP7_75t_R g2904 ( 
.A(n_2197),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2405),
.B(n_1911),
.Y(n_2905)
);

OR2x6_ASAP7_75t_L g2906 ( 
.A(n_2447),
.B(n_2028),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2245),
.B(n_1826),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_SL g2908 ( 
.A(n_2328),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2264),
.Y(n_2909)
);

BUFx3_ASAP7_75t_L g2910 ( 
.A(n_2063),
.Y(n_2910)
);

INVx2_ASAP7_75t_SL g2911 ( 
.A(n_2155),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2264),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_L g2913 ( 
.A1(n_2328),
.A2(n_2028),
.B1(n_1917),
.B2(n_1919),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2275),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2275),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2278),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2278),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2145),
.B(n_2037),
.Y(n_2918)
);

BUFx3_ASAP7_75t_L g2919 ( 
.A(n_2086),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2460),
.B(n_1913),
.Y(n_2920)
);

HB1xp67_ASAP7_75t_L g2921 ( 
.A(n_2160),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2289),
.Y(n_2922)
);

BUFx2_ASAP7_75t_L g2923 ( 
.A(n_2217),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2289),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2290),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2290),
.Y(n_2926)
);

AOI22xp33_ASAP7_75t_L g2927 ( 
.A1(n_2352),
.A2(n_1933),
.B1(n_1939),
.B2(n_1929),
.Y(n_2927)
);

NOR2xp33_ASAP7_75t_L g2928 ( 
.A(n_2507),
.B(n_2482),
.Y(n_2928)
);

NOR2xp33_ASAP7_75t_L g2929 ( 
.A(n_2535),
.B(n_2524),
.Y(n_2929)
);

INVx2_ASAP7_75t_SL g2930 ( 
.A(n_2690),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2815),
.Y(n_2931)
);

OR2x2_ASAP7_75t_L g2932 ( 
.A(n_2522),
.B(n_2279),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2524),
.B(n_2528),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2815),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2510),
.B(n_2460),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2821),
.Y(n_2936)
);

INVx3_ASAP7_75t_L g2937 ( 
.A(n_2486),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2821),
.Y(n_2938)
);

INVxp67_ASAP7_75t_L g2939 ( 
.A(n_2525),
.Y(n_2939)
);

AND2x6_ASAP7_75t_L g2940 ( 
.A(n_2542),
.B(n_2172),
.Y(n_2940)
);

BUFx6f_ASAP7_75t_L g2941 ( 
.A(n_2556),
.Y(n_2941)
);

AOI22xp33_ASAP7_75t_L g2942 ( 
.A1(n_2891),
.A2(n_2339),
.B1(n_2361),
.B2(n_2284),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2600),
.B(n_2352),
.Y(n_2943)
);

AND2x6_ASAP7_75t_L g2944 ( 
.A(n_2542),
.B(n_2172),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2600),
.B(n_2352),
.Y(n_2945)
);

NAND2xp33_ASAP7_75t_L g2946 ( 
.A(n_2822),
.B(n_2862),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_L g2947 ( 
.A(n_2528),
.B(n_2165),
.Y(n_2947)
);

INVx4_ASAP7_75t_SL g2948 ( 
.A(n_2621),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2489),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2489),
.Y(n_2950)
);

AND2x6_ASAP7_75t_L g2951 ( 
.A(n_2860),
.B(n_2175),
.Y(n_2951)
);

AO22x2_ASAP7_75t_L g2952 ( 
.A1(n_2494),
.A2(n_2150),
.B1(n_2247),
.B2(n_2023),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2525),
.B(n_2364),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2687),
.B(n_2364),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2491),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_2690),
.B(n_2195),
.Y(n_2956)
);

AND2x6_ASAP7_75t_L g2957 ( 
.A(n_2860),
.B(n_2175),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2590),
.B(n_2064),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_2690),
.B(n_2199),
.Y(n_2959)
);

INVx3_ASAP7_75t_L g2960 ( 
.A(n_2486),
.Y(n_2960)
);

AND2x6_ASAP7_75t_L g2961 ( 
.A(n_2874),
.B(n_2182),
.Y(n_2961)
);

INVx3_ASAP7_75t_L g2962 ( 
.A(n_2486),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2491),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_L g2964 ( 
.A(n_2556),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2825),
.Y(n_2965)
);

BUFx6f_ASAP7_75t_L g2966 ( 
.A(n_2556),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2500),
.Y(n_2967)
);

BUFx3_ASAP7_75t_L g2968 ( 
.A(n_2923),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2612),
.B(n_2364),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2500),
.Y(n_2970)
);

BUFx6f_ASAP7_75t_L g2971 ( 
.A(n_2556),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2612),
.B(n_2367),
.Y(n_2972)
);

BUFx3_ASAP7_75t_L g2973 ( 
.A(n_2923),
.Y(n_2973)
);

BUFx3_ASAP7_75t_L g2974 ( 
.A(n_2896),
.Y(n_2974)
);

BUFx3_ASAP7_75t_L g2975 ( 
.A(n_2896),
.Y(n_2975)
);

BUFx6f_ASAP7_75t_L g2976 ( 
.A(n_2556),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2501),
.Y(n_2977)
);

AO22x2_ASAP7_75t_L g2978 ( 
.A1(n_2638),
.A2(n_2150),
.B1(n_2023),
.B2(n_2339),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2486),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2622),
.B(n_2367),
.Y(n_2980)
);

INVx3_ASAP7_75t_L g2981 ( 
.A(n_2536),
.Y(n_2981)
);

AND2x4_ASAP7_75t_L g2982 ( 
.A(n_2492),
.B(n_2228),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2501),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2825),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2622),
.B(n_2367),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_2690),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2505),
.Y(n_2987)
);

BUFx6f_ASAP7_75t_L g2988 ( 
.A(n_2599),
.Y(n_2988)
);

OR2x2_ASAP7_75t_L g2989 ( 
.A(n_2670),
.B(n_2377),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2505),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2626),
.B(n_2377),
.Y(n_2991)
);

AND2x4_ASAP7_75t_L g2992 ( 
.A(n_2492),
.B(n_2274),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2692),
.B(n_2199),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2626),
.B(n_2377),
.Y(n_2994)
);

OR2x6_ASAP7_75t_L g2995 ( 
.A(n_2911),
.B(n_2385),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2508),
.Y(n_2996)
);

INVxp33_ASAP7_75t_L g2997 ( 
.A(n_2562),
.Y(n_2997)
);

INVx4_ASAP7_75t_SL g2998 ( 
.A(n_2621),
.Y(n_2998)
);

INVx5_ASAP7_75t_L g2999 ( 
.A(n_2621),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2504),
.B(n_2497),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2497),
.B(n_2066),
.Y(n_3001)
);

AND2x4_ASAP7_75t_L g3002 ( 
.A(n_2839),
.B(n_2782),
.Y(n_3002)
);

BUFx6f_ASAP7_75t_L g3003 ( 
.A(n_2599),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2508),
.Y(n_3004)
);

BUFx2_ASAP7_75t_L g3005 ( 
.A(n_2606),
.Y(n_3005)
);

AND2x4_ASAP7_75t_L g3006 ( 
.A(n_2839),
.B(n_2312),
.Y(n_3006)
);

INVx3_ASAP7_75t_L g3007 ( 
.A(n_2536),
.Y(n_3007)
);

INVx5_ASAP7_75t_L g3008 ( 
.A(n_2621),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2511),
.Y(n_3009)
);

BUFx6f_ASAP7_75t_L g3010 ( 
.A(n_2599),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2645),
.B(n_2393),
.Y(n_3011)
);

BUFx3_ASAP7_75t_L g3012 ( 
.A(n_2910),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2511),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2756),
.B(n_2316),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2512),
.Y(n_3015)
);

INVx5_ASAP7_75t_L g3016 ( 
.A(n_2621),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2826),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2645),
.B(n_2393),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2826),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2512),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2830),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2830),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2837),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2837),
.Y(n_3024)
);

INVx4_ASAP7_75t_L g3025 ( 
.A(n_2862),
.Y(n_3025)
);

BUFx2_ASAP7_75t_L g3026 ( 
.A(n_2606),
.Y(n_3026)
);

INVx1_ASAP7_75t_SL g3027 ( 
.A(n_2779),
.Y(n_3027)
);

OAI22xp33_ASAP7_75t_L g3028 ( 
.A1(n_2693),
.A2(n_2127),
.B1(n_2083),
.B2(n_2317),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2518),
.Y(n_3029)
);

INVx4_ASAP7_75t_L g3030 ( 
.A(n_2862),
.Y(n_3030)
);

AND2x4_ASAP7_75t_L g3031 ( 
.A(n_2839),
.B(n_2319),
.Y(n_3031)
);

BUFx6f_ASAP7_75t_L g3032 ( 
.A(n_2599),
.Y(n_3032)
);

BUFx2_ASAP7_75t_L g3033 ( 
.A(n_2797),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2687),
.B(n_2393),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2678),
.B(n_2394),
.Y(n_3035)
);

INVx3_ASAP7_75t_L g3036 ( 
.A(n_2536),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2838),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2678),
.B(n_2530),
.Y(n_3038)
);

BUFx6f_ASAP7_75t_L g3039 ( 
.A(n_2599),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2530),
.B(n_2394),
.Y(n_3040)
);

BUFx3_ASAP7_75t_L g3041 ( 
.A(n_2910),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2518),
.Y(n_3042)
);

AND2x2_ASAP7_75t_L g3043 ( 
.A(n_2792),
.B(n_2394),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_SL g3044 ( 
.A(n_2692),
.B(n_2199),
.Y(n_3044)
);

AND2x2_ASAP7_75t_SL g3045 ( 
.A(n_2891),
.B(n_2227),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2519),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2838),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_2559),
.B(n_2397),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_2754),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2842),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2519),
.Y(n_3051)
);

BUFx2_ASAP7_75t_L g3052 ( 
.A(n_2797),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2792),
.B(n_2421),
.Y(n_3053)
);

HB1xp67_ASAP7_75t_L g3054 ( 
.A(n_2902),
.Y(n_3054)
);

INVx1_ASAP7_75t_SL g3055 ( 
.A(n_2902),
.Y(n_3055)
);

AND2x4_ASAP7_75t_L g3056 ( 
.A(n_2839),
.B(n_2421),
.Y(n_3056)
);

INVx3_ASAP7_75t_L g3057 ( 
.A(n_2536),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2527),
.Y(n_3058)
);

INVx3_ASAP7_75t_L g3059 ( 
.A(n_2596),
.Y(n_3059)
);

BUFx2_ASAP7_75t_L g3060 ( 
.A(n_2921),
.Y(n_3060)
);

BUFx3_ASAP7_75t_L g3061 ( 
.A(n_2515),
.Y(n_3061)
);

INVx4_ASAP7_75t_SL g3062 ( 
.A(n_2621),
.Y(n_3062)
);

INVx4_ASAP7_75t_L g3063 ( 
.A(n_2862),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2731),
.B(n_2421),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2730),
.B(n_2459),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2842),
.Y(n_3066)
);

NAND2x1p5_ASAP7_75t_L g3067 ( 
.A(n_2615),
.B(n_2385),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2527),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2529),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2529),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2735),
.Y(n_3071)
);

AND2x4_ASAP7_75t_SL g3072 ( 
.A(n_2692),
.B(n_2459),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2735),
.Y(n_3073)
);

BUFx6f_ASAP7_75t_L g3074 ( 
.A(n_2607),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2845),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2774),
.B(n_2459),
.Y(n_3076)
);

INVx5_ASAP7_75t_L g3077 ( 
.A(n_2621),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2741),
.Y(n_3078)
);

INVx3_ASAP7_75t_L g3079 ( 
.A(n_2596),
.Y(n_3079)
);

OR2x2_ASAP7_75t_L g3080 ( 
.A(n_2670),
.B(n_2083),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2741),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2742),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2742),
.Y(n_3083)
);

BUFx6f_ASAP7_75t_L g3084 ( 
.A(n_2607),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2845),
.Y(n_3085)
);

BUFx6f_ASAP7_75t_L g3086 ( 
.A(n_2607),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_2730),
.B(n_2470),
.Y(n_3087)
);

AND2x4_ASAP7_75t_L g3088 ( 
.A(n_2782),
.B(n_2538),
.Y(n_3088)
);

BUFx10_ASAP7_75t_L g3089 ( 
.A(n_2623),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2752),
.Y(n_3090)
);

INVx6_ASAP7_75t_L g3091 ( 
.A(n_2692),
.Y(n_3091)
);

AND2x4_ASAP7_75t_L g3092 ( 
.A(n_2782),
.B(n_2470),
.Y(n_3092)
);

BUFx2_ASAP7_75t_L g3093 ( 
.A(n_2640),
.Y(n_3093)
);

INVx3_ASAP7_75t_L g3094 ( 
.A(n_2596),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2849),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2607),
.Y(n_3096)
);

INVx3_ASAP7_75t_L g3097 ( 
.A(n_2596),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2752),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2488),
.B(n_2748),
.Y(n_3099)
);

BUFx6f_ASAP7_75t_L g3100 ( 
.A(n_2607),
.Y(n_3100)
);

INVx4_ASAP7_75t_L g3101 ( 
.A(n_2862),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2526),
.B(n_2457),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_SL g3103 ( 
.A(n_2720),
.B(n_2199),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2849),
.Y(n_3104)
);

BUFx2_ASAP7_75t_L g3105 ( 
.A(n_2898),
.Y(n_3105)
);

OR2x6_ASAP7_75t_L g3106 ( 
.A(n_2911),
.B(n_2513),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2851),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2755),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2774),
.B(n_2470),
.Y(n_3109)
);

AND2x4_ASAP7_75t_L g3110 ( 
.A(n_2782),
.B(n_2202),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_2538),
.B(n_2202),
.Y(n_3111)
);

INVx2_ASAP7_75t_SL g3112 ( 
.A(n_2720),
.Y(n_3112)
);

CKINVDCx5p33_ASAP7_75t_R g3113 ( 
.A(n_2554),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2851),
.Y(n_3114)
);

NOR2x1p5_ASAP7_75t_L g3115 ( 
.A(n_2904),
.B(n_2127),
.Y(n_3115)
);

AND2x4_ASAP7_75t_L g3116 ( 
.A(n_2538),
.B(n_2266),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2755),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2884),
.B(n_2265),
.Y(n_3118)
);

INVx4_ASAP7_75t_L g3119 ( 
.A(n_2822),
.Y(n_3119)
);

INVx5_ASAP7_75t_L g3120 ( 
.A(n_2646),
.Y(n_3120)
);

BUFx2_ASAP7_75t_L g3121 ( 
.A(n_2503),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_SL g3122 ( 
.A(n_2720),
.B(n_2199),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2720),
.B(n_2221),
.Y(n_3123)
);

CKINVDCx11_ASAP7_75t_R g3124 ( 
.A(n_2904),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_SL g3125 ( 
.A(n_2745),
.B(n_2615),
.Y(n_3125)
);

AND2x2_ASAP7_75t_SL g3126 ( 
.A(n_2891),
.B(n_2323),
.Y(n_3126)
);

AND2x4_ASAP7_75t_L g3127 ( 
.A(n_2538),
.B(n_2266),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_2859),
.Y(n_3128)
);

BUFx3_ASAP7_75t_L g3129 ( 
.A(n_2515),
.Y(n_3129)
);

INVx4_ASAP7_75t_L g3130 ( 
.A(n_2822),
.Y(n_3130)
);

BUFx3_ASAP7_75t_L g3131 ( 
.A(n_2515),
.Y(n_3131)
);

NAND2xp33_ASAP7_75t_SL g3132 ( 
.A(n_2554),
.B(n_2190),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_2502),
.B(n_2401),
.Y(n_3133)
);

BUFx6f_ASAP7_75t_L g3134 ( 
.A(n_2610),
.Y(n_3134)
);

INVx4_ASAP7_75t_L g3135 ( 
.A(n_2822),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2859),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2766),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_2822),
.Y(n_3138)
);

OAI22xp5_ASAP7_75t_L g3139 ( 
.A1(n_2627),
.A2(n_2269),
.B1(n_2277),
.B2(n_2268),
.Y(n_3139)
);

INVx1_ASAP7_75t_SL g3140 ( 
.A(n_2503),
.Y(n_3140)
);

BUFx2_ASAP7_75t_L g3141 ( 
.A(n_2819),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2568),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2775),
.B(n_2363),
.Y(n_3143)
);

BUFx6f_ASAP7_75t_L g3144 ( 
.A(n_2610),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2740),
.B(n_2317),
.Y(n_3145)
);

BUFx3_ASAP7_75t_L g3146 ( 
.A(n_2515),
.Y(n_3146)
);

INVx3_ASAP7_75t_L g3147 ( 
.A(n_2863),
.Y(n_3147)
);

OAI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_2578),
.A2(n_2609),
.B1(n_2589),
.B2(n_2582),
.Y(n_3148)
);

OAI22xp5_ASAP7_75t_L g3149 ( 
.A1(n_2546),
.A2(n_2269),
.B1(n_2277),
.B2(n_2268),
.Y(n_3149)
);

NOR2xp33_ASAP7_75t_L g3150 ( 
.A(n_2502),
.B(n_2415),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2568),
.Y(n_3151)
);

BUFx3_ASAP7_75t_L g3152 ( 
.A(n_2544),
.Y(n_3152)
);

INVx2_ASAP7_75t_SL g3153 ( 
.A(n_2745),
.Y(n_3153)
);

AOI22xp5_ASAP7_75t_L g3154 ( 
.A1(n_2745),
.A2(n_2450),
.B1(n_2444),
.B2(n_2269),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2766),
.Y(n_3155)
);

AOI22xp5_ASAP7_75t_L g3156 ( 
.A1(n_2745),
.A2(n_2277),
.B1(n_2282),
.B2(n_2268),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2768),
.Y(n_3157)
);

HB1xp67_ASAP7_75t_L g3158 ( 
.A(n_2813),
.Y(n_3158)
);

OAI22xp5_ASAP7_75t_L g3159 ( 
.A1(n_2644),
.A2(n_2283),
.B1(n_2282),
.B2(n_2350),
.Y(n_3159)
);

CKINVDCx5p33_ASAP7_75t_R g3160 ( 
.A(n_2594),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2768),
.Y(n_3161)
);

AO21x2_ASAP7_75t_L g3162 ( 
.A1(n_2679),
.A2(n_2183),
.B(n_2182),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2775),
.B(n_2282),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2780),
.Y(n_3164)
);

INVx3_ASAP7_75t_L g3165 ( 
.A(n_2863),
.Y(n_3165)
);

NAND2x1p5_ASAP7_75t_L g3166 ( 
.A(n_2615),
.B(n_2283),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2740),
.B(n_1535),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2780),
.Y(n_3168)
);

INVx4_ASAP7_75t_L g3169 ( 
.A(n_2844),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_2665),
.B(n_2283),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2786),
.Y(n_3171)
);

INVx1_ASAP7_75t_SL g3172 ( 
.A(n_2770),
.Y(n_3172)
);

AND2x6_ASAP7_75t_L g3173 ( 
.A(n_2874),
.B(n_2183),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2786),
.Y(n_3174)
);

BUFx6f_ASAP7_75t_L g3175 ( 
.A(n_2610),
.Y(n_3175)
);

INVx1_ASAP7_75t_SL g3176 ( 
.A(n_2531),
.Y(n_3176)
);

NOR2xp33_ASAP7_75t_L g3177 ( 
.A(n_2539),
.B(n_2350),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2787),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2574),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_2665),
.B(n_1957),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2574),
.Y(n_3181)
);

BUFx3_ASAP7_75t_L g3182 ( 
.A(n_2544),
.Y(n_3182)
);

INVx5_ASAP7_75t_L g3183 ( 
.A(n_2646),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2575),
.Y(n_3184)
);

AND2x4_ASAP7_75t_L g3185 ( 
.A(n_2665),
.B(n_1959),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_2729),
.B(n_1575),
.Y(n_3186)
);

INVx4_ASAP7_75t_L g3187 ( 
.A(n_2844),
.Y(n_3187)
);

AND2x6_ASAP7_75t_L g3188 ( 
.A(n_2875),
.B(n_2185),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2787),
.Y(n_3189)
);

NAND2x1p5_ASAP7_75t_L g3190 ( 
.A(n_2844),
.B(n_2350),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2788),
.Y(n_3191)
);

AND2x4_ASAP7_75t_L g3192 ( 
.A(n_2665),
.B(n_1962),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2798),
.B(n_1582),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2788),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2790),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2804),
.B(n_1636),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2790),
.Y(n_3197)
);

BUFx6f_ASAP7_75t_L g3198 ( 
.A(n_2610),
.Y(n_3198)
);

OR2x6_ASAP7_75t_L g3199 ( 
.A(n_2513),
.B(n_2155),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2804),
.B(n_2565),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_2863),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2565),
.B(n_2155),
.Y(n_3202)
);

OR2x2_ASAP7_75t_L g3203 ( 
.A(n_2647),
.B(n_2234),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2575),
.Y(n_3204)
);

CKINVDCx16_ASAP7_75t_R g3205 ( 
.A(n_2771),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2576),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_2863),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_L g3208 ( 
.A(n_2558),
.B(n_2374),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2637),
.B(n_1636),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2791),
.Y(n_3210)
);

CKINVDCx5p33_ASAP7_75t_R g3211 ( 
.A(n_2594),
.Y(n_3211)
);

INVx8_ASAP7_75t_L g3212 ( 
.A(n_2646),
.Y(n_3212)
);

BUFx10_ASAP7_75t_L g3213 ( 
.A(n_2653),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_2648),
.B(n_2681),
.Y(n_3214)
);

BUFx2_ASAP7_75t_L g3215 ( 
.A(n_2819),
.Y(n_3215)
);

BUFx3_ASAP7_75t_L g3216 ( 
.A(n_2544),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2576),
.Y(n_3217)
);

NOR2x1p5_ASAP7_75t_L g3218 ( 
.A(n_2650),
.B(n_2063),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2791),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_2648),
.B(n_1994),
.Y(n_3220)
);

AO22x2_ASAP7_75t_L g3221 ( 
.A1(n_2638),
.A2(n_1805),
.B1(n_1961),
.B2(n_1485),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_2723),
.B(n_2374),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_SL g3223 ( 
.A(n_2650),
.B(n_2209),
.Y(n_3223)
);

INVx3_ASAP7_75t_L g3224 ( 
.A(n_2868),
.Y(n_3224)
);

NAND2x1p5_ASAP7_75t_L g3225 ( 
.A(n_2868),
.B(n_2374),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2803),
.Y(n_3226)
);

BUFx6f_ASAP7_75t_L g3227 ( 
.A(n_2610),
.Y(n_3227)
);

BUFx6f_ASAP7_75t_L g3228 ( 
.A(n_2662),
.Y(n_3228)
);

NAND2xp33_ASAP7_75t_L g3229 ( 
.A(n_2646),
.B(n_2751),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2803),
.Y(n_3230)
);

NOR2xp33_ASAP7_75t_L g3231 ( 
.A(n_2689),
.B(n_2391),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2577),
.Y(n_3232)
);

AND2x6_ASAP7_75t_L g3233 ( 
.A(n_2875),
.B(n_2185),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2805),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_2577),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2805),
.Y(n_3236)
);

BUFx6f_ASAP7_75t_L g3237 ( 
.A(n_2662),
.Y(n_3237)
);

INVx3_ASAP7_75t_L g3238 ( 
.A(n_2868),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_SL g3239 ( 
.A(n_2521),
.B(n_2221),
.Y(n_3239)
);

BUFx6f_ASAP7_75t_L g3240 ( 
.A(n_2662),
.Y(n_3240)
);

OR2x2_ASAP7_75t_L g3241 ( 
.A(n_2900),
.B(n_1483),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_2681),
.B(n_1688),
.Y(n_3242)
);

BUFx3_ASAP7_75t_L g3243 ( 
.A(n_2506),
.Y(n_3243)
);

AO22x2_ASAP7_75t_L g3244 ( 
.A1(n_2655),
.A2(n_1486),
.B1(n_1522),
.B2(n_1521),
.Y(n_3244)
);

INVx3_ASAP7_75t_L g3245 ( 
.A(n_2662),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_2809),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2579),
.Y(n_3247)
);

INVx3_ASAP7_75t_L g3248 ( 
.A(n_2662),
.Y(n_3248)
);

BUFx6f_ASAP7_75t_L g3249 ( 
.A(n_2784),
.Y(n_3249)
);

AND2x4_ASAP7_75t_L g3250 ( 
.A(n_2506),
.B(n_1996),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2708),
.B(n_2068),
.Y(n_3251)
);

NOR2xp33_ASAP7_75t_SL g3252 ( 
.A(n_2739),
.B(n_2209),
.Y(n_3252)
);

OAI22xp33_ASAP7_75t_L g3253 ( 
.A1(n_2714),
.A2(n_744),
.B1(n_1239),
.B2(n_1064),
.Y(n_3253)
);

AND2x4_ASAP7_75t_L g3254 ( 
.A(n_2584),
.B(n_2003),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_SL g3255 ( 
.A(n_2739),
.B(n_2209),
.Y(n_3255)
);

AND2x4_ASAP7_75t_L g3256 ( 
.A(n_2584),
.B(n_2006),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2809),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_SL g3258 ( 
.A(n_2521),
.B(n_2221),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2579),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_2708),
.B(n_2391),
.Y(n_3260)
);

AND2x4_ASAP7_75t_L g3261 ( 
.A(n_2819),
.B(n_2831),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2810),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2583),
.Y(n_3263)
);

INVx8_ASAP7_75t_L g3264 ( 
.A(n_2646),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2810),
.Y(n_3265)
);

CKINVDCx5p33_ASAP7_75t_R g3266 ( 
.A(n_2747),
.Y(n_3266)
);

INVx4_ASAP7_75t_L g3267 ( 
.A(n_2864),
.Y(n_3267)
);

NOR2xp33_ASAP7_75t_L g3268 ( 
.A(n_2683),
.B(n_2391),
.Y(n_3268)
);

BUFx6f_ASAP7_75t_L g3269 ( 
.A(n_2784),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2487),
.B(n_2049),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_SL g3271 ( 
.A(n_2521),
.B(n_2221),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2816),
.Y(n_3272)
);

NOR2xp33_ASAP7_75t_L g3273 ( 
.A(n_2603),
.B(n_2308),
.Y(n_3273)
);

INVx4_ASAP7_75t_L g3274 ( 
.A(n_2864),
.Y(n_3274)
);

NOR2xp33_ASAP7_75t_L g3275 ( 
.A(n_2890),
.B(n_2828),
.Y(n_3275)
);

BUFx3_ASAP7_75t_L g3276 ( 
.A(n_2819),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2816),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_2820),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2499),
.B(n_2059),
.Y(n_3279)
);

BUFx6f_ASAP7_75t_L g3280 ( 
.A(n_2784),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_2583),
.Y(n_3281)
);

BUFx2_ASAP7_75t_L g3282 ( 
.A(n_2819),
.Y(n_3282)
);

AND2x4_ASAP7_75t_L g3283 ( 
.A(n_2831),
.B(n_1743),
.Y(n_3283)
);

INVx4_ASAP7_75t_L g3284 ( 
.A(n_2864),
.Y(n_3284)
);

AND2x6_ASAP7_75t_L g3285 ( 
.A(n_2876),
.B(n_2714),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_L g3286 ( 
.A(n_2835),
.B(n_2308),
.Y(n_3286)
);

AND2x4_ASAP7_75t_L g3287 ( 
.A(n_2831),
.B(n_1745),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2820),
.Y(n_3288)
);

OAI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2593),
.A2(n_2194),
.B1(n_2072),
.B2(n_2074),
.Y(n_3289)
);

INVx2_ASAP7_75t_SL g3290 ( 
.A(n_2760),
.Y(n_3290)
);

AND2x4_ASAP7_75t_L g3291 ( 
.A(n_2831),
.B(n_1748),
.Y(n_3291)
);

INVx2_ASAP7_75t_L g3292 ( 
.A(n_2585),
.Y(n_3292)
);

INVx3_ASAP7_75t_L g3293 ( 
.A(n_2784),
.Y(n_3293)
);

AND2x6_ASAP7_75t_L g3294 ( 
.A(n_2876),
.B(n_2186),
.Y(n_3294)
);

AND2x4_ASAP7_75t_L g3295 ( 
.A(n_2831),
.B(n_1752),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_2572),
.B(n_1688),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_2585),
.Y(n_3297)
);

OR2x2_ASAP7_75t_SL g3298 ( 
.A(n_2570),
.B(n_1861),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2897),
.B(n_2412),
.Y(n_3299)
);

AO22x2_ASAP7_75t_L g3300 ( 
.A1(n_2655),
.A2(n_1890),
.B1(n_2013),
.B2(n_1826),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_2592),
.Y(n_3301)
);

BUFx3_ASAP7_75t_L g3302 ( 
.A(n_2747),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_2592),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_2601),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_2601),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2829),
.Y(n_3306)
);

AND2x2_ASAP7_75t_L g3307 ( 
.A(n_2677),
.B(n_1692),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2829),
.Y(n_3308)
);

AND2x4_ASAP7_75t_L g3309 ( 
.A(n_2795),
.B(n_1760),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2551),
.B(n_2412),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_2832),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_SL g3312 ( 
.A(n_2545),
.B(n_2221),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2832),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2833),
.Y(n_3314)
);

INVx4_ASAP7_75t_L g3315 ( 
.A(n_2864),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_L g3316 ( 
.A(n_2796),
.B(n_2313),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_2892),
.B(n_1692),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2905),
.B(n_2414),
.Y(n_3318)
);

BUFx3_ASAP7_75t_L g3319 ( 
.A(n_2771),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2833),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_SL g3321 ( 
.A(n_2771),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2840),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2840),
.Y(n_3323)
);

AND2x6_ASAP7_75t_L g3324 ( 
.A(n_2772),
.B(n_2186),
.Y(n_3324)
);

AND2x6_ASAP7_75t_L g3325 ( 
.A(n_2772),
.B(n_2060),
.Y(n_3325)
);

NOR2xp33_ASAP7_75t_L g3326 ( 
.A(n_2800),
.B(n_2313),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_L g3327 ( 
.A(n_2827),
.B(n_2318),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_SL g3328 ( 
.A(n_2545),
.B(n_2240),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_2895),
.B(n_1693),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_2920),
.B(n_2517),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2727),
.B(n_2414),
.Y(n_3331)
);

NAND2x1p5_ASAP7_75t_L g3332 ( 
.A(n_2864),
.B(n_2240),
.Y(n_3332)
);

AND2x4_ASAP7_75t_L g3333 ( 
.A(n_2795),
.B(n_1761),
.Y(n_3333)
);

BUFx6f_ASAP7_75t_L g3334 ( 
.A(n_2784),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2843),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_2602),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_2857),
.B(n_2318),
.Y(n_3337)
);

AND2x4_ASAP7_75t_L g3338 ( 
.A(n_2919),
.B(n_1763),
.Y(n_3338)
);

INVx2_ASAP7_75t_SL g3339 ( 
.A(n_2760),
.Y(n_3339)
);

AND2x4_ASAP7_75t_L g3340 ( 
.A(n_2919),
.B(n_1765),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_2843),
.Y(n_3341)
);

BUFx2_ASAP7_75t_L g3342 ( 
.A(n_2906),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_2602),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_2613),
.Y(n_3344)
);

INVx4_ASAP7_75t_L g3345 ( 
.A(n_2864),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_2765),
.B(n_2321),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_2907),
.B(n_2561),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_2853),
.Y(n_3348)
);

NOR2xp33_ASAP7_75t_L g3349 ( 
.A(n_2773),
.B(n_2321),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2853),
.Y(n_3350)
);

INVx5_ASAP7_75t_L g3351 ( 
.A(n_2646),
.Y(n_3351)
);

NAND2x1p5_ASAP7_75t_L g3352 ( 
.A(n_2919),
.B(n_2240),
.Y(n_3352)
);

BUFx6f_ASAP7_75t_L g3353 ( 
.A(n_2807),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2854),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_2613),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_2750),
.B(n_2416),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2854),
.Y(n_3357)
);

AO22x2_ASAP7_75t_L g3358 ( 
.A1(n_2591),
.A2(n_1890),
.B1(n_2013),
.B2(n_1826),
.Y(n_3358)
);

INVxp67_ASAP7_75t_L g3359 ( 
.A(n_2657),
.Y(n_3359)
);

INVx4_ASAP7_75t_L g3360 ( 
.A(n_2605),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2855),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2855),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2856),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2856),
.Y(n_3364)
);

BUFx6f_ASAP7_75t_L g3365 ( 
.A(n_2807),
.Y(n_3365)
);

AND2x4_ASAP7_75t_L g3366 ( 
.A(n_2513),
.B(n_1766),
.Y(n_3366)
);

BUFx6f_ASAP7_75t_L g3367 ( 
.A(n_2807),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_2801),
.B(n_2416),
.Y(n_3368)
);

AND2x4_ASAP7_75t_L g3369 ( 
.A(n_2513),
.B(n_1768),
.Y(n_3369)
);

BUFx6f_ASAP7_75t_L g3370 ( 
.A(n_2807),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_2717),
.B(n_2744),
.Y(n_3371)
);

OAI22xp5_ASAP7_75t_SL g3372 ( 
.A1(n_2671),
.A2(n_1693),
.B1(n_1935),
.B2(n_1713),
.Y(n_3372)
);

BUFx4f_ASAP7_75t_L g3373 ( 
.A(n_2646),
.Y(n_3373)
);

INVx5_ASAP7_75t_L g3374 ( 
.A(n_2751),
.Y(n_3374)
);

BUFx6f_ASAP7_75t_L g3375 ( 
.A(n_2807),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_2762),
.B(n_2325),
.Y(n_3376)
);

BUFx2_ASAP7_75t_L g3377 ( 
.A(n_2906),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_2879),
.B(n_1713),
.Y(n_3378)
);

OR2x6_ASAP7_75t_L g3379 ( 
.A(n_2513),
.B(n_2771),
.Y(n_3379)
);

INVx2_ASAP7_75t_SL g3380 ( 
.A(n_2760),
.Y(n_3380)
);

BUFx6f_ASAP7_75t_L g3381 ( 
.A(n_2873),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_2616),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2861),
.Y(n_3383)
);

NOR2xp33_ASAP7_75t_R g3384 ( 
.A(n_2498),
.B(n_1935),
.Y(n_3384)
);

AND2x6_ASAP7_75t_L g3385 ( 
.A(n_2836),
.B(n_2060),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_2563),
.B(n_1775),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_2616),
.Y(n_3387)
);

BUFx6f_ASAP7_75t_L g3388 ( 
.A(n_2873),
.Y(n_3388)
);

AND2x4_ASAP7_75t_L g3389 ( 
.A(n_2563),
.B(n_1777),
.Y(n_3389)
);

AND2x4_ASAP7_75t_L g3390 ( 
.A(n_2906),
.B(n_1797),
.Y(n_3390)
);

INVx1_ASAP7_75t_SL g3391 ( 
.A(n_2906),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_2629),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_L g3393 ( 
.A(n_2813),
.B(n_2325),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2929),
.B(n_2870),
.Y(n_3394)
);

AND2x4_ASAP7_75t_L g3395 ( 
.A(n_3002),
.B(n_2906),
.Y(n_3395)
);

INVxp67_ASAP7_75t_L g3396 ( 
.A(n_3054),
.Y(n_3396)
);

INVx8_ASAP7_75t_L g3397 ( 
.A(n_3261),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_2929),
.B(n_2913),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_2928),
.B(n_2625),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2928),
.B(n_2635),
.Y(n_3400)
);

NAND2xp33_ASAP7_75t_L g3401 ( 
.A(n_3212),
.B(n_2751),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2931),
.Y(n_3402)
);

O2A1O1Ixp33_ASAP7_75t_L g3403 ( 
.A1(n_2958),
.A2(n_2823),
.B(n_2704),
.C(n_2695),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3064),
.B(n_2927),
.Y(n_3404)
);

NOR2xp33_ASAP7_75t_L g3405 ( 
.A(n_3028),
.B(n_2813),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_2931),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3214),
.B(n_2532),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_3275),
.B(n_2908),
.Y(n_3408)
);

NOR2xp33_ASAP7_75t_L g3409 ( 
.A(n_3275),
.B(n_2908),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2954),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3034),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3118),
.B(n_2532),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3043),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2935),
.B(n_3222),
.Y(n_3414)
);

INVx2_ASAP7_75t_SL g3415 ( 
.A(n_2968),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3222),
.B(n_2757),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3065),
.B(n_2753),
.Y(n_3417)
);

BUFx2_ASAP7_75t_L g3418 ( 
.A(n_3105),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3053),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2949),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_SL g3421 ( 
.A(n_2999),
.B(n_2873),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_2934),
.Y(n_3422)
);

XOR2xp5_ASAP7_75t_L g3423 ( 
.A(n_3266),
.B(n_2052),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3087),
.B(n_2763),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_SL g3425 ( 
.A(n_2999),
.B(n_2873),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_2934),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2950),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_2936),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2955),
.Y(n_3429)
);

NAND2x1p5_ASAP7_75t_L g3430 ( 
.A(n_3169),
.B(n_3187),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_2963),
.Y(n_3431)
);

INVxp67_ASAP7_75t_L g3432 ( 
.A(n_3005),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3143),
.B(n_2571),
.Y(n_3433)
);

AND2x6_ASAP7_75t_SL g3434 ( 
.A(n_3209),
.B(n_2771),
.Y(n_3434)
);

NOR2xp67_ASAP7_75t_L g3435 ( 
.A(n_3049),
.B(n_2608),
.Y(n_3435)
);

AOI22xp33_ASAP7_75t_L g3436 ( 
.A1(n_2942),
.A2(n_2541),
.B1(n_2566),
.B2(n_2543),
.Y(n_3436)
);

INVx2_ASAP7_75t_L g3437 ( 
.A(n_2936),
.Y(n_3437)
);

AND2x2_ASAP7_75t_L g3438 ( 
.A(n_2953),
.B(n_2933),
.Y(n_3438)
);

NOR2x1p5_ASAP7_75t_L g3439 ( 
.A(n_3049),
.B(n_2235),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_3296),
.B(n_2850),
.Y(n_3440)
);

NOR3x1_ASAP7_75t_L g3441 ( 
.A(n_3026),
.B(n_2651),
.C(n_2674),
.Y(n_3441)
);

AOI22xp5_ASAP7_75t_L g3442 ( 
.A1(n_3307),
.A2(n_2908),
.B1(n_2850),
.B2(n_2872),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3200),
.B(n_2746),
.Y(n_3443)
);

INVx8_ASAP7_75t_L g3444 ( 
.A(n_3261),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_SL g3445 ( 
.A(n_2999),
.B(n_2873),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_2967),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_L g3447 ( 
.A(n_2939),
.B(n_2641),
.Y(n_3447)
);

INVx4_ASAP7_75t_L g3448 ( 
.A(n_3091),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_3000),
.B(n_2614),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3076),
.B(n_2719),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3109),
.B(n_2668),
.Y(n_3451)
);

OR2x2_ASAP7_75t_L g3452 ( 
.A(n_2932),
.B(n_2052),
.Y(n_3452)
);

NOR2xp67_ASAP7_75t_L g3453 ( 
.A(n_3266),
.B(n_2619),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_2970),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_2942),
.A2(n_3253),
.B1(n_2978),
.B2(n_3126),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_SL g3456 ( 
.A(n_2999),
.B(n_2557),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3040),
.B(n_2697),
.Y(n_3457)
);

AND2x4_ASAP7_75t_L g3458 ( 
.A(n_3002),
.B(n_2749),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3220),
.B(n_3251),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3220),
.B(n_3056),
.Y(n_3460)
);

BUFx8_ASAP7_75t_L g3461 ( 
.A(n_3321),
.Y(n_3461)
);

OAI22xp5_ASAP7_75t_L g3462 ( 
.A1(n_2958),
.A2(n_2812),
.B1(n_2817),
.B2(n_2672),
.Y(n_3462)
);

INVx2_ASAP7_75t_SL g3463 ( 
.A(n_2968),
.Y(n_3463)
);

BUFx6f_ASAP7_75t_L g3464 ( 
.A(n_2941),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2977),
.Y(n_3465)
);

NOR2xp33_ASAP7_75t_L g3466 ( 
.A(n_3000),
.B(n_2597),
.Y(n_3466)
);

NAND3xp33_ASAP7_75t_L g3467 ( 
.A(n_3048),
.B(n_2055),
.C(n_2041),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_2999),
.B(n_2557),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_2983),
.Y(n_3469)
);

INVx3_ASAP7_75t_L g3470 ( 
.A(n_3169),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3056),
.B(n_3092),
.Y(n_3471)
);

INVx3_ASAP7_75t_L g3472 ( 
.A(n_3169),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_2938),
.Y(n_3473)
);

OAI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3149),
.A2(n_2534),
.B(n_2705),
.Y(n_3474)
);

NOR2xp67_ASAP7_75t_L g3475 ( 
.A(n_3359),
.B(n_2847),
.Y(n_3475)
);

INVxp67_ASAP7_75t_L g3476 ( 
.A(n_3033),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3056),
.B(n_2566),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_2989),
.B(n_2597),
.Y(n_3478)
);

AND2x6_ASAP7_75t_SL g3479 ( 
.A(n_3186),
.B(n_1879),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3092),
.B(n_2595),
.Y(n_3480)
);

BUFx6f_ASAP7_75t_L g3481 ( 
.A(n_2941),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3092),
.B(n_2595),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3038),
.B(n_2624),
.Y(n_3483)
);

OAI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_3241),
.A2(n_744),
.B1(n_816),
.B2(n_751),
.Y(n_3484)
);

AOI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_2978),
.A2(n_2541),
.B1(n_2569),
.B2(n_2543),
.Y(n_3485)
);

NAND3xp33_ASAP7_75t_L g3486 ( 
.A(n_3048),
.B(n_3193),
.C(n_3150),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3140),
.B(n_2617),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_2987),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_2938),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_2965),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_2965),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_2990),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_2943),
.B(n_2617),
.Y(n_3493)
);

OAI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_3260),
.A2(n_2866),
.B(n_2814),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2996),
.Y(n_3495)
);

NOR2x2_ASAP7_75t_L g3496 ( 
.A(n_3379),
.B(n_1879),
.Y(n_3496)
);

AND2x6_ASAP7_75t_SL g3497 ( 
.A(n_3378),
.B(n_1915),
.Y(n_3497)
);

NAND2x1_ASAP7_75t_L g3498 ( 
.A(n_3267),
.B(n_2597),
.Y(n_3498)
);

INVx2_ASAP7_75t_SL g3499 ( 
.A(n_2973),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_SL g3500 ( 
.A(n_3008),
.B(n_2882),
.Y(n_3500)
);

A2O1A1Ixp33_ASAP7_75t_SL g3501 ( 
.A1(n_3102),
.A2(n_2706),
.B(n_2764),
.C(n_2669),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_2945),
.B(n_2624),
.Y(n_3502)
);

INVx4_ASAP7_75t_L g3503 ( 
.A(n_3091),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_2969),
.B(n_2628),
.Y(n_3504)
);

INVx4_ASAP7_75t_L g3505 ( 
.A(n_3091),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_2972),
.B(n_2628),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3008),
.B(n_2882),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_SL g3508 ( 
.A(n_3008),
.B(n_2569),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_2984),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_2997),
.B(n_2669),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_2984),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_2980),
.B(n_2588),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_2985),
.B(n_2588),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3017),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_SL g3515 ( 
.A(n_3223),
.B(n_2235),
.Y(n_3515)
);

A2O1A1Ixp33_ASAP7_75t_L g3516 ( 
.A1(n_3133),
.A2(n_3150),
.B(n_3330),
.C(n_3001),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_2991),
.B(n_2598),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_2997),
.B(n_2669),
.Y(n_3518)
);

XNOR2xp5_ASAP7_75t_L g3519 ( 
.A(n_3358),
.B(n_2858),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3008),
.B(n_2580),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3004),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_3052),
.B(n_3055),
.Y(n_3522)
);

AOI22xp5_ASAP7_75t_L g3523 ( 
.A1(n_3347),
.A2(n_2013),
.B1(n_1890),
.B2(n_2041),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3009),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_2994),
.B(n_2611),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_2947),
.B(n_2706),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3013),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_2947),
.B(n_2706),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3015),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3020),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3011),
.B(n_2611),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_SL g3532 ( 
.A(n_3008),
.B(n_2580),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3017),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3029),
.Y(n_3534)
);

OR2x2_ASAP7_75t_L g3535 ( 
.A(n_3242),
.B(n_2918),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3042),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3046),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3018),
.B(n_2702),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3035),
.B(n_3072),
.Y(n_3539)
);

O2A1O1Ixp33_ASAP7_75t_L g3540 ( 
.A1(n_3163),
.A2(n_904),
.B(n_1811),
.C(n_1803),
.Y(n_3540)
);

BUFx6f_ASAP7_75t_SL g3541 ( 
.A(n_3302),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_3016),
.B(n_2598),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3016),
.B(n_2604),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3072),
.B(n_2632),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3088),
.B(n_3371),
.Y(n_3545)
);

OAI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3045),
.A2(n_2841),
.B1(n_2759),
.B2(n_2761),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3167),
.B(n_2509),
.Y(n_3547)
);

OR2x2_ASAP7_75t_L g3548 ( 
.A(n_3196),
.B(n_3027),
.Y(n_3548)
);

AO22x1_ASAP7_75t_L g3549 ( 
.A1(n_3317),
.A2(n_2055),
.B1(n_2288),
.B2(n_2235),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3088),
.B(n_2604),
.Y(n_3550)
);

AOI22xp5_ASAP7_75t_L g3551 ( 
.A1(n_3001),
.A2(n_2055),
.B1(n_2306),
.B2(n_2288),
.Y(n_3551)
);

HB1xp67_ASAP7_75t_L g3552 ( 
.A(n_2973),
.Y(n_3552)
);

INVxp67_ASAP7_75t_SL g3553 ( 
.A(n_3229),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3019),
.Y(n_3554)
);

BUFx6f_ASAP7_75t_L g3555 ( 
.A(n_2941),
.Y(n_3555)
);

AND2x4_ASAP7_75t_L g3556 ( 
.A(n_3002),
.B(n_2749),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_SL g3557 ( 
.A(n_3016),
.B(n_3077),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3051),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3058),
.Y(n_3559)
);

A2O1A1Ixp33_ASAP7_75t_L g3560 ( 
.A1(n_3133),
.A2(n_2573),
.B(n_2633),
.C(n_2632),
.Y(n_3560)
);

NAND2x1p5_ASAP7_75t_L g3561 ( 
.A(n_3187),
.B(n_2759),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3088),
.B(n_2732),
.Y(n_3562)
);

NOR2xp33_ASAP7_75t_L g3563 ( 
.A(n_3080),
.B(n_2764),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3068),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3069),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3202),
.B(n_2732),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3070),
.Y(n_3567)
);

AOI22xp33_ASAP7_75t_L g3568 ( 
.A1(n_2978),
.A2(n_2633),
.B1(n_2649),
.B2(n_2643),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3071),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_L g3570 ( 
.A(n_3145),
.B(n_2764),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3019),
.Y(n_3571)
);

O2A1O1Ixp5_ASAP7_75t_L g3572 ( 
.A1(n_3102),
.A2(n_2824),
.B(n_2649),
.C(n_2654),
.Y(n_3572)
);

AOI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3329),
.A2(n_3160),
.B1(n_3211),
.B2(n_3113),
.Y(n_3573)
);

NAND2xp33_ASAP7_75t_SL g3574 ( 
.A(n_3025),
.B(n_2761),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3021),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3073),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_3021),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3202),
.B(n_2643),
.Y(n_3578)
);

CKINVDCx5p33_ASAP7_75t_R g3579 ( 
.A(n_3124),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3022),
.Y(n_3580)
);

AND2x4_ASAP7_75t_L g3581 ( 
.A(n_3276),
.B(n_2834),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_SL g3582 ( 
.A(n_3016),
.B(n_2654),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_L g3583 ( 
.A(n_3099),
.B(n_2767),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_L g3584 ( 
.A(n_3099),
.B(n_2767),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3078),
.Y(n_3585)
);

OR2x2_ASAP7_75t_L g3586 ( 
.A(n_3172),
.B(n_1915),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3286),
.B(n_3270),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3081),
.Y(n_3588)
);

OAI22xp33_ASAP7_75t_L g3589 ( 
.A1(n_3148),
.A2(n_968),
.B1(n_974),
.B2(n_890),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_3022),
.Y(n_3590)
);

NOR3xp33_ASAP7_75t_SL g3591 ( 
.A(n_3113),
.B(n_810),
.C(n_706),
.Y(n_3591)
);

OAI22x1_ASAP7_75t_L g3592 ( 
.A1(n_3261),
.A2(n_1930),
.B1(n_2014),
.B2(n_2010),
.Y(n_3592)
);

NOR3xp33_ASAP7_75t_L g3593 ( 
.A(n_3132),
.B(n_1822),
.C(n_1812),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3286),
.B(n_2702),
.Y(n_3594)
);

INVx4_ASAP7_75t_L g3595 ( 
.A(n_3187),
.Y(n_3595)
);

CKINVDCx16_ASAP7_75t_R g3596 ( 
.A(n_3252),
.Y(n_3596)
);

NOR2xp67_ASAP7_75t_L g3597 ( 
.A(n_3160),
.B(n_2847),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3121),
.B(n_2661),
.Y(n_3598)
);

BUFx3_ASAP7_75t_L g3599 ( 
.A(n_2974),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3093),
.B(n_2509),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3116),
.B(n_2661),
.Y(n_3601)
);

BUFx6f_ASAP7_75t_L g3602 ( 
.A(n_2941),
.Y(n_3602)
);

AND2x4_ASAP7_75t_L g3603 ( 
.A(n_3276),
.B(n_2834),
.Y(n_3603)
);

NAND2xp33_ASAP7_75t_L g3604 ( 
.A(n_3212),
.B(n_2751),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3023),
.Y(n_3605)
);

NAND2xp33_ASAP7_75t_L g3606 ( 
.A(n_3212),
.B(n_2751),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3116),
.B(n_2707),
.Y(n_3607)
);

INVx3_ASAP7_75t_L g3608 ( 
.A(n_3267),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3082),
.Y(n_3609)
);

INVx4_ASAP7_75t_L g3610 ( 
.A(n_3124),
.Y(n_3610)
);

OAI22xp33_ASAP7_75t_L g3611 ( 
.A1(n_3255),
.A2(n_968),
.B1(n_974),
.B2(n_890),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3116),
.B(n_2664),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3127),
.B(n_2664),
.Y(n_3613)
);

NOR2xp33_ASAP7_75t_L g3614 ( 
.A(n_3203),
.B(n_2767),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3127),
.B(n_2666),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3127),
.B(n_2666),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3302),
.B(n_2509),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_SL g3618 ( 
.A(n_3016),
.B(n_3077),
.Y(n_3618)
);

AOI21xp5_ASAP7_75t_L g3619 ( 
.A1(n_2946),
.A2(n_2709),
.B(n_2667),
.Y(n_3619)
);

NAND3xp33_ASAP7_75t_SL g3620 ( 
.A(n_3211),
.B(n_1181),
.C(n_1146),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3045),
.B(n_2707),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3023),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2946),
.A2(n_3229),
.B(n_3289),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_SL g3624 ( 
.A(n_3077),
.B(n_2680),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3126),
.B(n_2710),
.Y(n_3625)
);

AOI22xp33_ASAP7_75t_L g3626 ( 
.A1(n_3244),
.A2(n_2680),
.B1(n_2696),
.B2(n_2686),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3083),
.Y(n_3627)
);

NOR2xp33_ASAP7_75t_L g3628 ( 
.A(n_3177),
.B(n_2781),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3090),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3024),
.Y(n_3630)
);

NOR3x1_ASAP7_75t_L g3631 ( 
.A(n_3060),
.B(n_969),
.C(n_967),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3279),
.B(n_2696),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3180),
.B(n_2698),
.Y(n_3633)
);

O2A1O1Ixp5_ASAP7_75t_L g3634 ( 
.A1(n_3132),
.A2(n_3231),
.B(n_3258),
.C(n_3239),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3180),
.B(n_2698),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3180),
.B(n_2715),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3176),
.B(n_2509),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_L g3638 ( 
.A(n_3177),
.B(n_2781),
.Y(n_3638)
);

A2O1A1Ixp33_ASAP7_75t_L g3639 ( 
.A1(n_3373),
.A2(n_2700),
.B(n_2701),
.C(n_2686),
.Y(n_3639)
);

NOR2x2_ASAP7_75t_L g3640 ( 
.A(n_3379),
.B(n_1930),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3024),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3098),
.Y(n_3642)
);

BUFx3_ASAP7_75t_L g3643 ( 
.A(n_2974),
.Y(n_3643)
);

AOI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_3111),
.A2(n_2351),
.B1(n_2306),
.B2(n_2288),
.Y(n_3644)
);

AOI221xp5_ASAP7_75t_L g3645 ( 
.A1(n_3358),
.A2(n_1663),
.B1(n_1152),
.B2(n_1169),
.C(n_1064),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3108),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3117),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3137),
.Y(n_3648)
);

AOI21xp5_ASAP7_75t_L g3649 ( 
.A1(n_3373),
.A2(n_2194),
.B(n_2785),
.Y(n_3649)
);

AOI22xp33_ASAP7_75t_L g3650 ( 
.A1(n_3244),
.A2(n_2700),
.B1(n_2710),
.B2(n_2701),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3155),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3185),
.B(n_3192),
.Y(n_3652)
);

CKINVDCx5p33_ASAP7_75t_R g3653 ( 
.A(n_2975),
.Y(n_3653)
);

AOI22xp33_ASAP7_75t_L g3654 ( 
.A1(n_3244),
.A2(n_2711),
.B1(n_2715),
.B2(n_2712),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_3208),
.B(n_2781),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3037),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3037),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3157),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3185),
.B(n_2711),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3161),
.Y(n_3660)
);

AOI22xp33_ASAP7_75t_L g3661 ( 
.A1(n_2952),
.A2(n_2712),
.B1(n_2722),
.B2(n_2718),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_3047),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3164),
.Y(n_3663)
);

OR2x6_ASAP7_75t_L g3664 ( 
.A(n_3199),
.B(n_2688),
.Y(n_3664)
);

OR2x2_ASAP7_75t_L g3665 ( 
.A(n_3372),
.B(n_2014),
.Y(n_3665)
);

AOI22xp33_ASAP7_75t_L g3666 ( 
.A1(n_2952),
.A2(n_2718),
.B1(n_2724),
.B2(n_2722),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3047),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3185),
.B(n_2728),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3192),
.B(n_2728),
.Y(n_3669)
);

AOI22xp33_ASAP7_75t_SL g3670 ( 
.A1(n_3358),
.A2(n_2688),
.B1(n_2306),
.B2(n_2408),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3192),
.B(n_3208),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3168),
.Y(n_3672)
);

BUFx6f_ASAP7_75t_L g3673 ( 
.A(n_2964),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3171),
.Y(n_3674)
);

NOR2xp33_ASAP7_75t_L g3675 ( 
.A(n_3170),
.B(n_2793),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3170),
.B(n_2793),
.Y(n_3676)
);

NOR2xp33_ASAP7_75t_L g3677 ( 
.A(n_3170),
.B(n_2793),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_SL g3678 ( 
.A(n_3077),
.B(n_3120),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_SL g3679 ( 
.A(n_3077),
.B(n_2724),
.Y(n_3679)
);

INVx3_ASAP7_75t_L g3680 ( 
.A(n_3267),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3243),
.B(n_2726),
.Y(n_3681)
);

INVx4_ASAP7_75t_L g3682 ( 
.A(n_3152),
.Y(n_3682)
);

INVx2_ASAP7_75t_SL g3683 ( 
.A(n_2975),
.Y(n_3683)
);

NOR2xp33_ASAP7_75t_L g3684 ( 
.A(n_3213),
.B(n_2799),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3243),
.B(n_2726),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3141),
.B(n_2688),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3174),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_SL g3688 ( 
.A(n_3120),
.B(n_2734),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3215),
.B(n_2688),
.Y(n_3689)
);

AND2x6_ASAP7_75t_L g3690 ( 
.A(n_3224),
.B(n_2836),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3250),
.B(n_2734),
.Y(n_3691)
);

INVx2_ASAP7_75t_SL g3692 ( 
.A(n_3012),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3250),
.B(n_2861),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3250),
.B(n_2865),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3254),
.B(n_2865),
.Y(n_3695)
);

AND2x6_ASAP7_75t_SL g3696 ( 
.A(n_3379),
.B(n_2010),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3213),
.B(n_2799),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3254),
.B(n_2869),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3050),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3050),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3254),
.B(n_2869),
.Y(n_3701)
);

AOI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_3373),
.A2(n_2808),
.B(n_2806),
.Y(n_3702)
);

NOR2xp33_ASAP7_75t_L g3703 ( 
.A(n_3213),
.B(n_2799),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3178),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3066),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3189),
.Y(n_3706)
);

INVx2_ASAP7_75t_L g3707 ( 
.A(n_3066),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3256),
.B(n_2871),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3256),
.B(n_2871),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3256),
.B(n_2877),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3299),
.B(n_3191),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3075),
.Y(n_3712)
);

NOR2xp33_ASAP7_75t_L g3713 ( 
.A(n_3006),
.B(n_2818),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3194),
.B(n_3195),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_SL g3715 ( 
.A(n_3120),
.B(n_2818),
.Y(n_3715)
);

NOR3xp33_ASAP7_75t_L g3716 ( 
.A(n_3268),
.B(n_1827),
.C(n_1823),
.Y(n_3716)
);

INVxp33_ASAP7_75t_SL g3717 ( 
.A(n_3384),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3197),
.Y(n_3718)
);

BUFx3_ASAP7_75t_L g3719 ( 
.A(n_3012),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3075),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3210),
.Y(n_3721)
);

AND2x4_ASAP7_75t_L g3722 ( 
.A(n_3199),
.B(n_2818),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3219),
.B(n_2877),
.Y(n_3723)
);

NOR2xp67_ASAP7_75t_L g3724 ( 
.A(n_3158),
.B(n_2794),
.Y(n_3724)
);

NOR2xp33_ASAP7_75t_L g3725 ( 
.A(n_3006),
.B(n_2852),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3226),
.B(n_2880),
.Y(n_3726)
);

INVx2_ASAP7_75t_L g3727 ( 
.A(n_3085),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3230),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3282),
.B(n_1609),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3239),
.A2(n_2848),
.B(n_2846),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_L g3731 ( 
.A1(n_2952),
.A2(n_2883),
.B1(n_2887),
.B2(n_2878),
.Y(n_3731)
);

BUFx3_ASAP7_75t_L g3732 ( 
.A(n_3041),
.Y(n_3732)
);

AOI22xp5_ASAP7_75t_L g3733 ( 
.A1(n_3111),
.A2(n_2408),
.B1(n_2351),
.B2(n_2794),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3234),
.Y(n_3734)
);

INVx2_ASAP7_75t_L g3735 ( 
.A(n_3085),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3236),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3246),
.B(n_2880),
.Y(n_3737)
);

INVx2_ASAP7_75t_SL g3738 ( 
.A(n_3041),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3257),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3262),
.B(n_3265),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3095),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3095),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_SL g3743 ( 
.A(n_3120),
.B(n_2852),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3272),
.B(n_2885),
.Y(n_3744)
);

OAI22xp5_ASAP7_75t_L g3745 ( 
.A1(n_3025),
.A2(n_2867),
.B1(n_2881),
.B2(n_2852),
.Y(n_3745)
);

AND2x2_ASAP7_75t_SL g3746 ( 
.A(n_3205),
.B(n_2885),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3277),
.B(n_2886),
.Y(n_3747)
);

AND2x6_ASAP7_75t_SL g3748 ( 
.A(n_3379),
.B(n_2351),
.Y(n_3748)
);

AND2x4_ASAP7_75t_L g3749 ( 
.A(n_3199),
.B(n_2545),
.Y(n_3749)
);

INVxp33_ASAP7_75t_L g3750 ( 
.A(n_3384),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3278),
.B(n_2886),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3288),
.B(n_2889),
.Y(n_3752)
);

AOI22xp5_ASAP7_75t_L g3753 ( 
.A1(n_3111),
.A2(n_2408),
.B1(n_2751),
.B2(n_2586),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_SL g3754 ( 
.A(n_3120),
.B(n_2889),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3306),
.B(n_2899),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3308),
.B(n_2899),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3311),
.B(n_3313),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3314),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3104),
.Y(n_3759)
);

INVxp33_ASAP7_75t_L g3760 ( 
.A(n_3006),
.Y(n_3760)
);

AND2x2_ASAP7_75t_L g3761 ( 
.A(n_3221),
.B(n_1610),
.Y(n_3761)
);

NOR2x1_ASAP7_75t_R g3762 ( 
.A(n_3309),
.B(n_706),
.Y(n_3762)
);

OAI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3139),
.A2(n_2909),
.B(n_2901),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3320),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3104),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3322),
.Y(n_3766)
);

AOI22xp33_ASAP7_75t_L g3767 ( 
.A1(n_2940),
.A2(n_2883),
.B1(n_2887),
.B2(n_2878),
.Y(n_3767)
);

XOR2xp5_ASAP7_75t_L g3768 ( 
.A(n_3300),
.B(n_1587),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3323),
.B(n_2901),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3335),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3341),
.B(n_2909),
.Y(n_3771)
);

AOI22xp5_ASAP7_75t_L g3772 ( 
.A1(n_3110),
.A2(n_2751),
.B1(n_2581),
.B2(n_2658),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3348),
.B(n_2912),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_SL g3774 ( 
.A(n_3183),
.B(n_2912),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3107),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3350),
.B(n_2914),
.Y(n_3776)
);

AOI22xp5_ASAP7_75t_L g3777 ( 
.A1(n_3110),
.A2(n_3391),
.B1(n_3031),
.B2(n_3377),
.Y(n_3777)
);

INVx2_ASAP7_75t_SL g3778 ( 
.A(n_3218),
.Y(n_3778)
);

AND2x2_ASAP7_75t_SL g3779 ( 
.A(n_3342),
.B(n_2914),
.Y(n_3779)
);

NOR2xp33_ASAP7_75t_L g3780 ( 
.A(n_3031),
.B(n_3089),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3354),
.B(n_2915),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3107),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3357),
.Y(n_3783)
);

AOI22xp33_ASAP7_75t_L g3784 ( 
.A1(n_2940),
.A2(n_2893),
.B1(n_2894),
.B2(n_2888),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3183),
.B(n_2915),
.Y(n_3785)
);

AO22x1_ASAP7_75t_L g3786 ( 
.A1(n_3309),
.A2(n_1187),
.B1(n_1152),
.B2(n_1169),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3361),
.Y(n_3787)
);

AOI21xp5_ASAP7_75t_L g3788 ( 
.A1(n_3258),
.A2(n_2072),
.B(n_2074),
.Y(n_3788)
);

AOI22xp33_ASAP7_75t_L g3789 ( 
.A1(n_2940),
.A2(n_2893),
.B1(n_2894),
.B2(n_2888),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3114),
.Y(n_3790)
);

O2A1O1Ixp33_ASAP7_75t_L g3791 ( 
.A1(n_3268),
.A2(n_1831),
.B(n_1212),
.C(n_1239),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3438),
.B(n_3221),
.Y(n_3792)
);

INVx2_ASAP7_75t_SL g3793 ( 
.A(n_3653),
.Y(n_3793)
);

AOI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3486),
.A2(n_3283),
.B1(n_3291),
.B2(n_3287),
.Y(n_3794)
);

HB1xp67_ASAP7_75t_L g3795 ( 
.A(n_3552),
.Y(n_3795)
);

AND2x4_ASAP7_75t_L g3796 ( 
.A(n_3395),
.B(n_3199),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3402),
.Y(n_3797)
);

AOI22xp33_ASAP7_75t_L g3798 ( 
.A1(n_3455),
.A2(n_3221),
.B1(n_3300),
.B2(n_3386),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3420),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3414),
.B(n_3285),
.Y(n_3800)
);

BUFx6f_ASAP7_75t_L g3801 ( 
.A(n_3397),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3427),
.Y(n_3802)
);

BUFx6f_ASAP7_75t_L g3803 ( 
.A(n_3397),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3429),
.Y(n_3804)
);

HB1xp67_ASAP7_75t_L g3805 ( 
.A(n_3552),
.Y(n_3805)
);

INVx2_ASAP7_75t_L g3806 ( 
.A(n_3406),
.Y(n_3806)
);

BUFx3_ASAP7_75t_L g3807 ( 
.A(n_3418),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3431),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3446),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3454),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3423),
.B(n_3089),
.Y(n_3811)
);

NOR2xp33_ASAP7_75t_L g3812 ( 
.A(n_3408),
.B(n_3089),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3465),
.Y(n_3813)
);

BUFx6f_ASAP7_75t_L g3814 ( 
.A(n_3397),
.Y(n_3814)
);

NOR2xp33_ASAP7_75t_R g3815 ( 
.A(n_3579),
.B(n_3321),
.Y(n_3815)
);

BUFx6f_ASAP7_75t_L g3816 ( 
.A(n_3444),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3469),
.Y(n_3817)
);

HB1xp67_ASAP7_75t_L g3818 ( 
.A(n_3566),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3488),
.Y(n_3819)
);

OR2x4_ASAP7_75t_L g3820 ( 
.A(n_3620),
.B(n_3231),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3492),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3587),
.B(n_3516),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3516),
.B(n_3285),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3495),
.Y(n_3824)
);

INVx4_ASAP7_75t_L g3825 ( 
.A(n_3541),
.Y(n_3825)
);

OR2x6_ASAP7_75t_L g3826 ( 
.A(n_3444),
.B(n_3212),
.Y(n_3826)
);

BUFx3_ASAP7_75t_L g3827 ( 
.A(n_3599),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3521),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3440),
.B(n_3386),
.Y(n_3829)
);

INVx3_ASAP7_75t_L g3830 ( 
.A(n_3595),
.Y(n_3830)
);

AOI22xp5_ASAP7_75t_L g3831 ( 
.A1(n_3408),
.A2(n_3409),
.B1(n_3394),
.B2(n_3398),
.Y(n_3831)
);

INVx5_ASAP7_75t_L g3832 ( 
.A(n_3444),
.Y(n_3832)
);

CKINVDCx8_ASAP7_75t_R g3833 ( 
.A(n_3479),
.Y(n_3833)
);

INVx2_ASAP7_75t_L g3834 ( 
.A(n_3422),
.Y(n_3834)
);

BUFx3_ASAP7_75t_L g3835 ( 
.A(n_3599),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3426),
.Y(n_3836)
);

INVx4_ASAP7_75t_L g3837 ( 
.A(n_3541),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_SL g3838 ( 
.A(n_3399),
.B(n_2930),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3524),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3527),
.Y(n_3840)
);

NOR2xp33_ASAP7_75t_L g3841 ( 
.A(n_3409),
.B(n_3283),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3400),
.B(n_3779),
.Y(n_3842)
);

HB1xp67_ASAP7_75t_L g3843 ( 
.A(n_3578),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3529),
.Y(n_3844)
);

AOI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3405),
.A2(n_3283),
.B1(n_3291),
.B2(n_3287),
.Y(n_3845)
);

BUFx6f_ASAP7_75t_L g3846 ( 
.A(n_3643),
.Y(n_3846)
);

BUFx2_ASAP7_75t_L g3847 ( 
.A(n_3432),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3632),
.B(n_3285),
.Y(n_3848)
);

AND2x2_ASAP7_75t_SL g3849 ( 
.A(n_3455),
.B(n_3779),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3428),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3530),
.Y(n_3851)
);

BUFx2_ASAP7_75t_L g3852 ( 
.A(n_3476),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3449),
.B(n_3287),
.Y(n_3853)
);

O2A1O1Ixp33_ASAP7_75t_SL g3854 ( 
.A1(n_3501),
.A2(n_3290),
.B(n_3380),
.C(n_3339),
.Y(n_3854)
);

BUFx2_ASAP7_75t_L g3855 ( 
.A(n_3643),
.Y(n_3855)
);

HB1xp67_ASAP7_75t_L g3856 ( 
.A(n_3480),
.Y(n_3856)
);

INVx5_ASAP7_75t_L g3857 ( 
.A(n_3690),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3412),
.B(n_3285),
.Y(n_3858)
);

OR2x6_ASAP7_75t_L g3859 ( 
.A(n_3652),
.B(n_3264),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_SL g3860 ( 
.A(n_3459),
.B(n_3449),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3534),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3536),
.Y(n_3862)
);

NOR2x1p5_ASAP7_75t_L g3863 ( 
.A(n_3610),
.B(n_3319),
.Y(n_3863)
);

INVx5_ASAP7_75t_L g3864 ( 
.A(n_3690),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3711),
.B(n_3285),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3537),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3611),
.B(n_2930),
.Y(n_3867)
);

INVx4_ASAP7_75t_L g3868 ( 
.A(n_3448),
.Y(n_3868)
);

AOI22xp33_ASAP7_75t_L g3869 ( 
.A1(n_3589),
.A2(n_3300),
.B1(n_3285),
.B2(n_2940),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3729),
.B(n_3386),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3558),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3559),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3564),
.Y(n_3873)
);

INVx1_ASAP7_75t_SL g3874 ( 
.A(n_3548),
.Y(n_3874)
);

BUFx12f_ASAP7_75t_L g3875 ( 
.A(n_3610),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3565),
.Y(n_3876)
);

AND2x6_ASAP7_75t_L g3877 ( 
.A(n_3749),
.B(n_3224),
.Y(n_3877)
);

AO22x1_ASAP7_75t_L g3878 ( 
.A1(n_3461),
.A2(n_3319),
.B1(n_3369),
.B2(n_3366),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3437),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3473),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3567),
.Y(n_3881)
);

INVxp67_ASAP7_75t_L g3882 ( 
.A(n_3522),
.Y(n_3882)
);

NOR2xp67_ASAP7_75t_L g3883 ( 
.A(n_3778),
.B(n_3309),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3526),
.B(n_3362),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3526),
.B(n_3528),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_3528),
.B(n_3363),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3569),
.Y(n_3887)
);

BUFx6f_ASAP7_75t_L g3888 ( 
.A(n_3719),
.Y(n_3888)
);

AND2x4_ASAP7_75t_L g3889 ( 
.A(n_3395),
.B(n_3031),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3489),
.Y(n_3890)
);

AND3x1_ASAP7_75t_L g3891 ( 
.A(n_3515),
.B(n_980),
.C(n_969),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3576),
.Y(n_3892)
);

INVx3_ASAP7_75t_L g3893 ( 
.A(n_3595),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3585),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3490),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3588),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3609),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3627),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3629),
.Y(n_3899)
);

AOI211xp5_ASAP7_75t_L g3900 ( 
.A1(n_3403),
.A2(n_1212),
.B(n_1042),
.C(n_3291),
.Y(n_3900)
);

INVx2_ASAP7_75t_SL g3901 ( 
.A(n_3719),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3491),
.Y(n_3902)
);

INVx2_ASAP7_75t_SL g3903 ( 
.A(n_3732),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3509),
.Y(n_3904)
);

AND2x4_ASAP7_75t_L g3905 ( 
.A(n_3458),
.B(n_3556),
.Y(n_3905)
);

AOI211xp5_ASAP7_75t_L g3906 ( 
.A1(n_3611),
.A2(n_1042),
.B(n_3295),
.C(n_3333),
.Y(n_3906)
);

INVx1_ASAP7_75t_SL g3907 ( 
.A(n_3522),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_SL g3908 ( 
.A(n_3780),
.B(n_2986),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3511),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3466),
.B(n_3364),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3466),
.B(n_3383),
.Y(n_3911)
);

BUFx2_ASAP7_75t_L g3912 ( 
.A(n_3732),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3583),
.B(n_2940),
.Y(n_3913)
);

HB1xp67_ASAP7_75t_L g3914 ( 
.A(n_3482),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_SL g3915 ( 
.A1(n_3547),
.A2(n_2944),
.B1(n_2940),
.B2(n_3389),
.Y(n_3915)
);

AND2x2_ASAP7_75t_L g3916 ( 
.A(n_3600),
.B(n_3389),
.Y(n_3916)
);

INVx2_ASAP7_75t_L g3917 ( 
.A(n_3514),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3533),
.Y(n_3918)
);

OR2x6_ASAP7_75t_L g3919 ( 
.A(n_3549),
.B(n_3264),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3642),
.Y(n_3920)
);

NOR2xp33_ASAP7_75t_L g3921 ( 
.A(n_3452),
.B(n_3295),
.Y(n_3921)
);

AND3x1_ASAP7_75t_SL g3922 ( 
.A(n_3645),
.B(n_3115),
.C(n_985),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3554),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3583),
.B(n_2944),
.Y(n_3924)
);

INVx3_ASAP7_75t_L g3925 ( 
.A(n_3749),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3646),
.Y(n_3926)
);

BUFx8_ASAP7_75t_SL g3927 ( 
.A(n_3617),
.Y(n_3927)
);

AND2x4_ASAP7_75t_L g3928 ( 
.A(n_3458),
.B(n_3106),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3571),
.Y(n_3929)
);

OAI22xp5_ASAP7_75t_L g3930 ( 
.A1(n_3594),
.A2(n_3318),
.B1(n_3310),
.B2(n_3331),
.Y(n_3930)
);

AOI22xp5_ASAP7_75t_L g3931 ( 
.A1(n_3405),
.A2(n_3295),
.B1(n_3390),
.B2(n_3110),
.Y(n_3931)
);

HB1xp67_ASAP7_75t_L g3932 ( 
.A(n_3550),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3647),
.Y(n_3933)
);

HB1xp67_ASAP7_75t_L g3934 ( 
.A(n_3562),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3648),
.Y(n_3935)
);

INVx2_ASAP7_75t_SL g3936 ( 
.A(n_3439),
.Y(n_3936)
);

CKINVDCx5p33_ASAP7_75t_R g3937 ( 
.A(n_3497),
.Y(n_3937)
);

AOI211xp5_ASAP7_75t_L g3938 ( 
.A1(n_3484),
.A2(n_3333),
.B(n_3369),
.C(n_3366),
.Y(n_3938)
);

AND2x2_ASAP7_75t_SL g3939 ( 
.A(n_3746),
.B(n_3389),
.Y(n_3939)
);

BUFx4f_ASAP7_75t_L g3940 ( 
.A(n_3746),
.Y(n_3940)
);

INVx4_ASAP7_75t_L g3941 ( 
.A(n_3448),
.Y(n_3941)
);

OAI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3442),
.A2(n_3368),
.B1(n_3356),
.B2(n_3351),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3651),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3658),
.Y(n_3944)
);

A2O1A1Ixp33_ASAP7_75t_L g3945 ( 
.A1(n_3791),
.A2(n_3014),
.B(n_3273),
.C(n_3346),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3584),
.B(n_2944),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3584),
.B(n_2944),
.Y(n_3947)
);

BUFx6f_ASAP7_75t_L g3948 ( 
.A(n_3464),
.Y(n_3948)
);

AOI22xp5_ASAP7_75t_SL g3949 ( 
.A1(n_3768),
.A2(n_3298),
.B1(n_3333),
.B2(n_3366),
.Y(n_3949)
);

AND2x2_ASAP7_75t_SL g3950 ( 
.A(n_3731),
.B(n_3369),
.Y(n_3950)
);

HB1xp67_ASAP7_75t_L g3951 ( 
.A(n_3633),
.Y(n_3951)
);

AND2x4_ASAP7_75t_L g3952 ( 
.A(n_3556),
.B(n_3106),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3407),
.B(n_2944),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3483),
.B(n_2944),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3660),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3575),
.Y(n_3956)
);

BUFx12f_ASAP7_75t_L g3957 ( 
.A(n_3696),
.Y(n_3957)
);

INVx4_ASAP7_75t_L g3958 ( 
.A(n_3503),
.Y(n_3958)
);

INVxp67_ASAP7_75t_L g3959 ( 
.A(n_3563),
.Y(n_3959)
);

BUFx4f_ASAP7_75t_L g3960 ( 
.A(n_3430),
.Y(n_3960)
);

INVx4_ASAP7_75t_L g3961 ( 
.A(n_3503),
.Y(n_3961)
);

INVx1_ASAP7_75t_SL g3962 ( 
.A(n_3471),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3577),
.Y(n_3963)
);

BUFx2_ASAP7_75t_SL g3964 ( 
.A(n_3415),
.Y(n_3964)
);

INVxp67_ASAP7_75t_L g3965 ( 
.A(n_3563),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3436),
.B(n_3324),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3436),
.B(n_3324),
.Y(n_3967)
);

AOI22xp5_ASAP7_75t_SL g3968 ( 
.A1(n_3519),
.A2(n_817),
.B1(n_821),
.B2(n_810),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3580),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3433),
.B(n_3324),
.Y(n_3970)
);

AND2x4_ASAP7_75t_L g3971 ( 
.A(n_3722),
.B(n_3106),
.Y(n_3971)
);

AND2x6_ASAP7_75t_L g3972 ( 
.A(n_3722),
.B(n_3470),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3493),
.B(n_3324),
.Y(n_3973)
);

INVx2_ASAP7_75t_SL g3974 ( 
.A(n_3461),
.Y(n_3974)
);

AOI22xp5_ASAP7_75t_L g3975 ( 
.A1(n_3484),
.A2(n_3390),
.B1(n_3014),
.B2(n_2992),
.Y(n_3975)
);

BUFx2_ASAP7_75t_L g3976 ( 
.A(n_3463),
.Y(n_3976)
);

BUFx6f_ASAP7_75t_L g3977 ( 
.A(n_3464),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3502),
.B(n_3324),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3663),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3672),
.Y(n_3980)
);

AOI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_3570),
.A2(n_3390),
.B1(n_2992),
.B2(n_2982),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3674),
.Y(n_3982)
);

AOI22xp33_ASAP7_75t_L g3983 ( 
.A1(n_3589),
.A2(n_3324),
.B1(n_3321),
.B2(n_2992),
.Y(n_3983)
);

INVx3_ASAP7_75t_L g3984 ( 
.A(n_3430),
.Y(n_3984)
);

BUFx2_ASAP7_75t_L g3985 ( 
.A(n_3499),
.Y(n_3985)
);

HB1xp67_ASAP7_75t_L g3986 ( 
.A(n_3635),
.Y(n_3986)
);

BUFx2_ASAP7_75t_L g3987 ( 
.A(n_3396),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3590),
.Y(n_3988)
);

INVxp67_ASAP7_75t_SL g3989 ( 
.A(n_3763),
.Y(n_3989)
);

INVx4_ASAP7_75t_L g3990 ( 
.A(n_3505),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3460),
.B(n_3106),
.Y(n_3991)
);

INVx2_ASAP7_75t_SL g3992 ( 
.A(n_3683),
.Y(n_3992)
);

AND2x4_ASAP7_75t_L g3993 ( 
.A(n_3505),
.B(n_3061),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3605),
.Y(n_3994)
);

INVx2_ASAP7_75t_SL g3995 ( 
.A(n_3692),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3504),
.B(n_3506),
.Y(n_3996)
);

AND2x6_ASAP7_75t_SL g3997 ( 
.A(n_3447),
.B(n_980),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3622),
.Y(n_3998)
);

NOR2xp33_ASAP7_75t_L g3999 ( 
.A(n_3586),
.B(n_3338),
.Y(n_3999)
);

AOI22xp5_ASAP7_75t_L g4000 ( 
.A1(n_3570),
.A2(n_2982),
.B1(n_3340),
.B2(n_3338),
.Y(n_4000)
);

AND2x4_ASAP7_75t_L g4001 ( 
.A(n_3780),
.B(n_3061),
.Y(n_4001)
);

AND2x6_ASAP7_75t_L g4002 ( 
.A(n_3470),
.B(n_3224),
.Y(n_4002)
);

A2O1A1Ixp33_ASAP7_75t_L g4003 ( 
.A1(n_3475),
.A2(n_3273),
.B(n_3349),
.C(n_3346),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3630),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3687),
.Y(n_4005)
);

BUFx3_ASAP7_75t_L g4006 ( 
.A(n_3738),
.Y(n_4006)
);

INVx3_ASAP7_75t_L g4007 ( 
.A(n_3682),
.Y(n_4007)
);

INVx5_ASAP7_75t_L g4008 ( 
.A(n_3690),
.Y(n_4008)
);

HB1xp67_ASAP7_75t_L g4009 ( 
.A(n_3636),
.Y(n_4009)
);

INVx4_ASAP7_75t_L g4010 ( 
.A(n_3682),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3704),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_SL g4012 ( 
.A(n_3671),
.B(n_2986),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3512),
.B(n_3325),
.Y(n_4013)
);

INVx2_ASAP7_75t_SL g4014 ( 
.A(n_3596),
.Y(n_4014)
);

INVx4_ASAP7_75t_L g4015 ( 
.A(n_3464),
.Y(n_4015)
);

AND2x4_ASAP7_75t_L g4016 ( 
.A(n_3410),
.B(n_3129),
.Y(n_4016)
);

AND3x1_ASAP7_75t_SL g4017 ( 
.A(n_3411),
.B(n_989),
.C(n_985),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3706),
.Y(n_4018)
);

CKINVDCx5p33_ASAP7_75t_R g4019 ( 
.A(n_3573),
.Y(n_4019)
);

BUFx6f_ASAP7_75t_L g4020 ( 
.A(n_3464),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3718),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3721),
.Y(n_4022)
);

INVx2_ASAP7_75t_SL g4023 ( 
.A(n_3535),
.Y(n_4023)
);

INVx1_ASAP7_75t_SL g4024 ( 
.A(n_3598),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_L g4025 ( 
.A(n_3513),
.B(n_3325),
.Y(n_4025)
);

INVx3_ASAP7_75t_L g4026 ( 
.A(n_3472),
.Y(n_4026)
);

BUFx6f_ASAP7_75t_L g4027 ( 
.A(n_3481),
.Y(n_4027)
);

INVx2_ASAP7_75t_SL g4028 ( 
.A(n_3665),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3641),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3728),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3734),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_SL g4032 ( 
.A(n_3539),
.B(n_3112),
.Y(n_4032)
);

BUFx6f_ASAP7_75t_L g4033 ( 
.A(n_3481),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3656),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3517),
.B(n_3325),
.Y(n_4035)
);

BUFx6f_ASAP7_75t_L g4036 ( 
.A(n_3481),
.Y(n_4036)
);

OAI22xp33_ASAP7_75t_L g4037 ( 
.A1(n_3404),
.A2(n_3351),
.B1(n_3374),
.B2(n_3183),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_SL g4038 ( 
.A(n_3447),
.B(n_3112),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3736),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3739),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3753),
.B(n_3153),
.Y(n_4041)
);

BUFx2_ASAP7_75t_L g4042 ( 
.A(n_3762),
.Y(n_4042)
);

OAI22xp5_ASAP7_75t_L g4043 ( 
.A1(n_3723),
.A2(n_3183),
.B1(n_3374),
.B2(n_3351),
.Y(n_4043)
);

A2O1A1Ixp33_ASAP7_75t_SL g4044 ( 
.A1(n_3684),
.A2(n_3248),
.B(n_3293),
.C(n_3245),
.Y(n_4044)
);

BUFx2_ASAP7_75t_L g4045 ( 
.A(n_3581),
.Y(n_4045)
);

INVx1_ASAP7_75t_SL g4046 ( 
.A(n_3487),
.Y(n_4046)
);

NOR2x1p5_ASAP7_75t_L g4047 ( 
.A(n_3467),
.B(n_3238),
.Y(n_4047)
);

INVx2_ASAP7_75t_SL g4048 ( 
.A(n_3581),
.Y(n_4048)
);

BUFx3_ASAP7_75t_L g4049 ( 
.A(n_3717),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3758),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3764),
.Y(n_4051)
);

NOR2xp33_ASAP7_75t_L g4052 ( 
.A(n_3760),
.B(n_3338),
.Y(n_4052)
);

INVx2_ASAP7_75t_SL g4053 ( 
.A(n_3603),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3766),
.Y(n_4054)
);

BUFx2_ASAP7_75t_L g4055 ( 
.A(n_3603),
.Y(n_4055)
);

INVx2_ASAP7_75t_L g4056 ( 
.A(n_3657),
.Y(n_4056)
);

BUFx8_ASAP7_75t_L g4057 ( 
.A(n_3761),
.Y(n_4057)
);

OAI22xp5_ASAP7_75t_L g4058 ( 
.A1(n_3726),
.A2(n_3183),
.B1(n_3374),
.B2(n_3351),
.Y(n_4058)
);

CKINVDCx5p33_ASAP7_75t_R g4059 ( 
.A(n_3434),
.Y(n_4059)
);

INVx1_ASAP7_75t_SL g4060 ( 
.A(n_3659),
.Y(n_4060)
);

CKINVDCx8_ASAP7_75t_R g4061 ( 
.A(n_3748),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3770),
.Y(n_4062)
);

HB1xp67_ASAP7_75t_L g4063 ( 
.A(n_3668),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3783),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_SL g4065 ( 
.A(n_3628),
.B(n_3153),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3662),
.Y(n_4066)
);

BUFx6f_ASAP7_75t_L g4067 ( 
.A(n_3481),
.Y(n_4067)
);

NAND2x1p5_ASAP7_75t_L g4068 ( 
.A(n_3472),
.B(n_3152),
.Y(n_4068)
);

BUFx10_ASAP7_75t_L g4069 ( 
.A(n_3510),
.Y(n_4069)
);

HB1xp67_ASAP7_75t_L g4070 ( 
.A(n_3669),
.Y(n_4070)
);

NOR2xp33_ASAP7_75t_L g4071 ( 
.A(n_3760),
.B(n_3340),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3667),
.Y(n_4072)
);

AND2x4_ASAP7_75t_L g4073 ( 
.A(n_3413),
.B(n_3129),
.Y(n_4073)
);

INVx4_ASAP7_75t_L g4074 ( 
.A(n_3555),
.Y(n_4074)
);

INVxp67_ASAP7_75t_L g4075 ( 
.A(n_3510),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3699),
.Y(n_4076)
);

INVx5_ASAP7_75t_L g4077 ( 
.A(n_3690),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3700),
.Y(n_4078)
);

AOI22xp5_ASAP7_75t_L g4079 ( 
.A1(n_3614),
.A2(n_2982),
.B1(n_3340),
.B2(n_3125),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_SL g4080 ( 
.A(n_3628),
.B(n_3182),
.Y(n_4080)
);

AND2x4_ASAP7_75t_L g4081 ( 
.A(n_3419),
.B(n_3131),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3525),
.B(n_3325),
.Y(n_4082)
);

HB1xp67_ASAP7_75t_L g4083 ( 
.A(n_3477),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3531),
.B(n_3325),
.Y(n_4084)
);

HB1xp67_ASAP7_75t_L g4085 ( 
.A(n_3601),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3787),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3714),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3740),
.Y(n_4088)
);

A2O1A1Ixp33_ASAP7_75t_L g4089 ( 
.A1(n_3540),
.A2(n_3349),
.B(n_3316),
.C(n_3327),
.Y(n_4089)
);

INVx3_ASAP7_75t_L g4090 ( 
.A(n_3555),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3705),
.Y(n_4091)
);

NOR2xp33_ASAP7_75t_L g4092 ( 
.A(n_3750),
.B(n_3182),
.Y(n_4092)
);

OR2x6_ASAP7_75t_L g4093 ( 
.A(n_3545),
.B(n_3264),
.Y(n_4093)
);

BUFx6f_ASAP7_75t_L g4094 ( 
.A(n_3555),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3538),
.B(n_3325),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3757),
.Y(n_4096)
);

AND2x4_ASAP7_75t_L g4097 ( 
.A(n_3777),
.B(n_3131),
.Y(n_4097)
);

INVx2_ASAP7_75t_SL g4098 ( 
.A(n_3592),
.Y(n_4098)
);

BUFx3_ASAP7_75t_L g4099 ( 
.A(n_3637),
.Y(n_4099)
);

AOI22xp5_ASAP7_75t_L g4100 ( 
.A1(n_3614),
.A2(n_3690),
.B1(n_3597),
.B2(n_3713),
.Y(n_4100)
);

AND2x4_ASAP7_75t_L g4101 ( 
.A(n_3713),
.B(n_3725),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3707),
.Y(n_4102)
);

NOR2xp33_ASAP7_75t_L g4103 ( 
.A(n_3750),
.B(n_3216),
.Y(n_4103)
);

AOI22xp5_ASAP7_75t_L g4104 ( 
.A1(n_3725),
.A2(n_3125),
.B1(n_3393),
.B2(n_3376),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_3485),
.B(n_1114),
.Y(n_4105)
);

AND2x4_ASAP7_75t_L g4106 ( 
.A(n_3675),
.B(n_3146),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3712),
.Y(n_4107)
);

A2O1A1Ixp33_ASAP7_75t_L g4108 ( 
.A1(n_3638),
.A2(n_3316),
.B(n_3327),
.C(n_3326),
.Y(n_4108)
);

INVxp67_ASAP7_75t_L g4109 ( 
.A(n_3518),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3727),
.Y(n_4110)
);

INVx3_ASAP7_75t_L g4111 ( 
.A(n_3555),
.Y(n_4111)
);

INVx3_ASAP7_75t_L g4112 ( 
.A(n_3602),
.Y(n_4112)
);

INVx5_ASAP7_75t_L g4113 ( 
.A(n_3602),
.Y(n_4113)
);

HAxp5_ASAP7_75t_L g4114 ( 
.A(n_3591),
.B(n_817),
.CON(n_4114),
.SN(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_3741),
.Y(n_4115)
);

INVx4_ASAP7_75t_L g4116 ( 
.A(n_3602),
.Y(n_4116)
);

AOI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_3551),
.A2(n_3393),
.B1(n_3376),
.B2(n_3154),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3638),
.B(n_3655),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_3742),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3655),
.B(n_3385),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3759),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_3765),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3443),
.B(n_3385),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3775),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3737),
.B(n_3744),
.Y(n_4125)
);

BUFx6f_ASAP7_75t_L g4126 ( 
.A(n_3602),
.Y(n_4126)
);

INVxp67_ASAP7_75t_SL g4127 ( 
.A(n_3553),
.Y(n_4127)
);

CKINVDCx5p33_ASAP7_75t_R g4128 ( 
.A(n_3591),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3782),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_3485),
.B(n_1114),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3747),
.B(n_3385),
.Y(n_4131)
);

NOR2xp33_ASAP7_75t_L g4132 ( 
.A(n_3518),
.B(n_3216),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3751),
.B(n_3752),
.Y(n_4133)
);

INVx1_ASAP7_75t_SL g4134 ( 
.A(n_3691),
.Y(n_4134)
);

INVx3_ASAP7_75t_L g4135 ( 
.A(n_3673),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3790),
.Y(n_4136)
);

BUFx4f_ASAP7_75t_L g4137 ( 
.A(n_3673),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3693),
.Y(n_4138)
);

INVx4_ASAP7_75t_L g4139 ( 
.A(n_3673),
.Y(n_4139)
);

AND2x4_ASAP7_75t_L g4140 ( 
.A(n_3675),
.B(n_3146),
.Y(n_4140)
);

INVx2_ASAP7_75t_L g4141 ( 
.A(n_3720),
.Y(n_4141)
);

INVx2_ASAP7_75t_SL g4142 ( 
.A(n_3686),
.Y(n_4142)
);

AND2x2_ASAP7_75t_L g4143 ( 
.A(n_3568),
.B(n_1114),
.Y(n_4143)
);

INVx2_ASAP7_75t_SL g4144 ( 
.A(n_3689),
.Y(n_4144)
);

AND2x4_ASAP7_75t_L g4145 ( 
.A(n_3676),
.B(n_3238),
.Y(n_4145)
);

AOI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_3478),
.A2(n_3385),
.B1(n_3326),
.B2(n_3337),
.Y(n_4146)
);

AO22x1_ASAP7_75t_L g4147 ( 
.A1(n_3441),
.A2(n_3374),
.B1(n_3351),
.B2(n_824),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_3720),
.Y(n_4148)
);

BUFx2_ASAP7_75t_L g4149 ( 
.A(n_3673),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_3755),
.B(n_3756),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3694),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_SL g4152 ( 
.A(n_3478),
.B(n_3238),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_3568),
.B(n_1124),
.Y(n_4153)
);

INVx2_ASAP7_75t_L g4154 ( 
.A(n_3735),
.Y(n_4154)
);

INVx1_ASAP7_75t_SL g4155 ( 
.A(n_3695),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_3735),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_3769),
.B(n_3385),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_SL g4158 ( 
.A(n_3684),
.B(n_3374),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3698),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3771),
.B(n_3385),
.Y(n_4160)
);

AND2x4_ASAP7_75t_L g4161 ( 
.A(n_3676),
.B(n_2948),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_3681),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_3685),
.Y(n_4163)
);

AOI22xp33_ASAP7_75t_L g4164 ( 
.A1(n_3661),
.A2(n_2916),
.B1(n_2917),
.B2(n_2903),
.Y(n_4164)
);

AOI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3661),
.A2(n_2916),
.B1(n_2917),
.B2(n_2903),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3701),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3708),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_3709),
.Y(n_4168)
);

AND2x6_ASAP7_75t_L g4169 ( 
.A(n_3796),
.B(n_3823),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3822),
.B(n_3626),
.Y(n_4170)
);

HB1xp67_ASAP7_75t_L g4171 ( 
.A(n_3795),
.Y(n_4171)
);

OAI22xp5_ASAP7_75t_SL g4172 ( 
.A1(n_4019),
.A2(n_3670),
.B1(n_3523),
.B2(n_3664),
.Y(n_4172)
);

INVxp67_ASAP7_75t_L g4173 ( 
.A(n_3987),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3799),
.Y(n_4174)
);

NAND2x1p5_ASAP7_75t_L g4175 ( 
.A(n_3832),
.B(n_3960),
.Y(n_4175)
);

AOI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_4127),
.A2(n_3623),
.B(n_3553),
.Y(n_4176)
);

AOI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_4127),
.A2(n_3619),
.B(n_3416),
.Y(n_4177)
);

AOI22xp5_ASAP7_75t_L g4178 ( 
.A1(n_3900),
.A2(n_3733),
.B1(n_3644),
.B2(n_3786),
.Y(n_4178)
);

AOI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_3989),
.A2(n_3560),
.B(n_3401),
.Y(n_4179)
);

O2A1O1Ixp33_ASAP7_75t_L g4180 ( 
.A1(n_3860),
.A2(n_3593),
.B(n_3560),
.C(n_3639),
.Y(n_4180)
);

OAI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_3989),
.A2(n_3784),
.B1(n_3789),
.B2(n_3767),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_4046),
.B(n_3666),
.Y(n_4182)
);

NOR2xp33_ASAP7_75t_L g4183 ( 
.A(n_3882),
.B(n_3907),
.Y(n_4183)
);

OAI22xp5_ASAP7_75t_SL g4184 ( 
.A1(n_3869),
.A2(n_3664),
.B1(n_3666),
.B2(n_3731),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_R g4185 ( 
.A(n_3833),
.B(n_3574),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3802),
.Y(n_4186)
);

AOI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_4043),
.A2(n_3606),
.B(n_3604),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_4046),
.B(n_3710),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_3797),
.Y(n_4189)
);

AOI21xp5_ASAP7_75t_L g4190 ( 
.A1(n_4043),
.A2(n_3639),
.B(n_3462),
.Y(n_4190)
);

OAI22xp5_ASAP7_75t_L g4191 ( 
.A1(n_3885),
.A2(n_3784),
.B1(n_3789),
.B2(n_3767),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3806),
.Y(n_4192)
);

BUFx6f_ASAP7_75t_L g4193 ( 
.A(n_3801),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_3907),
.B(n_3631),
.Y(n_4194)
);

O2A1O1Ixp33_ASAP7_75t_L g4195 ( 
.A1(n_3945),
.A2(n_3593),
.B(n_3501),
.C(n_3716),
.Y(n_4195)
);

BUFx6f_ASAP7_75t_L g4196 ( 
.A(n_3801),
.Y(n_4196)
);

AOI21xp5_ASAP7_75t_L g4197 ( 
.A1(n_4058),
.A2(n_3702),
.B(n_3745),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_3882),
.B(n_3664),
.Y(n_4198)
);

NOR3xp33_ASAP7_75t_L g4199 ( 
.A(n_4038),
.B(n_3453),
.C(n_992),
.Y(n_4199)
);

INVx5_ASAP7_75t_L g4200 ( 
.A(n_3919),
.Y(n_4200)
);

BUFx6f_ASAP7_75t_L g4201 ( 
.A(n_3801),
.Y(n_4201)
);

O2A1O1Ixp33_ASAP7_75t_L g4202 ( 
.A1(n_4089),
.A2(n_3716),
.B(n_3424),
.C(n_3417),
.Y(n_4202)
);

BUFx3_ASAP7_75t_L g4203 ( 
.A(n_3807),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3822),
.B(n_3626),
.Y(n_4204)
);

NOR3xp33_ASAP7_75t_L g4205 ( 
.A(n_4147),
.B(n_992),
.C(n_989),
.Y(n_4205)
);

INVx3_ASAP7_75t_L g4206 ( 
.A(n_3803),
.Y(n_4206)
);

INVx2_ASAP7_75t_SL g4207 ( 
.A(n_3827),
.Y(n_4207)
);

O2A1O1Ixp33_ASAP7_75t_SL g4208 ( 
.A1(n_4118),
.A2(n_3703),
.B(n_3697),
.C(n_3625),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_SL g4209 ( 
.A(n_3812),
.B(n_3697),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4024),
.B(n_3650),
.Y(n_4210)
);

BUFx6f_ASAP7_75t_L g4211 ( 
.A(n_3803),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_L g4212 ( 
.A(n_3811),
.B(n_3703),
.Y(n_4212)
);

AOI21xp5_ASAP7_75t_L g4213 ( 
.A1(n_4058),
.A2(n_3930),
.B(n_3996),
.Y(n_4213)
);

BUFx2_ASAP7_75t_L g4214 ( 
.A(n_3855),
.Y(n_4214)
);

NOR2xp33_ASAP7_75t_L g4215 ( 
.A(n_4128),
.B(n_3435),
.Y(n_4215)
);

NOR2xp33_ASAP7_75t_L g4216 ( 
.A(n_3847),
.B(n_3677),
.Y(n_4216)
);

NOR2x1_ASAP7_75t_L g4217 ( 
.A(n_3825),
.B(n_3724),
.Y(n_4217)
);

OAI22xp5_ASAP7_75t_L g4218 ( 
.A1(n_3885),
.A2(n_3776),
.B1(n_3781),
.B2(n_3773),
.Y(n_4218)
);

OAI22xp5_ASAP7_75t_L g4219 ( 
.A1(n_4118),
.A2(n_4125),
.B1(n_4150),
.B2(n_4133),
.Y(n_4219)
);

BUFx2_ASAP7_75t_L g4220 ( 
.A(n_3912),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_3792),
.B(n_3650),
.Y(n_4221)
);

OAI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_4125),
.A2(n_3654),
.B1(n_3612),
.B2(n_3613),
.Y(n_4222)
);

A2O1A1Ixp33_ASAP7_75t_L g4223 ( 
.A1(n_3869),
.A2(n_3544),
.B(n_3634),
.C(n_3654),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_3834),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3836),
.Y(n_4225)
);

OA22x2_ASAP7_75t_L g4226 ( 
.A1(n_3831),
.A2(n_3621),
.B1(n_3640),
.B2(n_3496),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4024),
.B(n_3607),
.Y(n_4227)
);

NAND3xp33_ASAP7_75t_SL g4228 ( 
.A(n_3938),
.B(n_3906),
.C(n_3798),
.Y(n_4228)
);

HB1xp67_ASAP7_75t_L g4229 ( 
.A(n_3795),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3804),
.Y(n_4230)
);

A2O1A1Ixp33_ASAP7_75t_L g4231 ( 
.A1(n_4117),
.A2(n_3772),
.B(n_3451),
.C(n_3457),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_SL g4232 ( 
.A(n_3853),
.B(n_3561),
.Y(n_4232)
);

BUFx2_ASAP7_75t_L g4233 ( 
.A(n_3835),
.Y(n_4233)
);

O2A1O1Ixp33_ASAP7_75t_L g4234 ( 
.A1(n_3930),
.A2(n_993),
.B(n_999),
.C(n_998),
.Y(n_4234)
);

OR2x6_ASAP7_75t_L g4235 ( 
.A(n_3919),
.B(n_3264),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_3870),
.B(n_1124),
.Y(n_4236)
);

A2O1A1Ixp33_ASAP7_75t_L g4237 ( 
.A1(n_3975),
.A2(n_3983),
.B(n_4130),
.C(n_4105),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3808),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3818),
.B(n_3615),
.Y(n_4239)
);

NAND3xp33_ASAP7_75t_L g4240 ( 
.A(n_3983),
.B(n_998),
.C(n_993),
.Y(n_4240)
);

AO21x1_ASAP7_75t_L g4241 ( 
.A1(n_3942),
.A2(n_3546),
.B(n_3520),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_3996),
.A2(n_4150),
.B(n_4133),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_3818),
.B(n_3616),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_3843),
.B(n_3677),
.Y(n_4244)
);

BUFx2_ASAP7_75t_SL g4245 ( 
.A(n_3883),
.Y(n_4245)
);

AND2x4_ASAP7_75t_L g4246 ( 
.A(n_3796),
.B(n_3971),
.Y(n_4246)
);

INVx2_ASAP7_75t_SL g4247 ( 
.A(n_3846),
.Y(n_4247)
);

OAI22xp5_ASAP7_75t_SL g4248 ( 
.A1(n_3891),
.A2(n_3937),
.B1(n_3957),
.B2(n_3820),
.Y(n_4248)
);

AOI22xp33_ASAP7_75t_SL g4249 ( 
.A1(n_3849),
.A2(n_3450),
.B1(n_1190),
.B2(n_1246),
.Y(n_4249)
);

NOR2xp33_ASAP7_75t_R g4250 ( 
.A(n_3936),
.B(n_3793),
.Y(n_4250)
);

OAI21xp5_ASAP7_75t_L g4251 ( 
.A1(n_4108),
.A2(n_3572),
.B(n_3474),
.Y(n_4251)
);

AOI21xp5_ASAP7_75t_L g4252 ( 
.A1(n_4037),
.A2(n_3649),
.B(n_3520),
.Y(n_4252)
);

AO21x1_ASAP7_75t_L g4253 ( 
.A1(n_3942),
.A2(n_3532),
.B(n_3508),
.Y(n_4253)
);

INVx4_ASAP7_75t_L g4254 ( 
.A(n_4137),
.Y(n_4254)
);

AOI33xp33_ASAP7_75t_L g4255 ( 
.A1(n_3809),
.A2(n_1021),
.A3(n_1007),
.B1(n_1024),
.B2(n_1018),
.B3(n_999),
.Y(n_4255)
);

AOI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_4037),
.A2(n_3532),
.B(n_3508),
.Y(n_4256)
);

BUFx6f_ASAP7_75t_L g4257 ( 
.A(n_3803),
.Y(n_4257)
);

BUFx3_ASAP7_75t_L g4258 ( 
.A(n_3852),
.Y(n_4258)
);

BUFx6f_ASAP7_75t_L g4259 ( 
.A(n_3814),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3810),
.Y(n_4260)
);

NOR2xp33_ASAP7_75t_L g4261 ( 
.A(n_4075),
.B(n_821),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3843),
.B(n_2922),
.Y(n_4262)
);

O2A1O1Ixp33_ASAP7_75t_L g4263 ( 
.A1(n_4003),
.A2(n_1007),
.B(n_1021),
.C(n_1018),
.Y(n_4263)
);

NOR2xp33_ASAP7_75t_L g4264 ( 
.A(n_4075),
.B(n_824),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_3850),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_4131),
.A2(n_3543),
.B(n_3542),
.Y(n_4266)
);

O2A1O1Ixp33_ASAP7_75t_SL g4267 ( 
.A1(n_4044),
.A2(n_3498),
.B(n_3543),
.C(n_3542),
.Y(n_4267)
);

CKINVDCx20_ASAP7_75t_R g4268 ( 
.A(n_3815),
.Y(n_4268)
);

NOR2xp33_ASAP7_75t_L g4269 ( 
.A(n_4109),
.B(n_3997),
.Y(n_4269)
);

OAI22xp5_ASAP7_75t_L g4270 ( 
.A1(n_4146),
.A2(n_2926),
.B1(n_2922),
.B2(n_1025),
.Y(n_4270)
);

AOI21xp5_ASAP7_75t_L g4271 ( 
.A1(n_4131),
.A2(n_4160),
.B(n_4157),
.Y(n_4271)
);

A2O1A1Ixp33_ASAP7_75t_L g4272 ( 
.A1(n_4143),
.A2(n_3337),
.B(n_3730),
.C(n_3624),
.Y(n_4272)
);

INVx1_ASAP7_75t_SL g4273 ( 
.A(n_3805),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_3879),
.Y(n_4274)
);

OR2x2_ASAP7_75t_L g4275 ( 
.A(n_3874),
.B(n_3162),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3813),
.Y(n_4276)
);

INVx3_ASAP7_75t_L g4277 ( 
.A(n_3814),
.Y(n_4277)
);

CKINVDCx10_ASAP7_75t_R g4278 ( 
.A(n_3875),
.Y(n_4278)
);

NOR2xp33_ASAP7_75t_L g4279 ( 
.A(n_4109),
.B(n_825),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_4060),
.B(n_4087),
.Y(n_4280)
);

AOI21xp5_ASAP7_75t_L g4281 ( 
.A1(n_4157),
.A2(n_3624),
.B(n_3582),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_3817),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_3921),
.B(n_1124),
.Y(n_4283)
);

BUFx4f_ASAP7_75t_L g4284 ( 
.A(n_3814),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_3880),
.Y(n_4285)
);

AOI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4160),
.A2(n_3679),
.B(n_3582),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4060),
.B(n_2926),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_SL g4288 ( 
.A(n_3841),
.B(n_3561),
.Y(n_4288)
);

INVx1_ASAP7_75t_SL g4289 ( 
.A(n_3805),
.Y(n_4289)
);

A2O1A1Ixp33_ASAP7_75t_SL g4290 ( 
.A1(n_4007),
.A2(n_1025),
.B(n_1026),
.C(n_1024),
.Y(n_4290)
);

BUFx2_ASAP7_75t_L g4291 ( 
.A(n_3846),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_3829),
.B(n_1124),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_3819),
.Y(n_4293)
);

INVx1_ASAP7_75t_SL g4294 ( 
.A(n_4045),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_3890),
.Y(n_4295)
);

AOI21x1_ASAP7_75t_L g4296 ( 
.A1(n_4041),
.A2(n_3688),
.B(n_3679),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_L g4297 ( 
.A(n_3999),
.B(n_825),
.Y(n_4297)
);

AND2x4_ASAP7_75t_L g4298 ( 
.A(n_3971),
.B(n_3928),
.Y(n_4298)
);

AOI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_4013),
.A2(n_3754),
.B(n_3688),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_4088),
.B(n_3114),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_3895),
.Y(n_4301)
);

AOI22xp5_ASAP7_75t_L g4302 ( 
.A1(n_3931),
.A2(n_3845),
.B1(n_3794),
.B2(n_3922),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_3816),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4096),
.B(n_3128),
.Y(n_4304)
);

INVxp67_ASAP7_75t_L g4305 ( 
.A(n_3976),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_4134),
.B(n_3162),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_4134),
.B(n_2957),
.Y(n_4307)
);

BUFx2_ASAP7_75t_L g4308 ( 
.A(n_3846),
.Y(n_4308)
);

AOI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_4013),
.A2(n_4035),
.B(n_4025),
.Y(n_4309)
);

AOI21x1_ASAP7_75t_L g4310 ( 
.A1(n_4158),
.A2(n_3774),
.B(n_3754),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_L g4311 ( 
.A(n_4049),
.B(n_827),
.Y(n_4311)
);

A2O1A1Ixp33_ASAP7_75t_L g4312 ( 
.A1(n_4153),
.A2(n_3940),
.B(n_3823),
.C(n_3954),
.Y(n_4312)
);

O2A1O1Ixp33_ASAP7_75t_L g4313 ( 
.A1(n_3842),
.A2(n_1026),
.B(n_1032),
.C(n_1028),
.Y(n_4313)
);

O2A1O1Ixp33_ASAP7_75t_L g4314 ( 
.A1(n_4114),
.A2(n_1028),
.B(n_1041),
.C(n_1032),
.Y(n_4314)
);

NOR2xp33_ASAP7_75t_L g4315 ( 
.A(n_4101),
.B(n_3820),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3821),
.Y(n_4316)
);

AO32x1_ASAP7_75t_L g4317 ( 
.A1(n_4142),
.A2(n_3159),
.A3(n_3339),
.B1(n_3380),
.B2(n_3290),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_3902),
.Y(n_4318)
);

AOI21xp5_ASAP7_75t_L g4319 ( 
.A1(n_4025),
.A2(n_3785),
.B(n_3774),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_SL g4320 ( 
.A(n_3940),
.B(n_2964),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4155),
.B(n_2961),
.Y(n_4321)
);

O2A1O1Ixp33_ASAP7_75t_L g4322 ( 
.A1(n_3867),
.A2(n_1041),
.B(n_1046),
.C(n_1045),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_3824),
.Y(n_4323)
);

AOI21xp5_ASAP7_75t_L g4324 ( 
.A1(n_4035),
.A2(n_3785),
.B(n_3618),
.Y(n_4324)
);

OAI22xp5_ASAP7_75t_L g4325 ( 
.A1(n_3910),
.A2(n_1046),
.B1(n_1047),
.B2(n_1045),
.Y(n_4325)
);

BUFx2_ASAP7_75t_L g4326 ( 
.A(n_3888),
.Y(n_4326)
);

OAI22xp5_ASAP7_75t_L g4327 ( 
.A1(n_3910),
.A2(n_1054),
.B1(n_1057),
.B2(n_1047),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4155),
.B(n_3932),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_3932),
.B(n_3173),
.Y(n_4329)
);

OAI21x1_ASAP7_75t_L g4330 ( 
.A1(n_3865),
.A2(n_3788),
.B(n_3618),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_3904),
.Y(n_4331)
);

OAI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_3911),
.A2(n_1057),
.B1(n_1061),
.B2(n_1054),
.Y(n_4332)
);

A2O1A1Ixp33_ASAP7_75t_L g4333 ( 
.A1(n_3954),
.A2(n_2956),
.B(n_3044),
.C(n_2993),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_SL g4334 ( 
.A(n_4100),
.B(n_2964),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_3909),
.Y(n_4335)
);

INVx4_ASAP7_75t_L g4336 ( 
.A(n_4137),
.Y(n_4336)
);

CKINVDCx16_ASAP7_75t_R g4337 ( 
.A(n_4042),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_SL g4338 ( 
.A(n_3959),
.B(n_2964),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_4082),
.A2(n_3678),
.B(n_3557),
.Y(n_4339)
);

NOR2xp33_ASAP7_75t_L g4340 ( 
.A(n_4101),
.B(n_827),
.Y(n_4340)
);

OAI22xp5_ASAP7_75t_L g4341 ( 
.A1(n_3911),
.A2(n_1065),
.B1(n_1066),
.B2(n_1061),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_3934),
.B(n_2961),
.Y(n_4342)
);

A2O1A1Ixp33_ASAP7_75t_L g4343 ( 
.A1(n_3848),
.A2(n_2956),
.B(n_3044),
.C(n_2959),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_3828),
.Y(n_4344)
);

NOR2xp33_ASAP7_75t_L g4345 ( 
.A(n_3985),
.B(n_830),
.Y(n_4345)
);

A2O1A1Ixp33_ASAP7_75t_L g4346 ( 
.A1(n_3848),
.A2(n_2959),
.B(n_3122),
.C(n_2993),
.Y(n_4346)
);

O2A1O1Ixp33_ASAP7_75t_L g4347 ( 
.A1(n_3959),
.A2(n_3965),
.B(n_4152),
.C(n_3838),
.Y(n_4347)
);

CKINVDCx5p33_ASAP7_75t_R g4348 ( 
.A(n_3974),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_SL g4349 ( 
.A(n_3965),
.B(n_3857),
.Y(n_4349)
);

AOI21xp5_ASAP7_75t_L g4350 ( 
.A1(n_4082),
.A2(n_3678),
.B(n_3557),
.Y(n_4350)
);

BUFx2_ASAP7_75t_L g4351 ( 
.A(n_3888),
.Y(n_4351)
);

AOI21x1_ASAP7_75t_L g4352 ( 
.A1(n_4065),
.A2(n_3425),
.B(n_3421),
.Y(n_4352)
);

INVx3_ASAP7_75t_L g4353 ( 
.A(n_3816),
.Y(n_4353)
);

INVx3_ASAP7_75t_L g4354 ( 
.A(n_3816),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_3934),
.B(n_3233),
.Y(n_4355)
);

AOI21xp5_ASAP7_75t_L g4356 ( 
.A1(n_4084),
.A2(n_3743),
.B(n_3715),
.Y(n_4356)
);

OR2x2_ASAP7_75t_L g4357 ( 
.A(n_3874),
.B(n_1350),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_3916),
.B(n_1124),
.Y(n_4358)
);

NAND2x1p5_ASAP7_75t_L g4359 ( 
.A(n_3832),
.B(n_3456),
.Y(n_4359)
);

AOI21xp5_ASAP7_75t_L g4360 ( 
.A1(n_4084),
.A2(n_3743),
.B(n_3715),
.Y(n_4360)
);

AND2x4_ASAP7_75t_L g4361 ( 
.A(n_3928),
.B(n_3456),
.Y(n_4361)
);

OAI22xp5_ASAP7_75t_L g4362 ( 
.A1(n_3884),
.A2(n_1066),
.B1(n_1085),
.B2(n_1065),
.Y(n_4362)
);

OAI22xp5_ASAP7_75t_L g4363 ( 
.A1(n_3884),
.A2(n_1087),
.B1(n_1090),
.B2(n_1085),
.Y(n_4363)
);

OAI21xp33_ASAP7_75t_L g4364 ( 
.A1(n_3886),
.A2(n_1243),
.B(n_833),
.Y(n_4364)
);

AOI21x1_ASAP7_75t_L g4365 ( 
.A1(n_4080),
.A2(n_3425),
.B(n_3421),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_3886),
.B(n_2951),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_3951),
.B(n_2951),
.Y(n_4367)
);

BUFx12f_ASAP7_75t_L g4368 ( 
.A(n_3825),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3839),
.Y(n_4369)
);

BUFx2_ASAP7_75t_L g4370 ( 
.A(n_3888),
.Y(n_4370)
);

OAI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_3966),
.A2(n_1090),
.B1(n_1098),
.B2(n_1087),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_SL g4372 ( 
.A(n_3857),
.B(n_2966),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_3840),
.Y(n_4373)
);

INVx2_ASAP7_75t_L g4374 ( 
.A(n_3917),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_3951),
.B(n_3173),
.Y(n_4375)
);

BUFx2_ASAP7_75t_L g4376 ( 
.A(n_3901),
.Y(n_4376)
);

AOI21xp5_ASAP7_75t_L g4377 ( 
.A1(n_4095),
.A2(n_3978),
.B(n_3973),
.Y(n_4377)
);

O2A1O1Ixp33_ASAP7_75t_L g4378 ( 
.A1(n_4012),
.A2(n_1098),
.B(n_1102),
.C(n_1099),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_3918),
.Y(n_4379)
);

AOI21xp5_ASAP7_75t_L g4380 ( 
.A1(n_4095),
.A2(n_3445),
.B(n_3468),
.Y(n_4380)
);

AOI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_3973),
.A2(n_3445),
.B(n_3468),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_3844),
.Y(n_4382)
);

BUFx3_ASAP7_75t_L g4383 ( 
.A(n_4006),
.Y(n_4383)
);

AND2x4_ASAP7_75t_L g4384 ( 
.A(n_3952),
.B(n_3889),
.Y(n_4384)
);

A2O1A1Ixp33_ASAP7_75t_L g4385 ( 
.A1(n_3913),
.A2(n_3103),
.B(n_3123),
.C(n_3122),
.Y(n_4385)
);

CKINVDCx8_ASAP7_75t_R g4386 ( 
.A(n_3964),
.Y(n_4386)
);

BUFx6f_ASAP7_75t_L g4387 ( 
.A(n_3832),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_SL g4388 ( 
.A(n_3857),
.B(n_2966),
.Y(n_4388)
);

BUFx6f_ASAP7_75t_L g4389 ( 
.A(n_3832),
.Y(n_4389)
);

AOI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_3978),
.A2(n_4123),
.B(n_4120),
.Y(n_4390)
);

INVx1_ASAP7_75t_SL g4391 ( 
.A(n_4055),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_3986),
.B(n_3128),
.Y(n_4392)
);

AOI22xp33_ASAP7_75t_L g4393 ( 
.A1(n_3950),
.A2(n_3142),
.B1(n_3151),
.B2(n_3136),
.Y(n_4393)
);

BUFx3_ASAP7_75t_L g4394 ( 
.A(n_4014),
.Y(n_4394)
);

AOI21xp5_ASAP7_75t_L g4395 ( 
.A1(n_4123),
.A2(n_4120),
.B(n_3970),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_3851),
.Y(n_4396)
);

O2A1O1Ixp5_ASAP7_75t_SL g4397 ( 
.A1(n_3861),
.A2(n_1356),
.B(n_1357),
.C(n_1352),
.Y(n_4397)
);

OAI22xp5_ASAP7_75t_L g4398 ( 
.A1(n_3966),
.A2(n_1102),
.B1(n_1104),
.B2(n_1099),
.Y(n_4398)
);

AOI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_3970),
.A2(n_3507),
.B(n_3500),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_SL g4400 ( 
.A(n_3857),
.B(n_2966),
.Y(n_4400)
);

AOI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_3800),
.A2(n_3507),
.B(n_3500),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_3862),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_3866),
.Y(n_4403)
);

O2A1O1Ixp33_ASAP7_75t_SL g4404 ( 
.A1(n_3913),
.A2(n_3123),
.B(n_3103),
.C(n_3271),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_3923),
.Y(n_4405)
);

OAI22xp5_ASAP7_75t_SL g4406 ( 
.A1(n_4061),
.A2(n_833),
.B1(n_834),
.B2(n_830),
.Y(n_4406)
);

O2A1O1Ixp33_ASAP7_75t_L g4407 ( 
.A1(n_3924),
.A2(n_1109),
.B(n_1112),
.C(n_1104),
.Y(n_4407)
);

INVx3_ASAP7_75t_L g4408 ( 
.A(n_3960),
.Y(n_4408)
);

BUFx2_ASAP7_75t_L g4409 ( 
.A(n_3903),
.Y(n_4409)
);

O2A1O1Ixp33_ASAP7_75t_SL g4410 ( 
.A1(n_3924),
.A2(n_3312),
.B(n_3328),
.C(n_3271),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_3929),
.Y(n_4411)
);

AOI22xp5_ASAP7_75t_L g4412 ( 
.A1(n_3922),
.A2(n_3981),
.B1(n_4000),
.B2(n_4028),
.Y(n_4412)
);

O2A1O1Ixp33_ASAP7_75t_L g4413 ( 
.A1(n_3946),
.A2(n_1112),
.B(n_1118),
.C(n_1109),
.Y(n_4413)
);

AOI21xp5_ASAP7_75t_L g4414 ( 
.A1(n_3800),
.A2(n_2960),
.B(n_2937),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_3986),
.B(n_3136),
.Y(n_4415)
);

HB1xp67_ASAP7_75t_L g4416 ( 
.A(n_4009),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_4009),
.B(n_3142),
.Y(n_4417)
);

AND2x4_ASAP7_75t_L g4418 ( 
.A(n_3952),
.B(n_3245),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_3956),
.Y(n_4419)
);

A2O1A1Ixp33_ASAP7_75t_L g4420 ( 
.A1(n_3946),
.A2(n_3494),
.B(n_2620),
.C(n_3156),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_3963),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_SL g4422 ( 
.A(n_3864),
.B(n_2966),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_3871),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_SL g4424 ( 
.A(n_3864),
.B(n_2971),
.Y(n_4424)
);

O2A1O1Ixp5_ASAP7_75t_SL g4425 ( 
.A1(n_3872),
.A2(n_1356),
.B(n_1357),
.C(n_1352),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_3854),
.A2(n_2960),
.B(n_2937),
.Y(n_4426)
);

CKINVDCx20_ASAP7_75t_R g4427 ( 
.A(n_4057),
.Y(n_4427)
);

AOI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_3947),
.A2(n_2960),
.B(n_2937),
.Y(n_4428)
);

A2O1A1Ixp33_ASAP7_75t_L g4429 ( 
.A1(n_3947),
.A2(n_2925),
.B(n_2924),
.C(n_1132),
.Y(n_4429)
);

BUFx8_ASAP7_75t_L g4430 ( 
.A(n_4098),
.Y(n_4430)
);

A2O1A1Ixp33_ASAP7_75t_L g4431 ( 
.A1(n_3967),
.A2(n_3949),
.B(n_3865),
.C(n_3858),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_SL g4432 ( 
.A(n_3864),
.B(n_2971),
.Y(n_4432)
);

OAI22xp5_ASAP7_75t_L g4433 ( 
.A1(n_3967),
.A2(n_1132),
.B1(n_1133),
.B2(n_1118),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_SL g4434 ( 
.A(n_3864),
.B(n_2971),
.Y(n_4434)
);

NOR2x1p5_ASAP7_75t_SL g4435 ( 
.A(n_3873),
.B(n_2824),
.Y(n_4435)
);

O2A1O1Ixp33_ASAP7_75t_L g4436 ( 
.A1(n_4032),
.A2(n_1136),
.B(n_1144),
.C(n_1133),
.Y(n_4436)
);

INVx3_ASAP7_75t_L g4437 ( 
.A(n_3972),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_3876),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_3881),
.Y(n_4439)
);

AOI21xp5_ASAP7_75t_L g4440 ( 
.A1(n_3858),
.A2(n_4077),
.B(n_4008),
.Y(n_4440)
);

NOR2xp33_ASAP7_75t_L g4441 ( 
.A(n_4069),
.B(n_834),
.Y(n_4441)
);

BUFx2_ASAP7_75t_L g4442 ( 
.A(n_3972),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4063),
.B(n_3151),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_3969),
.Y(n_4444)
);

INVxp67_ASAP7_75t_L g4445 ( 
.A(n_4023),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_SL g4446 ( 
.A(n_4008),
.B(n_2971),
.Y(n_4446)
);

INVx4_ASAP7_75t_L g4447 ( 
.A(n_4113),
.Y(n_4447)
);

AOI21xp5_ASAP7_75t_L g4448 ( 
.A1(n_4008),
.A2(n_2979),
.B(n_2962),
.Y(n_4448)
);

OR2x6_ASAP7_75t_L g4449 ( 
.A(n_3919),
.B(n_2995),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_3988),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_3887),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4063),
.B(n_3179),
.Y(n_4452)
);

BUFx6f_ASAP7_75t_L g4453 ( 
.A(n_3889),
.Y(n_4453)
);

BUFx12f_ASAP7_75t_L g4454 ( 
.A(n_3837),
.Y(n_4454)
);

INVxp67_ASAP7_75t_SL g4455 ( 
.A(n_4070),
.Y(n_4455)
);

NOR2xp33_ASAP7_75t_L g4456 ( 
.A(n_4069),
.B(n_965),
.Y(n_4456)
);

OAI21xp5_ASAP7_75t_L g4457 ( 
.A1(n_3953),
.A2(n_3328),
.B(n_3312),
.Y(n_4457)
);

AOI22x1_ASAP7_75t_L g4458 ( 
.A1(n_3830),
.A2(n_1111),
.B1(n_1113),
.B2(n_965),
.Y(n_4458)
);

AND2x4_ASAP7_75t_L g4459 ( 
.A(n_3863),
.B(n_3925),
.Y(n_4459)
);

INVx2_ASAP7_75t_L g4460 ( 
.A(n_3994),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_SL g4461 ( 
.A(n_4008),
.B(n_2976),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_3892),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_4070),
.B(n_3179),
.Y(n_4463)
);

NOR3xp33_ASAP7_75t_SL g4464 ( 
.A(n_4092),
.B(n_1113),
.C(n_1111),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_3894),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_3896),
.Y(n_4466)
);

CKINVDCx8_ASAP7_75t_R g4467 ( 
.A(n_4059),
.Y(n_4467)
);

NOR2xp33_ASAP7_75t_L g4468 ( 
.A(n_4106),
.B(n_1116),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_4138),
.B(n_3181),
.Y(n_4469)
);

AOI22xp5_ASAP7_75t_L g4470 ( 
.A1(n_4052),
.A2(n_1190),
.B1(n_1246),
.B2(n_1241),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4151),
.B(n_3181),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4159),
.B(n_3184),
.Y(n_4472)
);

AOI21xp5_ASAP7_75t_L g4473 ( 
.A1(n_4077),
.A2(n_2979),
.B(n_2962),
.Y(n_4473)
);

A2O1A1Ixp33_ASAP7_75t_L g4474 ( 
.A1(n_3953),
.A2(n_4132),
.B(n_4079),
.C(n_4104),
.Y(n_4474)
);

BUFx2_ASAP7_75t_L g4475 ( 
.A(n_3972),
.Y(n_4475)
);

BUFx12f_ASAP7_75t_L g4476 ( 
.A(n_3837),
.Y(n_4476)
);

A2O1A1Ixp33_ASAP7_75t_L g4477 ( 
.A1(n_3915),
.A2(n_4166),
.B(n_4168),
.C(n_4167),
.Y(n_4477)
);

AOI22xp33_ASAP7_75t_L g4478 ( 
.A1(n_3915),
.A2(n_3387),
.B1(n_3392),
.B2(n_3382),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_3856),
.B(n_3184),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_3968),
.B(n_1190),
.Y(n_4480)
);

OAI22xp5_ASAP7_75t_SL g4481 ( 
.A1(n_4077),
.A2(n_1241),
.B1(n_1242),
.B2(n_1116),
.Y(n_4481)
);

OAI21xp33_ASAP7_75t_SL g4482 ( 
.A1(n_4026),
.A2(n_3248),
.B(n_3245),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_SL g4483 ( 
.A(n_4077),
.B(n_2976),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_3856),
.B(n_3204),
.Y(n_4484)
);

NOR2xp33_ASAP7_75t_L g4485 ( 
.A(n_4106),
.B(n_1242),
.Y(n_4485)
);

OAI21x1_ASAP7_75t_L g4486 ( 
.A1(n_4090),
.A2(n_3067),
.B(n_3608),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_3914),
.B(n_3204),
.Y(n_4487)
);

A2O1A1Ixp33_ASAP7_75t_L g4488 ( 
.A1(n_4071),
.A2(n_2925),
.B(n_2924),
.C(n_1144),
.Y(n_4488)
);

BUFx4f_ASAP7_75t_SL g4489 ( 
.A(n_4057),
.Y(n_4489)
);

AO32x2_ASAP7_75t_L g4490 ( 
.A1(n_4144),
.A2(n_2679),
.A3(n_3315),
.B1(n_3284),
.B2(n_3274),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_3998),
.Y(n_4491)
);

AO32x2_ASAP7_75t_L g4492 ( 
.A1(n_4048),
.A2(n_2679),
.A3(n_3315),
.B1(n_3284),
.B2(n_3274),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_3905),
.B(n_1190),
.Y(n_4493)
);

AOI22xp5_ASAP7_75t_L g4494 ( 
.A1(n_3939),
.A2(n_1246),
.B1(n_1190),
.B2(n_1244),
.Y(n_4494)
);

INVx2_ASAP7_75t_SL g4495 ( 
.A(n_3992),
.Y(n_4495)
);

AOI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_4093),
.A2(n_2979),
.B(n_2962),
.Y(n_4496)
);

A2O1A1Ixp33_ASAP7_75t_L g4497 ( 
.A1(n_4103),
.A2(n_1149),
.B(n_1153),
.C(n_1136),
.Y(n_4497)
);

CKINVDCx8_ASAP7_75t_R g4498 ( 
.A(n_3972),
.Y(n_4498)
);

AOI21xp5_ASAP7_75t_L g4499 ( 
.A1(n_4093),
.A2(n_3007),
.B(n_2981),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_3914),
.B(n_3206),
.Y(n_4500)
);

AOI22xp5_ASAP7_75t_L g4501 ( 
.A1(n_4017),
.A2(n_1244),
.B1(n_1245),
.B2(n_1243),
.Y(n_4501)
);

INVx3_ASAP7_75t_L g4502 ( 
.A(n_4113),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_SL g4503 ( 
.A(n_4001),
.B(n_2976),
.Y(n_4503)
);

AOI22xp5_ASAP7_75t_L g4504 ( 
.A1(n_4017),
.A2(n_1248),
.B1(n_1245),
.B2(n_761),
.Y(n_4504)
);

INVx4_ASAP7_75t_L g4505 ( 
.A(n_4113),
.Y(n_4505)
);

AOI21xp5_ASAP7_75t_L g4506 ( 
.A1(n_4093),
.A2(n_3007),
.B(n_2981),
.Y(n_4506)
);

BUFx2_ASAP7_75t_L g4507 ( 
.A(n_4010),
.Y(n_4507)
);

NOR2xp33_ASAP7_75t_L g4508 ( 
.A(n_4140),
.B(n_1248),
.Y(n_4508)
);

A2O1A1Ixp33_ASAP7_75t_L g4509 ( 
.A1(n_4162),
.A2(n_1153),
.B(n_1156),
.C(n_1149),
.Y(n_4509)
);

NAND2xp5_ASAP7_75t_SL g4510 ( 
.A(n_4001),
.B(n_2976),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_3905),
.B(n_1156),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_4004),
.Y(n_4512)
);

INVx2_ASAP7_75t_L g4513 ( 
.A(n_4029),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4083),
.B(n_3206),
.Y(n_4514)
);

BUFx2_ASAP7_75t_L g4515 ( 
.A(n_4010),
.Y(n_4515)
);

CKINVDCx8_ASAP7_75t_R g4516 ( 
.A(n_3993),
.Y(n_4516)
);

AOI21xp5_ASAP7_75t_L g4517 ( 
.A1(n_3859),
.A2(n_3007),
.B(n_2981),
.Y(n_4517)
);

INVx2_ASAP7_75t_L g4518 ( 
.A(n_4034),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_3897),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4083),
.B(n_3217),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4085),
.B(n_3217),
.Y(n_4521)
);

HB1xp67_ASAP7_75t_L g4522 ( 
.A(n_4085),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_3898),
.Y(n_4523)
);

BUFx3_ASAP7_75t_L g4524 ( 
.A(n_3995),
.Y(n_4524)
);

A2O1A1Ixp33_ASAP7_75t_L g4525 ( 
.A1(n_4163),
.A2(n_1163),
.B(n_1165),
.C(n_1157),
.Y(n_4525)
);

AOI21xp5_ASAP7_75t_L g4526 ( 
.A1(n_3859),
.A2(n_3057),
.B(n_3036),
.Y(n_4526)
);

HB1xp67_ASAP7_75t_L g4527 ( 
.A(n_3899),
.Y(n_4527)
);

NAND3xp33_ASAP7_75t_SL g4528 ( 
.A(n_3920),
.B(n_759),
.C(n_753),
.Y(n_4528)
);

HB1xp67_ASAP7_75t_L g4529 ( 
.A(n_3926),
.Y(n_4529)
);

NOR2xp33_ASAP7_75t_L g4530 ( 
.A(n_4140),
.B(n_4145),
.Y(n_4530)
);

O2A1O1Ixp33_ASAP7_75t_L g4531 ( 
.A1(n_3908),
.A2(n_1157),
.B(n_1165),
.C(n_1163),
.Y(n_4531)
);

OAI22xp5_ASAP7_75t_L g4532 ( 
.A1(n_4164),
.A2(n_1180),
.B1(n_1192),
.B2(n_1174),
.Y(n_4532)
);

OAI21xp5_ASAP7_75t_L g4533 ( 
.A1(n_4164),
.A2(n_3225),
.B(n_3190),
.Y(n_4533)
);

AOI21xp5_ASAP7_75t_L g4534 ( 
.A1(n_3859),
.A2(n_3057),
.B(n_3036),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_3933),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_3935),
.Y(n_4536)
);

O2A1O1Ixp5_ASAP7_75t_L g4537 ( 
.A1(n_4015),
.A2(n_3680),
.B(n_3608),
.C(n_3293),
.Y(n_4537)
);

BUFx2_ASAP7_75t_L g4538 ( 
.A(n_3948),
.Y(n_4538)
);

OAI22x1_ASAP7_75t_L g4539 ( 
.A1(n_4047),
.A2(n_1180),
.B1(n_1192),
.B2(n_1174),
.Y(n_4539)
);

A2O1A1Ixp33_ASAP7_75t_L g4540 ( 
.A1(n_3962),
.A2(n_1198),
.B(n_1199),
.C(n_1193),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_SL g4541 ( 
.A(n_4145),
.B(n_2988),
.Y(n_4541)
);

NOR2xp33_ASAP7_75t_L g4542 ( 
.A(n_4016),
.B(n_765),
.Y(n_4542)
);

O2A1O1Ixp33_ASAP7_75t_L g4543 ( 
.A1(n_3943),
.A2(n_1193),
.B(n_1199),
.C(n_1198),
.Y(n_4543)
);

OAI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_4165),
.A2(n_1206),
.B1(n_1209),
.B2(n_1202),
.Y(n_4544)
);

AOI21xp33_ASAP7_75t_L g4545 ( 
.A1(n_4165),
.A2(n_2493),
.B(n_2995),
.Y(n_4545)
);

NAND2x1p5_ASAP7_75t_L g4546 ( 
.A(n_4113),
.B(n_3248),
.Y(n_4546)
);

NOR2xp33_ASAP7_75t_L g4547 ( 
.A(n_4016),
.B(n_766),
.Y(n_4547)
);

INVxp67_ASAP7_75t_L g4548 ( 
.A(n_4073),
.Y(n_4548)
);

CKINVDCx20_ASAP7_75t_R g4549 ( 
.A(n_3927),
.Y(n_4549)
);

OAI22xp5_ASAP7_75t_L g4550 ( 
.A1(n_3944),
.A2(n_1206),
.B1(n_1209),
.B2(n_1202),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_4056),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_SL g4552 ( 
.A(n_4007),
.B(n_2988),
.Y(n_4552)
);

AOI21xp5_ASAP7_75t_L g4553 ( 
.A1(n_4026),
.A2(n_3057),
.B(n_3036),
.Y(n_4553)
);

BUFx2_ASAP7_75t_L g4554 ( 
.A(n_3948),
.Y(n_4554)
);

AOI21xp5_ASAP7_75t_L g4555 ( 
.A1(n_3826),
.A2(n_3079),
.B(n_3059),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_3955),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_3979),
.Y(n_4557)
);

AOI21xp5_ASAP7_75t_L g4558 ( 
.A1(n_3826),
.A2(n_3079),
.B(n_3059),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_3980),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4066),
.Y(n_4560)
);

AOI21xp5_ASAP7_75t_L g4561 ( 
.A1(n_3826),
.A2(n_3079),
.B(n_3059),
.Y(n_4561)
);

AOI21xp5_ASAP7_75t_L g4562 ( 
.A1(n_4068),
.A2(n_3097),
.B(n_3094),
.Y(n_4562)
);

AOI22xp5_ASAP7_75t_L g4563 ( 
.A1(n_3877),
.A2(n_774),
.B1(n_778),
.B2(n_767),
.Y(n_4563)
);

NOR2xp33_ASAP7_75t_L g4564 ( 
.A(n_4073),
.B(n_769),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4068),
.A2(n_3097),
.B(n_3094),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4072),
.Y(n_4566)
);

NAND3xp33_ASAP7_75t_SL g4567 ( 
.A(n_3982),
.B(n_784),
.C(n_780),
.Y(n_4567)
);

OAI21x1_ASAP7_75t_L g4568 ( 
.A1(n_4090),
.A2(n_3067),
.B(n_3680),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4099),
.B(n_1210),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_3962),
.B(n_2957),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4527),
.Y(n_4571)
);

AOI22xp33_ASAP7_75t_SL g4572 ( 
.A1(n_4184),
.A2(n_4097),
.B1(n_4011),
.B2(n_4018),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4219),
.B(n_4005),
.Y(n_4573)
);

INVx3_ASAP7_75t_L g4574 ( 
.A(n_4437),
.Y(n_4574)
);

OR2x6_ASAP7_75t_L g4575 ( 
.A(n_4440),
.B(n_3878),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_SL g4576 ( 
.A(n_4219),
.B(n_4212),
.Y(n_4576)
);

AND2x2_ASAP7_75t_L g4577 ( 
.A(n_4183),
.B(n_4021),
.Y(n_4577)
);

CKINVDCx5p33_ASAP7_75t_R g4578 ( 
.A(n_4278),
.Y(n_4578)
);

INVx2_ASAP7_75t_L g4579 ( 
.A(n_4189),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4529),
.Y(n_4580)
);

O2A1O1Ixp33_ASAP7_75t_SL g4581 ( 
.A1(n_4549),
.A2(n_1216),
.B(n_1218),
.C(n_1210),
.Y(n_4581)
);

O2A1O1Ixp33_ASAP7_75t_L g4582 ( 
.A1(n_4234),
.A2(n_1216),
.B(n_1220),
.C(n_1218),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4416),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4522),
.Y(n_4584)
);

BUFx12f_ASAP7_75t_L g4585 ( 
.A(n_4348),
.Y(n_4585)
);

INVx4_ASAP7_75t_L g4586 ( 
.A(n_4408),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4242),
.B(n_4022),
.Y(n_4587)
);

INVxp67_ASAP7_75t_SL g4588 ( 
.A(n_4455),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4174),
.Y(n_4589)
);

INVx2_ASAP7_75t_SL g4590 ( 
.A(n_4383),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4186),
.Y(n_4591)
);

INVx3_ASAP7_75t_L g4592 ( 
.A(n_4437),
.Y(n_4592)
);

BUFx8_ASAP7_75t_L g4593 ( 
.A(n_4233),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4192),
.Y(n_4594)
);

INVx4_ASAP7_75t_L g4595 ( 
.A(n_4408),
.Y(n_4595)
);

INVx3_ASAP7_75t_L g4596 ( 
.A(n_4502),
.Y(n_4596)
);

NOR2xp33_ASAP7_75t_L g4597 ( 
.A(n_4203),
.B(n_3868),
.Y(n_4597)
);

BUFx6f_ASAP7_75t_L g4598 ( 
.A(n_4453),
.Y(n_4598)
);

INVx3_ASAP7_75t_L g4599 ( 
.A(n_4502),
.Y(n_4599)
);

BUFx2_ASAP7_75t_L g4600 ( 
.A(n_4214),
.Y(n_4600)
);

AOI21xp5_ASAP7_75t_L g4601 ( 
.A1(n_4176),
.A2(n_3097),
.B(n_3094),
.Y(n_4601)
);

INVx3_ASAP7_75t_L g4602 ( 
.A(n_4447),
.Y(n_4602)
);

AOI22xp33_ASAP7_75t_L g4603 ( 
.A1(n_4228),
.A2(n_4097),
.B1(n_4076),
.B2(n_4091),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4230),
.Y(n_4604)
);

BUFx12f_ASAP7_75t_L g4605 ( 
.A(n_4368),
.Y(n_4605)
);

OAI22xp5_ASAP7_75t_L g4606 ( 
.A1(n_4237),
.A2(n_4030),
.B1(n_4039),
.B2(n_4031),
.Y(n_4606)
);

AND2x4_ASAP7_75t_L g4607 ( 
.A(n_4198),
.B(n_3925),
.Y(n_4607)
);

A2O1A1Ixp33_ASAP7_75t_L g4608 ( 
.A1(n_4178),
.A2(n_4053),
.B(n_4040),
.C(n_4051),
.Y(n_4608)
);

BUFx2_ASAP7_75t_L g4609 ( 
.A(n_4220),
.Y(n_4609)
);

OAI22xp5_ASAP7_75t_L g4610 ( 
.A1(n_4302),
.A2(n_4050),
.B1(n_4062),
.B2(n_4054),
.Y(n_4610)
);

HB1xp67_ASAP7_75t_L g4611 ( 
.A(n_4171),
.Y(n_4611)
);

OAI221xp5_ASAP7_75t_L g4612 ( 
.A1(n_4249),
.A2(n_1224),
.B1(n_1233),
.B2(n_1222),
.C(n_1220),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4238),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4224),
.Y(n_4614)
);

O2A1O1Ixp33_ASAP7_75t_L g4615 ( 
.A1(n_4195),
.A2(n_1222),
.B(n_1233),
.C(n_1224),
.Y(n_4615)
);

BUFx2_ASAP7_75t_L g4616 ( 
.A(n_4258),
.Y(n_4616)
);

BUFx12f_ASAP7_75t_L g4617 ( 
.A(n_4454),
.Y(n_4617)
);

CKINVDCx6p67_ASAP7_75t_R g4618 ( 
.A(n_4427),
.Y(n_4618)
);

INVx3_ASAP7_75t_L g4619 ( 
.A(n_4447),
.Y(n_4619)
);

AOI22xp33_ASAP7_75t_L g4620 ( 
.A1(n_4172),
.A2(n_4078),
.B1(n_4107),
.B2(n_4102),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_4273),
.B(n_4064),
.Y(n_4621)
);

A2O1A1Ixp33_ASAP7_75t_L g4622 ( 
.A1(n_4494),
.A2(n_4086),
.B(n_3991),
.C(n_4081),
.Y(n_4622)
);

BUFx6f_ASAP7_75t_L g4623 ( 
.A(n_4453),
.Y(n_4623)
);

HB1xp67_ASAP7_75t_L g4624 ( 
.A(n_4229),
.Y(n_4624)
);

BUFx6f_ASAP7_75t_L g4625 ( 
.A(n_4453),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4225),
.Y(n_4626)
);

NOR2xp33_ASAP7_75t_L g4627 ( 
.A(n_4216),
.B(n_3868),
.Y(n_4627)
);

INVx2_ASAP7_75t_L g4628 ( 
.A(n_4265),
.Y(n_4628)
);

BUFx6f_ASAP7_75t_L g4629 ( 
.A(n_4516),
.Y(n_4629)
);

AO22x1_ASAP7_75t_L g4630 ( 
.A1(n_4430),
.A2(n_4217),
.B1(n_4269),
.B2(n_4194),
.Y(n_4630)
);

AOI22xp33_ASAP7_75t_L g4631 ( 
.A1(n_4480),
.A2(n_4119),
.B1(n_4122),
.B2(n_4115),
.Y(n_4631)
);

NAND2x1p5_ASAP7_75t_L g4632 ( 
.A(n_4200),
.B(n_4442),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_4294),
.B(n_4149),
.Y(n_4633)
);

AND2x4_ASAP7_75t_L g4634 ( 
.A(n_4200),
.B(n_4015),
.Y(n_4634)
);

INVxp67_ASAP7_75t_L g4635 ( 
.A(n_4273),
.Y(n_4635)
);

AOI22xp5_ASAP7_75t_L g4636 ( 
.A1(n_4412),
.A2(n_3877),
.B1(n_4161),
.B2(n_4081),
.Y(n_4636)
);

OAI22xp33_ASAP7_75t_L g4637 ( 
.A1(n_4226),
.A2(n_1240),
.B1(n_1238),
.B2(n_2995),
.Y(n_4637)
);

CKINVDCx20_ASAP7_75t_R g4638 ( 
.A(n_4268),
.Y(n_4638)
);

INVx1_ASAP7_75t_SL g4639 ( 
.A(n_4289),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4260),
.Y(n_4640)
);

AOI22xp33_ASAP7_75t_L g4641 ( 
.A1(n_4226),
.A2(n_4121),
.B1(n_4124),
.B2(n_4110),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_4289),
.B(n_4111),
.Y(n_4642)
);

NAND2x1p5_ASAP7_75t_L g4643 ( 
.A(n_4200),
.B(n_3984),
.Y(n_4643)
);

BUFx6f_ASAP7_75t_L g4644 ( 
.A(n_4284),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4274),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4276),
.Y(n_4646)
);

BUFx12f_ASAP7_75t_L g4647 ( 
.A(n_4476),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4282),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4293),
.Y(n_4649)
);

INVx2_ASAP7_75t_L g4650 ( 
.A(n_4285),
.Y(n_4650)
);

AOI22xp33_ASAP7_75t_L g4651 ( 
.A1(n_4182),
.A2(n_4136),
.B1(n_4129),
.B2(n_4141),
.Y(n_4651)
);

INVxp67_ASAP7_75t_SL g4652 ( 
.A(n_4253),
.Y(n_4652)
);

OR2x6_ASAP7_75t_L g4653 ( 
.A(n_4449),
.B(n_4235),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4316),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4323),
.Y(n_4655)
);

BUFx2_ASAP7_75t_L g4656 ( 
.A(n_4291),
.Y(n_4656)
);

BUFx6f_ASAP7_75t_L g4657 ( 
.A(n_4284),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4344),
.Y(n_4658)
);

INVx4_ASAP7_75t_L g4659 ( 
.A(n_4193),
.Y(n_4659)
);

INVx2_ASAP7_75t_SL g4660 ( 
.A(n_4524),
.Y(n_4660)
);

NOR2xp33_ASAP7_75t_L g4661 ( 
.A(n_4340),
.B(n_3941),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4369),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_4295),
.Y(n_4663)
);

OAI22x1_ASAP7_75t_L g4664 ( 
.A1(n_4315),
.A2(n_1240),
.B1(n_1238),
.B2(n_4161),
.Y(n_4664)
);

BUFx6f_ASAP7_75t_L g4665 ( 
.A(n_4386),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4170),
.B(n_4111),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4301),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4170),
.B(n_4112),
.Y(n_4668)
);

BUFx2_ASAP7_75t_SL g4669 ( 
.A(n_4467),
.Y(n_4669)
);

CKINVDCx5p33_ASAP7_75t_R g4670 ( 
.A(n_4250),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_4318),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4331),
.Y(n_4672)
);

INVx2_ASAP7_75t_L g4673 ( 
.A(n_4335),
.Y(n_4673)
);

OAI22xp5_ASAP7_75t_SL g4674 ( 
.A1(n_4489),
.A2(n_3958),
.B1(n_3961),
.B2(n_3941),
.Y(n_4674)
);

OAI22xp33_ASAP7_75t_L g4675 ( 
.A1(n_4240),
.A2(n_2995),
.B1(n_3961),
.B2(n_3958),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4204),
.B(n_4112),
.Y(n_4676)
);

AO21x1_ASAP7_75t_L g4677 ( 
.A1(n_4325),
.A2(n_1361),
.B(n_1359),
.Y(n_4677)
);

AOI22xp5_ASAP7_75t_L g4678 ( 
.A1(n_4297),
.A2(n_3877),
.B1(n_4002),
.B2(n_3993),
.Y(n_4678)
);

NAND3xp33_ASAP7_75t_L g4679 ( 
.A(n_4325),
.B(n_1529),
.C(n_1528),
.Y(n_4679)
);

BUFx12f_ASAP7_75t_L g4680 ( 
.A(n_4207),
.Y(n_4680)
);

INVx1_ASAP7_75t_SL g4681 ( 
.A(n_4308),
.Y(n_4681)
);

BUFx6f_ASAP7_75t_L g4682 ( 
.A(n_4193),
.Y(n_4682)
);

OAI22xp33_ASAP7_75t_L g4683 ( 
.A1(n_4470),
.A2(n_4181),
.B1(n_4191),
.B2(n_4501),
.Y(n_4683)
);

OAI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_4270),
.A2(n_3893),
.B1(n_3830),
.B2(n_3990),
.Y(n_4684)
);

INVx1_ASAP7_75t_SL g4685 ( 
.A(n_4326),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4204),
.B(n_4135),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_SL g4687 ( 
.A(n_4218),
.B(n_3948),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4213),
.B(n_4135),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_4218),
.B(n_4148),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4373),
.Y(n_4690)
);

AND2x6_ASAP7_75t_L g4691 ( 
.A(n_4361),
.B(n_3984),
.Y(n_4691)
);

BUFx2_ASAP7_75t_L g4692 ( 
.A(n_4351),
.Y(n_4692)
);

INVx4_ASAP7_75t_L g4693 ( 
.A(n_4193),
.Y(n_4693)
);

BUFx2_ASAP7_75t_L g4694 ( 
.A(n_4370),
.Y(n_4694)
);

INVx2_ASAP7_75t_SL g4695 ( 
.A(n_4394),
.Y(n_4695)
);

CKINVDCx5p33_ASAP7_75t_R g4696 ( 
.A(n_4337),
.Y(n_4696)
);

HB1xp67_ASAP7_75t_L g4697 ( 
.A(n_4329),
.Y(n_4697)
);

AOI21xp5_ASAP7_75t_L g4698 ( 
.A1(n_4177),
.A2(n_3165),
.B(n_3147),
.Y(n_4698)
);

AOI21xp5_ASAP7_75t_L g4699 ( 
.A1(n_4179),
.A2(n_3165),
.B(n_3147),
.Y(n_4699)
);

AND2x4_ASAP7_75t_L g4700 ( 
.A(n_4200),
.B(n_4074),
.Y(n_4700)
);

AOI21xp33_ASAP7_75t_L g4701 ( 
.A1(n_4180),
.A2(n_2493),
.B(n_4154),
.Y(n_4701)
);

NOR2xp33_ASAP7_75t_L g4702 ( 
.A(n_4311),
.B(n_3990),
.Y(n_4702)
);

INVx4_ASAP7_75t_L g4703 ( 
.A(n_4196),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4294),
.B(n_3977),
.Y(n_4704)
);

NAND2x2_ASAP7_75t_L g4705 ( 
.A(n_4495),
.B(n_4),
.Y(n_4705)
);

INVx2_ASAP7_75t_L g4706 ( 
.A(n_4374),
.Y(n_4706)
);

NOR2xp33_ASAP7_75t_L g4707 ( 
.A(n_4173),
.B(n_785),
.Y(n_4707)
);

CKINVDCx8_ASAP7_75t_R g4708 ( 
.A(n_4245),
.Y(n_4708)
);

NOR2xp33_ASAP7_75t_SL g4709 ( 
.A(n_4498),
.B(n_3877),
.Y(n_4709)
);

BUFx4f_ASAP7_75t_L g4710 ( 
.A(n_4175),
.Y(n_4710)
);

HB1xp67_ASAP7_75t_L g4711 ( 
.A(n_4329),
.Y(n_4711)
);

OAI21x1_ASAP7_75t_L g4712 ( 
.A1(n_4197),
.A2(n_3893),
.B(n_4156),
.Y(n_4712)
);

AND2x4_ASAP7_75t_L g4713 ( 
.A(n_4449),
.B(n_4235),
.Y(n_4713)
);

INVx8_ASAP7_75t_L g4714 ( 
.A(n_4459),
.Y(n_4714)
);

BUFx4f_ASAP7_75t_L g4715 ( 
.A(n_4175),
.Y(n_4715)
);

AOI22xp5_ASAP7_75t_L g4716 ( 
.A1(n_4248),
.A2(n_4002),
.B1(n_789),
.B2(n_790),
.Y(n_4716)
);

INVx5_ASAP7_75t_L g4717 ( 
.A(n_4235),
.Y(n_4717)
);

INVx3_ASAP7_75t_L g4718 ( 
.A(n_4505),
.Y(n_4718)
);

INVx1_ASAP7_75t_SL g4719 ( 
.A(n_4391),
.Y(n_4719)
);

INVx3_ASAP7_75t_L g4720 ( 
.A(n_4505),
.Y(n_4720)
);

NOR3xp33_ASAP7_75t_L g4721 ( 
.A(n_4263),
.B(n_1612),
.C(n_1611),
.Y(n_4721)
);

AND2x2_ASAP7_75t_L g4722 ( 
.A(n_4391),
.B(n_3977),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4382),
.Y(n_4723)
);

AOI22xp33_ASAP7_75t_L g4724 ( 
.A1(n_4221),
.A2(n_3235),
.B1(n_3247),
.B2(n_3232),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4379),
.Y(n_4725)
);

AOI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_4190),
.A2(n_3165),
.B(n_3147),
.Y(n_4726)
);

BUFx3_ASAP7_75t_L g4727 ( 
.A(n_4376),
.Y(n_4727)
);

BUFx3_ASAP7_75t_L g4728 ( 
.A(n_4409),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4396),
.Y(n_4729)
);

INVx2_ASAP7_75t_L g4730 ( 
.A(n_4405),
.Y(n_4730)
);

INVx2_ASAP7_75t_L g4731 ( 
.A(n_4411),
.Y(n_4731)
);

AOI22xp33_ASAP7_75t_SL g4732 ( 
.A1(n_4181),
.A2(n_794),
.B1(n_795),
.B2(n_788),
.Y(n_4732)
);

INVx5_ASAP7_75t_L g4733 ( 
.A(n_4449),
.Y(n_4733)
);

BUFx6f_ASAP7_75t_L g4734 ( 
.A(n_4196),
.Y(n_4734)
);

OR2x2_ASAP7_75t_L g4735 ( 
.A(n_4328),
.B(n_3977),
.Y(n_4735)
);

NOR2xp67_ASAP7_75t_SL g4736 ( 
.A(n_4387),
.B(n_4020),
.Y(n_4736)
);

CKINVDCx8_ASAP7_75t_R g4737 ( 
.A(n_4384),
.Y(n_4737)
);

BUFx2_ASAP7_75t_L g4738 ( 
.A(n_4305),
.Y(n_4738)
);

BUFx3_ASAP7_75t_L g4739 ( 
.A(n_4430),
.Y(n_4739)
);

NOR2xp33_ASAP7_75t_L g4740 ( 
.A(n_4215),
.B(n_793),
.Y(n_4740)
);

INVx5_ASAP7_75t_L g4741 ( 
.A(n_4387),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4402),
.Y(n_4742)
);

HB1xp67_ASAP7_75t_L g4743 ( 
.A(n_4342),
.Y(n_4743)
);

HB1xp67_ASAP7_75t_L g4744 ( 
.A(n_4342),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4419),
.Y(n_4745)
);

CKINVDCx5p33_ASAP7_75t_R g4746 ( 
.A(n_4185),
.Y(n_4746)
);

BUFx5_ASAP7_75t_L g4747 ( 
.A(n_4169),
.Y(n_4747)
);

AND2x2_ASAP7_75t_SL g4748 ( 
.A(n_4475),
.B(n_4074),
.Y(n_4748)
);

NOR2xp33_ASAP7_75t_SL g4749 ( 
.A(n_4477),
.B(n_4116),
.Y(n_4749)
);

INVx2_ASAP7_75t_SL g4750 ( 
.A(n_4247),
.Y(n_4750)
);

AO31x2_ASAP7_75t_L g4751 ( 
.A1(n_4241),
.A2(n_3235),
.A3(n_3247),
.B(n_3232),
.Y(n_4751)
);

CKINVDCx8_ASAP7_75t_R g4752 ( 
.A(n_4384),
.Y(n_4752)
);

BUFx3_ASAP7_75t_L g4753 ( 
.A(n_4196),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4328),
.B(n_4020),
.Y(n_4754)
);

AO22x1_ASAP7_75t_L g4755 ( 
.A1(n_4459),
.A2(n_4002),
.B1(n_4139),
.B2(n_4116),
.Y(n_4755)
);

INVx5_ASAP7_75t_L g4756 ( 
.A(n_4387),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4403),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4423),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4239),
.B(n_4020),
.Y(n_4759)
);

INVx6_ASAP7_75t_L g4760 ( 
.A(n_4254),
.Y(n_4760)
);

BUFx3_ASAP7_75t_L g4761 ( 
.A(n_4201),
.Y(n_4761)
);

BUFx12f_ASAP7_75t_L g4762 ( 
.A(n_4201),
.Y(n_4762)
);

AND2x2_ASAP7_75t_SL g4763 ( 
.A(n_4246),
.B(n_4139),
.Y(n_4763)
);

OAI22xp5_ASAP7_75t_L g4764 ( 
.A1(n_4270),
.A2(n_798),
.B1(n_799),
.B2(n_796),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4243),
.B(n_4390),
.Y(n_4765)
);

OAI22xp33_ASAP7_75t_L g4766 ( 
.A1(n_4191),
.A2(n_801),
.B1(n_807),
.B2(n_797),
.Y(n_4766)
);

CKINVDCx8_ASAP7_75t_R g4767 ( 
.A(n_4201),
.Y(n_4767)
);

OR2x6_ASAP7_75t_L g4768 ( 
.A(n_4395),
.B(n_4027),
.Y(n_4768)
);

INVx3_ASAP7_75t_L g4769 ( 
.A(n_4389),
.Y(n_4769)
);

AOI22xp33_ASAP7_75t_L g4770 ( 
.A1(n_4236),
.A2(n_3263),
.B1(n_3281),
.B2(n_3259),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_L g4771 ( 
.A(n_4309),
.B(n_4027),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4438),
.Y(n_4772)
);

BUFx3_ASAP7_75t_L g4773 ( 
.A(n_4211),
.Y(n_4773)
);

INVx2_ASAP7_75t_L g4774 ( 
.A(n_4421),
.Y(n_4774)
);

BUFx12f_ASAP7_75t_L g4775 ( 
.A(n_4211),
.Y(n_4775)
);

AOI21xp5_ASAP7_75t_L g4776 ( 
.A1(n_4187),
.A2(n_3207),
.B(n_3201),
.Y(n_4776)
);

INVx2_ASAP7_75t_SL g4777 ( 
.A(n_4211),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4439),
.Y(n_4778)
);

INVx3_ASAP7_75t_L g4779 ( 
.A(n_4389),
.Y(n_4779)
);

OR2x6_ASAP7_75t_SL g4780 ( 
.A(n_4550),
.B(n_836),
.Y(n_4780)
);

INVx1_ASAP7_75t_SL g4781 ( 
.A(n_4538),
.Y(n_4781)
);

AND2x2_ASAP7_75t_L g4782 ( 
.A(n_4530),
.B(n_4027),
.Y(n_4782)
);

INVx8_ASAP7_75t_L g4783 ( 
.A(n_4418),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4444),
.Y(n_4784)
);

O2A1O1Ixp5_ASAP7_75t_L g4785 ( 
.A1(n_4251),
.A2(n_4252),
.B(n_4334),
.C(n_4256),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4451),
.Y(n_4786)
);

AOI21xp5_ASAP7_75t_L g4787 ( 
.A1(n_4251),
.A2(n_3207),
.B(n_3201),
.Y(n_4787)
);

INVx2_ASAP7_75t_L g4788 ( 
.A(n_4450),
.Y(n_4788)
);

HB1xp67_ASAP7_75t_L g4789 ( 
.A(n_4355),
.Y(n_4789)
);

AND2x4_ASAP7_75t_L g4790 ( 
.A(n_4298),
.B(n_4033),
.Y(n_4790)
);

BUFx8_ASAP7_75t_L g4791 ( 
.A(n_4511),
.Y(n_4791)
);

INVx1_ASAP7_75t_SL g4792 ( 
.A(n_4554),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4460),
.Y(n_4793)
);

BUFx2_ASAP7_75t_L g4794 ( 
.A(n_4507),
.Y(n_4794)
);

BUFx3_ASAP7_75t_L g4795 ( 
.A(n_4257),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_4491),
.Y(n_4796)
);

INVx2_ASAP7_75t_L g4797 ( 
.A(n_4512),
.Y(n_4797)
);

HB1xp67_ASAP7_75t_L g4798 ( 
.A(n_4355),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4462),
.Y(n_4799)
);

NAND2xp5_ASAP7_75t_L g4800 ( 
.A(n_4377),
.B(n_4033),
.Y(n_4800)
);

INVx2_ASAP7_75t_L g4801 ( 
.A(n_4513),
.Y(n_4801)
);

BUFx6f_ASAP7_75t_L g4802 ( 
.A(n_4257),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4465),
.Y(n_4803)
);

INVx3_ASAP7_75t_L g4804 ( 
.A(n_4389),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4466),
.Y(n_4805)
);

BUFx6f_ASAP7_75t_L g4806 ( 
.A(n_4257),
.Y(n_4806)
);

O2A1O1Ixp33_ASAP7_75t_L g4807 ( 
.A1(n_4231),
.A2(n_4202),
.B(n_4332),
.C(n_4327),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4519),
.Y(n_4808)
);

OAI22xp5_ASAP7_75t_L g4809 ( 
.A1(n_4474),
.A2(n_840),
.B1(n_842),
.B2(n_837),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_L g4810 ( 
.A(n_4271),
.B(n_4227),
.Y(n_4810)
);

BUFx2_ASAP7_75t_L g4811 ( 
.A(n_4515),
.Y(n_4811)
);

HB1xp67_ASAP7_75t_L g4812 ( 
.A(n_4367),
.Y(n_4812)
);

BUFx6f_ASAP7_75t_L g4813 ( 
.A(n_4259),
.Y(n_4813)
);

BUFx8_ASAP7_75t_SL g4814 ( 
.A(n_4259),
.Y(n_4814)
);

AND2x4_ASAP7_75t_L g4815 ( 
.A(n_4298),
.B(n_4033),
.Y(n_4815)
);

INVx2_ASAP7_75t_L g4816 ( 
.A(n_4518),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4523),
.Y(n_4817)
);

OR2x6_ASAP7_75t_L g4818 ( 
.A(n_4367),
.B(n_4036),
.Y(n_4818)
);

INVx5_ASAP7_75t_L g4819 ( 
.A(n_4169),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4551),
.Y(n_4820)
);

A2O1A1Ixp33_ASAP7_75t_L g4821 ( 
.A1(n_4364),
.A2(n_1614),
.B(n_1617),
.C(n_1613),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4535),
.Y(n_4822)
);

AOI21xp5_ASAP7_75t_L g4823 ( 
.A1(n_4426),
.A2(n_3207),
.B(n_3201),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_L g4824 ( 
.A(n_4222),
.B(n_4036),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4536),
.Y(n_4825)
);

CKINVDCx8_ASAP7_75t_R g4826 ( 
.A(n_4259),
.Y(n_4826)
);

AND2x2_ASAP7_75t_L g4827 ( 
.A(n_4244),
.B(n_4036),
.Y(n_4827)
);

BUFx6f_ASAP7_75t_L g4828 ( 
.A(n_4303),
.Y(n_4828)
);

CKINVDCx5p33_ASAP7_75t_R g4829 ( 
.A(n_4445),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4548),
.B(n_4067),
.Y(n_4830)
);

AND3x1_ASAP7_75t_SL g4831 ( 
.A(n_4556),
.B(n_1620),
.C(n_1619),
.Y(n_4831)
);

INVx4_ASAP7_75t_L g4832 ( 
.A(n_4303),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4557),
.Y(n_4833)
);

INVx3_ASAP7_75t_L g4834 ( 
.A(n_4365),
.Y(n_4834)
);

OAI221xp5_ASAP7_75t_L g4835 ( 
.A1(n_4504),
.A2(n_892),
.B1(n_911),
.B2(n_855),
.C(n_843),
.Y(n_4835)
);

INVx6_ASAP7_75t_L g4836 ( 
.A(n_4254),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4222),
.B(n_4067),
.Y(n_4837)
);

INVx2_ASAP7_75t_L g4838 ( 
.A(n_4560),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4559),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4275),
.Y(n_4840)
);

AND2x2_ASAP7_75t_SL g4841 ( 
.A(n_4246),
.B(n_4067),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4280),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4210),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4569),
.B(n_4094),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4392),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4415),
.Y(n_4846)
);

AND2x4_ASAP7_75t_L g4847 ( 
.A(n_4169),
.B(n_4094),
.Y(n_4847)
);

HB1xp67_ASAP7_75t_L g4848 ( 
.A(n_4375),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4417),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4366),
.B(n_4188),
.Y(n_4850)
);

INVx1_ASAP7_75t_SL g4851 ( 
.A(n_4349),
.Y(n_4851)
);

NAND2x1p5_ASAP7_75t_L g4852 ( 
.A(n_4372),
.B(n_4094),
.Y(n_4852)
);

AND2x4_ASAP7_75t_L g4853 ( 
.A(n_4169),
.B(n_4126),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4443),
.Y(n_4854)
);

NAND2xp5_ASAP7_75t_L g4855 ( 
.A(n_4366),
.B(n_4126),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4452),
.Y(n_4856)
);

AOI22xp33_ASAP7_75t_SL g4857 ( 
.A1(n_4532),
.A2(n_846),
.B1(n_847),
.B2(n_838),
.Y(n_4857)
);

INVxp67_ASAP7_75t_L g4858 ( 
.A(n_4375),
.Y(n_4858)
);

BUFx3_ASAP7_75t_L g4859 ( 
.A(n_4303),
.Y(n_4859)
);

BUFx2_ASAP7_75t_L g4860 ( 
.A(n_4262),
.Y(n_4860)
);

BUFx3_ASAP7_75t_L g4861 ( 
.A(n_4206),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4306),
.B(n_4126),
.Y(n_4862)
);

INVx2_ASAP7_75t_L g4863 ( 
.A(n_4566),
.Y(n_4863)
);

HB1xp67_ASAP7_75t_L g4864 ( 
.A(n_4330),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4463),
.Y(n_4865)
);

NOR2xp67_ASAP7_75t_SL g4866 ( 
.A(n_4336),
.B(n_2988),
.Y(n_4866)
);

INVxp67_ASAP7_75t_L g4867 ( 
.A(n_4307),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_L g4868 ( 
.A(n_4306),
.B(n_4002),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4479),
.Y(n_4869)
);

BUFx6f_ASAP7_75t_L g4870 ( 
.A(n_4418),
.Y(n_4870)
);

HB1xp67_ASAP7_75t_L g4871 ( 
.A(n_4307),
.Y(n_4871)
);

A2O1A1Ixp33_ASAP7_75t_L g4872 ( 
.A1(n_4407),
.A2(n_1623),
.B(n_1626),
.C(n_1621),
.Y(n_4872)
);

A2O1A1Ixp33_ASAP7_75t_L g4873 ( 
.A1(n_4413),
.A2(n_1629),
.B(n_1631),
.C(n_1628),
.Y(n_4873)
);

NOR2xp33_ASAP7_75t_L g4874 ( 
.A(n_4468),
.B(n_844),
.Y(n_4874)
);

INVx4_ASAP7_75t_L g4875 ( 
.A(n_4336),
.Y(n_4875)
);

BUFx6f_ASAP7_75t_L g4876 ( 
.A(n_4206),
.Y(n_4876)
);

OAI22xp5_ASAP7_75t_L g4877 ( 
.A1(n_4327),
.A2(n_852),
.B1(n_853),
.B2(n_849),
.Y(n_4877)
);

INVxp67_ASAP7_75t_SL g4878 ( 
.A(n_4321),
.Y(n_4878)
);

BUFx3_ASAP7_75t_L g4879 ( 
.A(n_4277),
.Y(n_4879)
);

AND2x2_ASAP7_75t_L g4880 ( 
.A(n_4358),
.B(n_1359),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4292),
.B(n_1361),
.Y(n_4881)
);

OR2x2_ASAP7_75t_L g4882 ( 
.A(n_4357),
.B(n_4321),
.Y(n_4882)
);

AND2x2_ASAP7_75t_L g4883 ( 
.A(n_4485),
.B(n_1362),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4484),
.Y(n_4884)
);

AND2x2_ASAP7_75t_L g4885 ( 
.A(n_4508),
.B(n_1362),
.Y(n_4885)
);

BUFx3_ASAP7_75t_L g4886 ( 
.A(n_4277),
.Y(n_4886)
);

INVx2_ASAP7_75t_L g4887 ( 
.A(n_4487),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4500),
.Y(n_4888)
);

A2O1A1Ixp33_ASAP7_75t_L g4889 ( 
.A1(n_4255),
.A2(n_1635),
.B(n_1637),
.C(n_1632),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4514),
.Y(n_4890)
);

BUFx6f_ASAP7_75t_L g4891 ( 
.A(n_4353),
.Y(n_4891)
);

INVx4_ASAP7_75t_L g4892 ( 
.A(n_4353),
.Y(n_4892)
);

CKINVDCx11_ASAP7_75t_R g4893 ( 
.A(n_4361),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4520),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4431),
.B(n_2951),
.Y(n_4895)
);

AND2x4_ASAP7_75t_L g4896 ( 
.A(n_4503),
.B(n_3293),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_SL g4897 ( 
.A(n_4209),
.B(n_3353),
.Y(n_4897)
);

AOI22xp5_ASAP7_75t_L g4898 ( 
.A1(n_4532),
.A2(n_864),
.B1(n_865),
.B2(n_850),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4521),
.Y(n_4899)
);

INVx5_ASAP7_75t_L g4900 ( 
.A(n_4354),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4300),
.Y(n_4901)
);

NAND2xp5_ASAP7_75t_L g4902 ( 
.A(n_4287),
.B(n_2951),
.Y(n_4902)
);

INVx3_ASAP7_75t_L g4903 ( 
.A(n_4359),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4304),
.Y(n_4904)
);

AOI22xp33_ASAP7_75t_L g4905 ( 
.A1(n_4371),
.A2(n_3263),
.B1(n_3281),
.B2(n_3259),
.Y(n_4905)
);

BUFx3_ASAP7_75t_L g4906 ( 
.A(n_4354),
.Y(n_4906)
);

BUFx6f_ASAP7_75t_L g4907 ( 
.A(n_4510),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4469),
.Y(n_4908)
);

AND2x2_ASAP7_75t_SL g4909 ( 
.A(n_4283),
.B(n_3025),
.Y(n_4909)
);

AOI21xp5_ASAP7_75t_L g4910 ( 
.A1(n_4448),
.A2(n_3003),
.B(n_2988),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4570),
.Y(n_4911)
);

AOI22xp5_ASAP7_75t_L g4912 ( 
.A1(n_4544),
.A2(n_871),
.B1(n_877),
.B2(n_869),
.Y(n_4912)
);

BUFx2_ASAP7_75t_L g4913 ( 
.A(n_4482),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4570),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4471),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_L g4916 ( 
.A(n_4312),
.B(n_2951),
.Y(n_4916)
);

BUFx6f_ASAP7_75t_L g4917 ( 
.A(n_4546),
.Y(n_4917)
);

NAND2x1_ASAP7_75t_L g4918 ( 
.A(n_4266),
.B(n_3003),
.Y(n_4918)
);

INVx2_ASAP7_75t_L g4919 ( 
.A(n_4472),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_4371),
.B(n_2951),
.Y(n_4920)
);

INVx5_ASAP7_75t_L g4921 ( 
.A(n_4493),
.Y(n_4921)
);

AND2x4_ASAP7_75t_L g4922 ( 
.A(n_4541),
.B(n_3003),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4435),
.Y(n_4923)
);

AND2x4_ASAP7_75t_L g4924 ( 
.A(n_4288),
.B(n_3003),
.Y(n_4924)
);

AND2x2_ASAP7_75t_L g4925 ( 
.A(n_4542),
.B(n_1365),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4338),
.Y(n_4926)
);

HB1xp67_ASAP7_75t_L g4927 ( 
.A(n_4457),
.Y(n_4927)
);

OAI22xp5_ASAP7_75t_L g4928 ( 
.A1(n_4332),
.A2(n_893),
.B1(n_896),
.B2(n_881),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_4490),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4347),
.Y(n_4930)
);

NAND2x1p5_ASAP7_75t_L g4931 ( 
.A(n_4388),
.B(n_3010),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_L g4932 ( 
.A(n_4398),
.B(n_2957),
.Y(n_4932)
);

INVx2_ASAP7_75t_L g4933 ( 
.A(n_4490),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4490),
.Y(n_4934)
);

OAI222xp33_ASAP7_75t_L g4935 ( 
.A1(n_4544),
.A2(n_902),
.B1(n_898),
.B2(n_905),
.C1(n_901),
.C2(n_885),
.Y(n_4935)
);

AND2x2_ASAP7_75t_L g4936 ( 
.A(n_4547),
.B(n_1365),
.Y(n_4936)
);

BUFx6f_ASAP7_75t_L g4937 ( 
.A(n_4546),
.Y(n_4937)
);

HB1xp67_ASAP7_75t_L g4938 ( 
.A(n_4457),
.Y(n_4938)
);

INVx2_ASAP7_75t_SL g4939 ( 
.A(n_4320),
.Y(n_4939)
);

INVx4_ASAP7_75t_L g4940 ( 
.A(n_4359),
.Y(n_4940)
);

AND2x6_ASAP7_75t_SL g4941 ( 
.A(n_4441),
.B(n_1638),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4296),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_SL g4943 ( 
.A(n_4232),
.B(n_3375),
.Y(n_4943)
);

INVx3_ASAP7_75t_L g4944 ( 
.A(n_4352),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4310),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4492),
.Y(n_4946)
);

NAND2xp5_ASAP7_75t_L g4947 ( 
.A(n_4398),
.B(n_2957),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4564),
.B(n_4223),
.Y(n_4948)
);

INVx1_ASAP7_75t_SL g4949 ( 
.A(n_4400),
.Y(n_4949)
);

AOI22xp33_ASAP7_75t_L g4950 ( 
.A1(n_4433),
.A2(n_3297),
.B1(n_3301),
.B2(n_3292),
.Y(n_4950)
);

CKINVDCx11_ASAP7_75t_R g4951 ( 
.A(n_4550),
.Y(n_4951)
);

OAI22xp5_ASAP7_75t_L g4952 ( 
.A1(n_4341),
.A2(n_913),
.B1(n_917),
.B2(n_910),
.Y(n_4952)
);

BUFx3_ASAP7_75t_L g4953 ( 
.A(n_4345),
.Y(n_4953)
);

NAND2x1p5_ASAP7_75t_L g4954 ( 
.A(n_4422),
.B(n_3010),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4356),
.Y(n_4955)
);

INVx4_ASAP7_75t_L g4956 ( 
.A(n_4552),
.Y(n_4956)
);

OR2x6_ASAP7_75t_L g4957 ( 
.A(n_4399),
.B(n_3010),
.Y(n_4957)
);

INVxp67_ASAP7_75t_L g4958 ( 
.A(n_4281),
.Y(n_4958)
);

CKINVDCx5p33_ASAP7_75t_R g4959 ( 
.A(n_4464),
.Y(n_4959)
);

BUFx8_ASAP7_75t_SL g4960 ( 
.A(n_4456),
.Y(n_4960)
);

AND2x2_ASAP7_75t_L g4961 ( 
.A(n_4539),
.B(n_4261),
.Y(n_4961)
);

AOI21x1_ASAP7_75t_L g4962 ( 
.A1(n_4433),
.A2(n_1532),
.B(n_1531),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4492),
.Y(n_4963)
);

A2O1A1Ixp33_ASAP7_75t_L g4964 ( 
.A1(n_4543),
.A2(n_1640),
.B(n_1643),
.C(n_1639),
.Y(n_4964)
);

A2O1A1Ixp33_ASAP7_75t_L g4965 ( 
.A1(n_4264),
.A2(n_1647),
.B(n_1648),
.C(n_1645),
.Y(n_4965)
);

INVx2_ASAP7_75t_SL g4966 ( 
.A(n_4424),
.Y(n_4966)
);

BUFx6f_ASAP7_75t_L g4967 ( 
.A(n_4432),
.Y(n_4967)
);

BUFx6f_ASAP7_75t_L g4968 ( 
.A(n_4434),
.Y(n_4968)
);

BUFx3_ASAP7_75t_L g4969 ( 
.A(n_4486),
.Y(n_4969)
);

BUFx3_ASAP7_75t_L g4970 ( 
.A(n_4568),
.Y(n_4970)
);

OAI22xp5_ASAP7_75t_L g4971 ( 
.A1(n_4341),
.A2(n_925),
.B1(n_926),
.B2(n_912),
.Y(n_4971)
);

AND2x2_ASAP7_75t_L g4972 ( 
.A(n_4279),
.B(n_1366),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4360),
.Y(n_4973)
);

O2A1O1Ixp33_ASAP7_75t_L g4974 ( 
.A1(n_4362),
.A2(n_1650),
.B(n_1652),
.C(n_1649),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4492),
.Y(n_4975)
);

AOI22xp33_ASAP7_75t_L g4976 ( 
.A1(n_4205),
.A2(n_3297),
.B1(n_3301),
.B2(n_3292),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4286),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4299),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4362),
.B(n_2957),
.Y(n_4979)
);

OR2x2_ASAP7_75t_L g4980 ( 
.A(n_4363),
.B(n_1366),
.Y(n_4980)
);

INVxp67_ASAP7_75t_L g4981 ( 
.A(n_4319),
.Y(n_4981)
);

INVx4_ASAP7_75t_L g4982 ( 
.A(n_4537),
.Y(n_4982)
);

AOI22xp33_ASAP7_75t_L g4983 ( 
.A1(n_4393),
.A2(n_4363),
.B1(n_4481),
.B2(n_4478),
.Y(n_4983)
);

AND2x4_ASAP7_75t_L g4984 ( 
.A(n_4446),
.B(n_3010),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4385),
.B(n_1367),
.Y(n_4985)
);

BUFx2_ASAP7_75t_SL g4986 ( 
.A(n_4461),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4333),
.B(n_1367),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4380),
.Y(n_4988)
);

INVx2_ASAP7_75t_L g4989 ( 
.A(n_4317),
.Y(n_4989)
);

AO21x1_ASAP7_75t_L g4990 ( 
.A1(n_4576),
.A2(n_4683),
.B(n_4766),
.Y(n_4990)
);

O2A1O1Ixp33_ASAP7_75t_L g4991 ( 
.A1(n_4809),
.A2(n_4497),
.B(n_4199),
.C(n_4509),
.Y(n_4991)
);

A2O1A1Ixp33_ASAP7_75t_L g4992 ( 
.A1(n_4807),
.A2(n_4563),
.B(n_4322),
.C(n_4540),
.Y(n_4992)
);

OAI21x1_ASAP7_75t_L g4993 ( 
.A1(n_4698),
.A2(n_4425),
.B(n_4397),
.Y(n_4993)
);

CKINVDCx20_ASAP7_75t_R g4994 ( 
.A(n_4638),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4860),
.B(n_4381),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4611),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4577),
.B(n_4401),
.Y(n_4997)
);

BUFx10_ASAP7_75t_L g4998 ( 
.A(n_4746),
.Y(n_4998)
);

AOI21xp5_ASAP7_75t_L g4999 ( 
.A1(n_4652),
.A2(n_4208),
.B(n_4410),
.Y(n_4999)
);

INVx1_ASAP7_75t_SL g5000 ( 
.A(n_4696),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4611),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4624),
.Y(n_5002)
);

A2O1A1Ixp33_ASAP7_75t_L g5003 ( 
.A1(n_4807),
.A2(n_4314),
.B(n_4525),
.C(n_4313),
.Y(n_5003)
);

HB1xp67_ASAP7_75t_L g5004 ( 
.A(n_4624),
.Y(n_5004)
);

BUFx2_ASAP7_75t_L g5005 ( 
.A(n_4593),
.Y(n_5005)
);

O2A1O1Ixp33_ASAP7_75t_L g5006 ( 
.A1(n_4809),
.A2(n_4528),
.B(n_4567),
.C(n_4531),
.Y(n_5006)
);

A2O1A1Ixp33_ASAP7_75t_L g5007 ( 
.A1(n_4615),
.A2(n_4948),
.B(n_4732),
.C(n_4652),
.Y(n_5007)
);

O2A1O1Ixp5_ASAP7_75t_L g5008 ( 
.A1(n_4766),
.A2(n_4483),
.B(n_4324),
.C(n_4272),
.Y(n_5008)
);

AOI21xp5_ASAP7_75t_L g5009 ( 
.A1(n_4785),
.A2(n_4267),
.B(n_4404),
.Y(n_5009)
);

AO31x2_ASAP7_75t_L g5010 ( 
.A1(n_4989),
.A2(n_4346),
.A3(n_4343),
.B(n_4339),
.Y(n_5010)
);

NOR2xp33_ASAP7_75t_L g5011 ( 
.A(n_4953),
.B(n_4406),
.Y(n_5011)
);

AO32x2_ASAP7_75t_L g5012 ( 
.A1(n_4610),
.A2(n_4317),
.A3(n_4545),
.B1(n_4350),
.B2(n_4290),
.Y(n_5012)
);

AOI221xp5_ASAP7_75t_L g5013 ( 
.A1(n_4877),
.A2(n_4378),
.B1(n_4436),
.B2(n_930),
.C(n_932),
.Y(n_5013)
);

CKINVDCx20_ASAP7_75t_R g5014 ( 
.A(n_4618),
.Y(n_5014)
);

AOI22xp33_ASAP7_75t_SL g5015 ( 
.A1(n_4606),
.A2(n_4458),
.B1(n_4533),
.B2(n_4317),
.Y(n_5015)
);

AOI21xp5_ASAP7_75t_L g5016 ( 
.A1(n_4785),
.A2(n_4726),
.B(n_4699),
.Y(n_5016)
);

BUFx2_ASAP7_75t_L g5017 ( 
.A(n_4593),
.Y(n_5017)
);

BUFx3_ASAP7_75t_L g5018 ( 
.A(n_4680),
.Y(n_5018)
);

O2A1O1Ixp33_ASAP7_75t_L g5019 ( 
.A1(n_4615),
.A2(n_4488),
.B(n_4429),
.C(n_1654),
.Y(n_5019)
);

AO21x1_ASAP7_75t_L g5020 ( 
.A1(n_4610),
.A2(n_4606),
.B(n_4573),
.Y(n_5020)
);

AOI21xp5_ASAP7_75t_L g5021 ( 
.A1(n_4726),
.A2(n_4473),
.B(n_4496),
.Y(n_5021)
);

INVxp67_ASAP7_75t_SL g5022 ( 
.A(n_4588),
.Y(n_5022)
);

OAI221xp5_ASAP7_75t_L g5023 ( 
.A1(n_4732),
.A2(n_934),
.B1(n_937),
.B2(n_927),
.C(n_921),
.Y(n_5023)
);

AND2x4_ASAP7_75t_L g5024 ( 
.A(n_4819),
.B(n_4533),
.Y(n_5024)
);

CKINVDCx5p33_ASAP7_75t_R g5025 ( 
.A(n_4578),
.Y(n_5025)
);

OAI21x1_ASAP7_75t_L g5026 ( 
.A1(n_4698),
.A2(n_4414),
.B(n_4428),
.Y(n_5026)
);

AOI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4699),
.A2(n_4506),
.B(n_4499),
.Y(n_5027)
);

NOR2xp33_ASAP7_75t_L g5028 ( 
.A(n_4960),
.B(n_4590),
.Y(n_5028)
);

INVx2_ASAP7_75t_L g5029 ( 
.A(n_4579),
.Y(n_5029)
);

CKINVDCx9p33_ASAP7_75t_R g5030 ( 
.A(n_4702),
.Y(n_5030)
);

NOR2xp33_ASAP7_75t_L g5031 ( 
.A(n_4740),
.B(n_4670),
.Y(n_5031)
);

AOI22xp33_ASAP7_75t_L g5032 ( 
.A1(n_4951),
.A2(n_4572),
.B1(n_4843),
.B2(n_4637),
.Y(n_5032)
);

AO31x2_ASAP7_75t_L g5033 ( 
.A1(n_4946),
.A2(n_4420),
.A3(n_4526),
.B(n_4517),
.Y(n_5033)
);

AOI22xp33_ASAP7_75t_L g5034 ( 
.A1(n_4572),
.A2(n_4545),
.B1(n_2493),
.B2(n_3304),
.Y(n_5034)
);

NAND3xp33_ASAP7_75t_SL g5035 ( 
.A(n_4874),
.B(n_940),
.C(n_939),
.Y(n_5035)
);

INVx2_ASAP7_75t_L g5036 ( 
.A(n_4594),
.Y(n_5036)
);

OAI21x1_ASAP7_75t_L g5037 ( 
.A1(n_4910),
.A2(n_4601),
.B(n_4787),
.Y(n_5037)
);

A2O1A1Ixp33_ASAP7_75t_L g5038 ( 
.A1(n_4582),
.A2(n_1534),
.B(n_1536),
.C(n_1533),
.Y(n_5038)
);

NAND3xp33_ASAP7_75t_L g5039 ( 
.A(n_4930),
.B(n_1538),
.C(n_1537),
.Y(n_5039)
);

OAI22xp5_ASAP7_75t_L g5040 ( 
.A1(n_4780),
.A2(n_4534),
.B1(n_4558),
.B2(n_4555),
.Y(n_5040)
);

AO31x2_ASAP7_75t_L g5041 ( 
.A1(n_4963),
.A2(n_4565),
.A3(n_4562),
.B(n_1369),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4571),
.Y(n_5042)
);

NOR2xp33_ASAP7_75t_L g5043 ( 
.A(n_4660),
.B(n_45),
.Y(n_5043)
);

A2O1A1Ixp33_ASAP7_75t_L g5044 ( 
.A1(n_4582),
.A2(n_1544),
.B(n_1545),
.C(n_1541),
.Y(n_5044)
);

OAI21x1_ASAP7_75t_L g5045 ( 
.A1(n_4910),
.A2(n_4561),
.B(n_4553),
.Y(n_5045)
);

O2A1O1Ixp33_ASAP7_75t_SL g5046 ( 
.A1(n_4695),
.A2(n_1657),
.B(n_1658),
.C(n_1653),
.Y(n_5046)
);

O2A1O1Ixp33_ASAP7_75t_SL g5047 ( 
.A1(n_4661),
.A2(n_1662),
.B(n_1664),
.C(n_1660),
.Y(n_5047)
);

OAI21xp5_ASAP7_75t_L g5048 ( 
.A1(n_4877),
.A2(n_1370),
.B(n_1369),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4580),
.Y(n_5049)
);

AND2x4_ASAP7_75t_L g5050 ( 
.A(n_4819),
.B(n_1370),
.Y(n_5050)
);

AOI21xp5_ASAP7_75t_L g5051 ( 
.A1(n_4776),
.A2(n_3063),
.B(n_3030),
.Y(n_5051)
);

HB1xp67_ASAP7_75t_L g5052 ( 
.A(n_4635),
.Y(n_5052)
);

AND2x2_ASAP7_75t_L g5053 ( 
.A(n_4616),
.B(n_1371),
.Y(n_5053)
);

OAI22xp33_ASAP7_75t_L g5054 ( 
.A1(n_4749),
.A2(n_3039),
.B1(n_3074),
.B2(n_3032),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4589),
.Y(n_5055)
);

NOR2xp33_ASAP7_75t_L g5056 ( 
.A(n_4597),
.B(n_4669),
.Y(n_5056)
);

AND2x2_ASAP7_75t_L g5057 ( 
.A(n_4719),
.B(n_1371),
.Y(n_5057)
);

OR2x2_ASAP7_75t_L g5058 ( 
.A(n_4639),
.B(n_1374),
.Y(n_5058)
);

OAI21xp5_ASAP7_75t_L g5059 ( 
.A1(n_4928),
.A2(n_1375),
.B(n_1374),
.Y(n_5059)
);

BUFx2_ASAP7_75t_L g5060 ( 
.A(n_4794),
.Y(n_5060)
);

A2O1A1Ixp33_ASAP7_75t_L g5061 ( 
.A1(n_4612),
.A2(n_1547),
.B(n_1551),
.C(n_1546),
.Y(n_5061)
);

A2O1A1Ixp33_ASAP7_75t_L g5062 ( 
.A1(n_4612),
.A2(n_1553),
.B(n_1554),
.C(n_1552),
.Y(n_5062)
);

AOI21xp5_ASAP7_75t_L g5063 ( 
.A1(n_4776),
.A2(n_4749),
.B(n_4601),
.Y(n_5063)
);

NOR2xp67_ASAP7_75t_SL g5064 ( 
.A(n_4708),
.B(n_3032),
.Y(n_5064)
);

BUFx2_ASAP7_75t_L g5065 ( 
.A(n_4811),
.Y(n_5065)
);

AOI21xp5_ASAP7_75t_L g5066 ( 
.A1(n_4687),
.A2(n_3063),
.B(n_3030),
.Y(n_5066)
);

AO21x2_ASAP7_75t_L g5067 ( 
.A1(n_4701),
.A2(n_1556),
.B(n_1555),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_4591),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_4604),
.Y(n_5069)
);

AOI21xp5_ASAP7_75t_L g5070 ( 
.A1(n_4958),
.A2(n_3063),
.B(n_3030),
.Y(n_5070)
);

OAI22xp33_ASAP7_75t_L g5071 ( 
.A1(n_4705),
.A2(n_3039),
.B1(n_3074),
.B2(n_3032),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4639),
.B(n_4635),
.Y(n_5072)
);

INVx2_ASAP7_75t_L g5073 ( 
.A(n_4614),
.Y(n_5073)
);

NAND2xp5_ASAP7_75t_L g5074 ( 
.A(n_4719),
.B(n_1375),
.Y(n_5074)
);

OR2x6_ASAP7_75t_L g5075 ( 
.A(n_4653),
.B(n_3032),
.Y(n_5075)
);

A2O1A1Ixp33_ASAP7_75t_L g5076 ( 
.A1(n_4608),
.A2(n_1559),
.B(n_1560),
.C(n_1557),
.Y(n_5076)
);

AO32x2_ASAP7_75t_L g5077 ( 
.A1(n_4982),
.A2(n_3315),
.A3(n_3345),
.B1(n_3284),
.B2(n_3274),
.Y(n_5077)
);

A2O1A1Ixp33_ASAP7_75t_L g5078 ( 
.A1(n_4835),
.A2(n_1562),
.B(n_1563),
.C(n_1561),
.Y(n_5078)
);

OAI21x1_ASAP7_75t_L g5079 ( 
.A1(n_4787),
.A2(n_3352),
.B(n_2676),
.Y(n_5079)
);

INVxp67_ASAP7_75t_L g5080 ( 
.A(n_4600),
.Y(n_5080)
);

AOI21xp5_ASAP7_75t_L g5081 ( 
.A1(n_4958),
.A2(n_3119),
.B(n_3101),
.Y(n_5081)
);

O2A1O1Ixp33_ASAP7_75t_L g5082 ( 
.A1(n_4935),
.A2(n_1666),
.B(n_1667),
.C(n_1665),
.Y(n_5082)
);

OR2x2_ASAP7_75t_L g5083 ( 
.A(n_4583),
.B(n_1376),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4613),
.Y(n_5084)
);

INVx2_ASAP7_75t_L g5085 ( 
.A(n_4626),
.Y(n_5085)
);

NAND2x1_ASAP7_75t_L g5086 ( 
.A(n_4913),
.B(n_4596),
.Y(n_5086)
);

AOI21xp5_ASAP7_75t_L g5087 ( 
.A1(n_4981),
.A2(n_3119),
.B(n_3101),
.Y(n_5087)
);

BUFx6f_ASAP7_75t_L g5088 ( 
.A(n_4629),
.Y(n_5088)
);

OAI21x1_ASAP7_75t_L g5089 ( 
.A1(n_4712),
.A2(n_3352),
.B(n_2676),
.Y(n_5089)
);

A2O1A1Ixp33_ASAP7_75t_L g5090 ( 
.A1(n_4835),
.A2(n_1568),
.B(n_1567),
.C(n_1377),
.Y(n_5090)
);

AO31x2_ASAP7_75t_L g5091 ( 
.A1(n_4929),
.A2(n_1376),
.A3(n_1378),
.B(n_1377),
.Y(n_5091)
);

OAI22xp5_ASAP7_75t_L g5092 ( 
.A1(n_4983),
.A2(n_4857),
.B1(n_4764),
.B2(n_4678),
.Y(n_5092)
);

INVx4_ASAP7_75t_L g5093 ( 
.A(n_4682),
.Y(n_5093)
);

OAI22xp5_ASAP7_75t_L g5094 ( 
.A1(n_4857),
.A2(n_3166),
.B1(n_3074),
.B2(n_3084),
.Y(n_5094)
);

AND2x4_ASAP7_75t_L g5095 ( 
.A(n_4819),
.B(n_1378),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4981),
.A2(n_4588),
.B(n_4688),
.Y(n_5096)
);

BUFx6f_ASAP7_75t_L g5097 ( 
.A(n_4629),
.Y(n_5097)
);

AOI21xp5_ASAP7_75t_SL g5098 ( 
.A1(n_4684),
.A2(n_3119),
.B(n_3101),
.Y(n_5098)
);

INVx2_ASAP7_75t_L g5099 ( 
.A(n_4628),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4640),
.Y(n_5100)
);

AOI21xp5_ASAP7_75t_L g5101 ( 
.A1(n_4688),
.A2(n_3135),
.B(n_3130),
.Y(n_5101)
);

OAI21xp5_ASAP7_75t_L g5102 ( 
.A1(n_4928),
.A2(n_1384),
.B(n_1380),
.Y(n_5102)
);

HB1xp67_ASAP7_75t_L g5103 ( 
.A(n_4584),
.Y(n_5103)
);

AOI21xp5_ASAP7_75t_L g5104 ( 
.A1(n_4823),
.A2(n_3135),
.B(n_3130),
.Y(n_5104)
);

CKINVDCx5p33_ASAP7_75t_R g5105 ( 
.A(n_4585),
.Y(n_5105)
);

NOR2xp33_ASAP7_75t_L g5106 ( 
.A(n_4665),
.B(n_4829),
.Y(n_5106)
);

AOI22xp5_ASAP7_75t_L g5107 ( 
.A1(n_4764),
.A2(n_941),
.B1(n_944),
.B2(n_943),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4646),
.Y(n_5108)
);

OAI21x1_ASAP7_75t_SL g5109 ( 
.A1(n_4573),
.A2(n_1669),
.B(n_1668),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4648),
.Y(n_5110)
);

BUFx2_ASAP7_75t_L g5111 ( 
.A(n_4656),
.Y(n_5111)
);

OAI222xp33_ASAP7_75t_L g5112 ( 
.A1(n_4620),
.A2(n_1391),
.B1(n_1384),
.B2(n_1393),
.C1(n_1390),
.C2(n_1380),
.Y(n_5112)
);

A2O1A1Ixp33_ASAP7_75t_L g5113 ( 
.A1(n_4952),
.A2(n_1391),
.B(n_1393),
.C(n_1390),
.Y(n_5113)
);

OR2x2_ASAP7_75t_L g5114 ( 
.A(n_4621),
.B(n_1394),
.Y(n_5114)
);

AND2x6_ASAP7_75t_SL g5115 ( 
.A(n_4707),
.B(n_1670),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4649),
.Y(n_5116)
);

AOI21xp5_ASAP7_75t_L g5117 ( 
.A1(n_4823),
.A2(n_3135),
.B(n_3130),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4654),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_L g5119 ( 
.A(n_4850),
.B(n_1394),
.Y(n_5119)
);

NOR2xp33_ASAP7_75t_SL g5120 ( 
.A(n_4737),
.B(n_3345),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_4655),
.Y(n_5121)
);

AND2x6_ASAP7_75t_L g5122 ( 
.A(n_4713),
.B(n_3039),
.Y(n_5122)
);

OAI21xp5_ASAP7_75t_L g5123 ( 
.A1(n_4952),
.A2(n_1397),
.B(n_1396),
.Y(n_5123)
);

BUFx3_ASAP7_75t_L g5124 ( 
.A(n_4605),
.Y(n_5124)
);

AOI22xp5_ASAP7_75t_L g5125 ( 
.A1(n_4971),
.A2(n_946),
.B1(n_948),
.B2(n_947),
.Y(n_5125)
);

O2A1O1Ixp33_ASAP7_75t_SL g5126 ( 
.A1(n_4627),
.A2(n_1673),
.B(n_47),
.C(n_48),
.Y(n_5126)
);

AND2x2_ASAP7_75t_L g5127 ( 
.A(n_4609),
.B(n_1396),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_4658),
.Y(n_5128)
);

A2O1A1Ixp33_ASAP7_75t_L g5129 ( 
.A1(n_4971),
.A2(n_1472),
.B(n_1397),
.C(n_949),
.Y(n_5129)
);

O2A1O1Ixp33_ASAP7_75t_L g5130 ( 
.A1(n_4935),
.A2(n_4581),
.B(n_4622),
.C(n_4965),
.Y(n_5130)
);

OAI22xp5_ASAP7_75t_L g5131 ( 
.A1(n_4636),
.A2(n_3166),
.B1(n_3074),
.B2(n_3084),
.Y(n_5131)
);

AOI21xp5_ASAP7_75t_L g5132 ( 
.A1(n_4771),
.A2(n_4800),
.B(n_4918),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_4633),
.B(n_1472),
.Y(n_5133)
);

AO31x2_ASAP7_75t_L g5134 ( 
.A1(n_4933),
.A2(n_3304),
.A3(n_3305),
.B(n_3303),
.Y(n_5134)
);

AND2x4_ASAP7_75t_L g5135 ( 
.A(n_4819),
.B(n_2948),
.Y(n_5135)
);

AOI221xp5_ASAP7_75t_L g5136 ( 
.A1(n_4880),
.A2(n_952),
.B1(n_955),
.B2(n_953),
.C(n_950),
.Y(n_5136)
);

OAI22x1_ASAP7_75t_L g5137 ( 
.A1(n_4921),
.A2(n_4842),
.B1(n_4961),
.B2(n_4690),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4662),
.Y(n_5138)
);

A2O1A1Ixp33_ASAP7_75t_L g5139 ( 
.A1(n_4716),
.A2(n_957),
.B(n_960),
.C(n_958),
.Y(n_5139)
);

BUFx3_ASAP7_75t_L g5140 ( 
.A(n_4617),
.Y(n_5140)
);

INVx1_ASAP7_75t_SL g5141 ( 
.A(n_4727),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_4723),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_L g5143 ( 
.A(n_4850),
.B(n_4),
.Y(n_5143)
);

OAI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_4921),
.A2(n_3084),
.B1(n_3086),
.B2(n_3039),
.Y(n_5144)
);

BUFx2_ASAP7_75t_L g5145 ( 
.A(n_4692),
.Y(n_5145)
);

NOR2xp33_ASAP7_75t_L g5146 ( 
.A(n_4665),
.B(n_4728),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_4621),
.B(n_5),
.Y(n_5147)
);

NOR2xp33_ASAP7_75t_L g5148 ( 
.A(n_4665),
.B(n_46),
.Y(n_5148)
);

CKINVDCx20_ASAP7_75t_R g5149 ( 
.A(n_4814),
.Y(n_5149)
);

A2O1A1Ixp33_ASAP7_75t_L g5150 ( 
.A1(n_4898),
.A2(n_959),
.B(n_964),
.C(n_963),
.Y(n_5150)
);

OAI22xp5_ASAP7_75t_L g5151 ( 
.A1(n_4921),
.A2(n_3086),
.B1(n_3096),
.B2(n_3084),
.Y(n_5151)
);

AOI22xp33_ASAP7_75t_L g5152 ( 
.A1(n_4603),
.A2(n_3387),
.B1(n_3392),
.B2(n_3382),
.Y(n_5152)
);

OAI21xp5_ASAP7_75t_L g5153 ( 
.A1(n_4912),
.A2(n_971),
.B(n_970),
.Y(n_5153)
);

A2O1A1Ixp33_ASAP7_75t_L g5154 ( 
.A1(n_4895),
.A2(n_972),
.B(n_975),
.C(n_973),
.Y(n_5154)
);

NAND3xp33_ASAP7_75t_L g5155 ( 
.A(n_4587),
.B(n_978),
.C(n_976),
.Y(n_5155)
);

O2A1O1Ixp33_ASAP7_75t_L g5156 ( 
.A1(n_4821),
.A2(n_938),
.B(n_3225),
.C(n_3190),
.Y(n_5156)
);

AOI21xp5_ASAP7_75t_L g5157 ( 
.A1(n_4771),
.A2(n_3096),
.B(n_3086),
.Y(n_5157)
);

O2A1O1Ixp5_ASAP7_75t_L g5158 ( 
.A1(n_4956),
.A2(n_2380),
.B(n_2384),
.C(n_2370),
.Y(n_5158)
);

A2O1A1Ixp33_ASAP7_75t_L g5159 ( 
.A1(n_4895),
.A2(n_981),
.B(n_983),
.C(n_979),
.Y(n_5159)
);

NOR2xp33_ASAP7_75t_SL g5160 ( 
.A(n_4752),
.B(n_3345),
.Y(n_5160)
);

OAI22xp33_ASAP7_75t_L g5161 ( 
.A1(n_4921),
.A2(n_3096),
.B1(n_3100),
.B2(n_3086),
.Y(n_5161)
);

CKINVDCx5p33_ASAP7_75t_R g5162 ( 
.A(n_4647),
.Y(n_5162)
);

BUFx2_ASAP7_75t_L g5163 ( 
.A(n_4694),
.Y(n_5163)
);

OAI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_4985),
.A2(n_994),
.B(n_987),
.Y(n_5164)
);

AOI221x1_ASAP7_75t_L g5165 ( 
.A1(n_4664),
.A2(n_1936),
.B1(n_3370),
.B2(n_3375),
.C(n_3367),
.Y(n_5165)
);

O2A1O1Ixp33_ASAP7_75t_L g5166 ( 
.A1(n_4974),
.A2(n_2380),
.B(n_2384),
.C(n_2370),
.Y(n_5166)
);

CKINVDCx20_ASAP7_75t_R g5167 ( 
.A(n_4791),
.Y(n_5167)
);

OAI221xp5_ASAP7_75t_L g5168 ( 
.A1(n_4641),
.A2(n_4631),
.B1(n_4959),
.B2(n_4889),
.C(n_4936),
.Y(n_5168)
);

OA21x2_ASAP7_75t_L g5169 ( 
.A1(n_4934),
.A2(n_2079),
.B(n_2077),
.Y(n_5169)
);

A2O1A1Ixp33_ASAP7_75t_L g5170 ( 
.A1(n_4974),
.A2(n_997),
.B(n_1002),
.C(n_995),
.Y(n_5170)
);

NOR2xp67_ASAP7_75t_L g5171 ( 
.A(n_4982),
.B(n_47),
.Y(n_5171)
);

AOI21xp5_ASAP7_75t_L g5172 ( 
.A1(n_4800),
.A2(n_3100),
.B(n_3096),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_4765),
.B(n_5),
.Y(n_5173)
);

AOI22xp33_ASAP7_75t_SL g5174 ( 
.A1(n_4909),
.A2(n_1008),
.B1(n_1010),
.B2(n_1005),
.Y(n_5174)
);

CKINVDCx5p33_ASAP7_75t_R g5175 ( 
.A(n_4739),
.Y(n_5175)
);

INVx2_ASAP7_75t_L g5176 ( 
.A(n_4645),
.Y(n_5176)
);

A2O1A1Ixp33_ASAP7_75t_L g5177 ( 
.A1(n_4925),
.A2(n_1013),
.B(n_1015),
.C(n_1012),
.Y(n_5177)
);

AOI21xp5_ASAP7_75t_L g5178 ( 
.A1(n_4587),
.A2(n_3134),
.B(n_3100),
.Y(n_5178)
);

BUFx6f_ASAP7_75t_L g5179 ( 
.A(n_4629),
.Y(n_5179)
);

BUFx3_ASAP7_75t_L g5180 ( 
.A(n_4738),
.Y(n_5180)
);

NAND2x1p5_ASAP7_75t_L g5181 ( 
.A(n_4710),
.B(n_4715),
.Y(n_5181)
);

BUFx10_ASAP7_75t_L g5182 ( 
.A(n_4644),
.Y(n_5182)
);

NAND2xp5_ASAP7_75t_SL g5183 ( 
.A(n_4748),
.B(n_3100),
.Y(n_5183)
);

INVx2_ASAP7_75t_SL g5184 ( 
.A(n_4844),
.Y(n_5184)
);

AOI21xp5_ASAP7_75t_L g5185 ( 
.A1(n_4684),
.A2(n_3144),
.B(n_3134),
.Y(n_5185)
);

O2A1O1Ixp33_ASAP7_75t_SL g5186 ( 
.A1(n_4897),
.A2(n_51),
.B(n_53),
.C(n_49),
.Y(n_5186)
);

A2O1A1Ixp33_ASAP7_75t_L g5187 ( 
.A1(n_4972),
.A2(n_1019),
.B(n_1027),
.C(n_1016),
.Y(n_5187)
);

NOR2xp33_ASAP7_75t_L g5188 ( 
.A(n_4791),
.B(n_49),
.Y(n_5188)
);

AOI22xp33_ASAP7_75t_L g5189 ( 
.A1(n_4840),
.A2(n_4881),
.B1(n_4882),
.B2(n_4883),
.Y(n_5189)
);

OR2x2_ASAP7_75t_L g5190 ( 
.A(n_4765),
.B(n_5),
.Y(n_5190)
);

INVx2_ASAP7_75t_L g5191 ( 
.A(n_4650),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4729),
.Y(n_5192)
);

AOI22xp5_ASAP7_75t_L g5193 ( 
.A1(n_4721),
.A2(n_1031),
.B1(n_1034),
.B2(n_1030),
.Y(n_5193)
);

AOI21xp5_ASAP7_75t_L g5194 ( 
.A1(n_4709),
.A2(n_3144),
.B(n_3134),
.Y(n_5194)
);

OAI22xp5_ASAP7_75t_L g5195 ( 
.A1(n_4979),
.A2(n_3144),
.B1(n_3175),
.B2(n_3134),
.Y(n_5195)
);

AOI21xp5_ASAP7_75t_L g5196 ( 
.A1(n_4709),
.A2(n_3175),
.B(n_3144),
.Y(n_5196)
);

OAI21xp5_ASAP7_75t_L g5197 ( 
.A1(n_4987),
.A2(n_1036),
.B(n_1035),
.Y(n_5197)
);

AOI21xp5_ASAP7_75t_L g5198 ( 
.A1(n_4955),
.A2(n_3198),
.B(n_3175),
.Y(n_5198)
);

OR2x2_ASAP7_75t_L g5199 ( 
.A(n_4862),
.B(n_6),
.Y(n_5199)
);

AO21x1_ASAP7_75t_L g5200 ( 
.A1(n_4810),
.A2(n_6),
.B(n_7),
.Y(n_5200)
);

OAI21x1_ASAP7_75t_L g5201 ( 
.A1(n_4944),
.A2(n_2736),
.B(n_2630),
.Y(n_5201)
);

O2A1O1Ixp33_ASAP7_75t_L g5202 ( 
.A1(n_4721),
.A2(n_2409),
.B(n_2410),
.C(n_2388),
.Y(n_5202)
);

O2A1O1Ixp33_ASAP7_75t_SL g5203 ( 
.A1(n_4926),
.A2(n_55),
.B(n_56),
.C(n_53),
.Y(n_5203)
);

BUFx6f_ASAP7_75t_SL g5204 ( 
.A(n_4644),
.Y(n_5204)
);

NOR2xp33_ASAP7_75t_L g5205 ( 
.A(n_4630),
.B(n_4941),
.Y(n_5205)
);

A2O1A1Ixp33_ASAP7_75t_L g5206 ( 
.A1(n_4979),
.A2(n_1043),
.B(n_1044),
.C(n_1040),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_4663),
.Y(n_5207)
);

NAND3xp33_ASAP7_75t_L g5208 ( 
.A(n_4885),
.B(n_1050),
.C(n_1048),
.Y(n_5208)
);

INVx2_ASAP7_75t_SL g5209 ( 
.A(n_4704),
.Y(n_5209)
);

OR2x2_ASAP7_75t_L g5210 ( 
.A(n_4862),
.B(n_7),
.Y(n_5210)
);

AOI21xp5_ASAP7_75t_L g5211 ( 
.A1(n_4973),
.A2(n_3198),
.B(n_3175),
.Y(n_5211)
);

INVx2_ASAP7_75t_L g5212 ( 
.A(n_4667),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_4671),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_4672),
.Y(n_5214)
);

AOI21xp5_ASAP7_75t_L g5215 ( 
.A1(n_4977),
.A2(n_3227),
.B(n_3198),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_4742),
.Y(n_5216)
);

AND2x2_ASAP7_75t_L g5217 ( 
.A(n_4722),
.B(n_7),
.Y(n_5217)
);

HB1xp67_ASAP7_75t_L g5218 ( 
.A(n_4697),
.Y(n_5218)
);

OAI21xp5_ASAP7_75t_L g5219 ( 
.A1(n_4689),
.A2(n_1053),
.B(n_1052),
.Y(n_5219)
);

AOI22xp33_ASAP7_75t_L g5220 ( 
.A1(n_4724),
.A2(n_4911),
.B1(n_4914),
.B2(n_4770),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_4810),
.B(n_8),
.Y(n_5221)
);

AO31x2_ASAP7_75t_L g5222 ( 
.A1(n_4975),
.A2(n_3305),
.A3(n_3336),
.B(n_3303),
.Y(n_5222)
);

OAI21x1_ASAP7_75t_L g5223 ( 
.A1(n_4944),
.A2(n_2736),
.B(n_2630),
.Y(n_5223)
);

O2A1O1Ixp33_ASAP7_75t_L g5224 ( 
.A1(n_4872),
.A2(n_2409),
.B(n_2410),
.C(n_2388),
.Y(n_5224)
);

A2O1A1Ixp33_ASAP7_75t_L g5225 ( 
.A1(n_4916),
.A2(n_1058),
.B(n_1059),
.C(n_1056),
.Y(n_5225)
);

O2A1O1Ixp33_ASAP7_75t_L g5226 ( 
.A1(n_4873),
.A2(n_2337),
.B(n_2338),
.C(n_2329),
.Y(n_5226)
);

AO21x1_ASAP7_75t_L g5227 ( 
.A1(n_4689),
.A2(n_8),
.B(n_9),
.Y(n_5227)
);

NOR2xp33_ASAP7_75t_L g5228 ( 
.A(n_4586),
.B(n_57),
.Y(n_5228)
);

OAI21x1_ASAP7_75t_L g5229 ( 
.A1(n_4834),
.A2(n_3343),
.B(n_3336),
.Y(n_5229)
);

AOI22xp5_ASAP7_75t_L g5230 ( 
.A1(n_4831),
.A2(n_1063),
.B1(n_1067),
.B2(n_1062),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_4681),
.B(n_9),
.Y(n_5231)
);

AO32x2_ASAP7_75t_L g5232 ( 
.A1(n_4956),
.A2(n_12),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_5232)
);

HB1xp67_ASAP7_75t_L g5233 ( 
.A(n_4697),
.Y(n_5233)
);

NOR2x1_ASAP7_75t_SL g5234 ( 
.A(n_4653),
.B(n_3198),
.Y(n_5234)
);

AND2x4_ASAP7_75t_L g5235 ( 
.A(n_4653),
.B(n_4713),
.Y(n_5235)
);

A2O1A1Ixp33_ASAP7_75t_L g5236 ( 
.A1(n_4916),
.A2(n_1069),
.B(n_1075),
.C(n_1074),
.Y(n_5236)
);

AOI21xp5_ASAP7_75t_L g5237 ( 
.A1(n_4978),
.A2(n_3228),
.B(n_3227),
.Y(n_5237)
);

INVxp67_ASAP7_75t_SL g5238 ( 
.A(n_4927),
.Y(n_5238)
);

A2O1A1Ixp33_ASAP7_75t_L g5239 ( 
.A1(n_4980),
.A2(n_1077),
.B(n_1082),
.C(n_1078),
.Y(n_5239)
);

CKINVDCx5p33_ASAP7_75t_R g5240 ( 
.A(n_4762),
.Y(n_5240)
);

HB1xp67_ASAP7_75t_L g5241 ( 
.A(n_4711),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_4757),
.Y(n_5242)
);

OAI22xp5_ASAP7_75t_L g5243 ( 
.A1(n_4710),
.A2(n_3228),
.B1(n_3237),
.B2(n_3227),
.Y(n_5243)
);

OAI21x1_ASAP7_75t_L g5244 ( 
.A1(n_4834),
.A2(n_3344),
.B(n_3343),
.Y(n_5244)
);

INVx1_ASAP7_75t_SL g5245 ( 
.A(n_4893),
.Y(n_5245)
);

AND2x4_ASAP7_75t_SL g5246 ( 
.A(n_4644),
.B(n_3227),
.Y(n_5246)
);

O2A1O1Ixp33_ASAP7_75t_L g5247 ( 
.A1(n_4964),
.A2(n_2337),
.B(n_2338),
.C(n_2329),
.Y(n_5247)
);

OA21x2_ASAP7_75t_L g5248 ( 
.A1(n_4923),
.A2(n_2079),
.B(n_2077),
.Y(n_5248)
);

OAI22xp5_ASAP7_75t_L g5249 ( 
.A1(n_4715),
.A2(n_3237),
.B1(n_3240),
.B2(n_3228),
.Y(n_5249)
);

A2O1A1Ixp33_ASAP7_75t_L g5250 ( 
.A1(n_4824),
.A2(n_1083),
.B(n_1086),
.C(n_1084),
.Y(n_5250)
);

A2O1A1Ixp33_ASAP7_75t_L g5251 ( 
.A1(n_4824),
.A2(n_1088),
.B(n_1092),
.C(n_1091),
.Y(n_5251)
);

OAI21xp5_ASAP7_75t_L g5252 ( 
.A1(n_4837),
.A2(n_1096),
.B(n_1068),
.Y(n_5252)
);

O2A1O1Ixp33_ASAP7_75t_SL g5253 ( 
.A1(n_4781),
.A2(n_59),
.B(n_61),
.C(n_57),
.Y(n_5253)
);

A2O1A1Ixp33_ASAP7_75t_L g5254 ( 
.A1(n_4837),
.A2(n_1103),
.B(n_1106),
.C(n_1097),
.Y(n_5254)
);

A2O1A1Ixp33_ASAP7_75t_L g5255 ( 
.A1(n_4920),
.A2(n_1107),
.B(n_1115),
.C(n_1105),
.Y(n_5255)
);

AOI21xp5_ASAP7_75t_L g5256 ( 
.A1(n_4988),
.A2(n_4768),
.B(n_4957),
.Y(n_5256)
);

INVx2_ASAP7_75t_L g5257 ( 
.A(n_4673),
.Y(n_5257)
);

INVx2_ASAP7_75t_SL g5258 ( 
.A(n_4861),
.Y(n_5258)
);

AOI22xp5_ASAP7_75t_L g5259 ( 
.A1(n_4677),
.A2(n_1120),
.B1(n_1121),
.B2(n_1108),
.Y(n_5259)
);

AOI21xp33_ASAP7_75t_L g5260 ( 
.A1(n_4942),
.A2(n_3355),
.B(n_3344),
.Y(n_5260)
);

AO31x2_ASAP7_75t_L g5261 ( 
.A1(n_4945),
.A2(n_3355),
.A3(n_2495),
.B(n_2496),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_4758),
.Y(n_5262)
);

AOI21xp33_ASAP7_75t_L g5263 ( 
.A1(n_4867),
.A2(n_1123),
.B(n_1122),
.Y(n_5263)
);

O2A1O1Ixp33_ASAP7_75t_L g5264 ( 
.A1(n_4675),
.A2(n_2343),
.B(n_2344),
.C(n_2342),
.Y(n_5264)
);

O2A1O1Ixp33_ASAP7_75t_L g5265 ( 
.A1(n_4927),
.A2(n_2343),
.B(n_2344),
.C(n_2342),
.Y(n_5265)
);

AOI22xp33_ASAP7_75t_L g5266 ( 
.A1(n_4651),
.A2(n_2490),
.B1(n_2496),
.B2(n_2495),
.Y(n_5266)
);

OAI21xp5_ASAP7_75t_L g5267 ( 
.A1(n_4938),
.A2(n_1130),
.B(n_1128),
.Y(n_5267)
);

AOI22xp33_ASAP7_75t_L g5268 ( 
.A1(n_4884),
.A2(n_2490),
.B1(n_2516),
.B2(n_2514),
.Y(n_5268)
);

INVx2_ASAP7_75t_L g5269 ( 
.A(n_4706),
.Y(n_5269)
);

AOI21xp5_ASAP7_75t_L g5270 ( 
.A1(n_4768),
.A2(n_3237),
.B(n_3228),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_L g5271 ( 
.A(n_4681),
.B(n_10),
.Y(n_5271)
);

OAI21xp5_ASAP7_75t_L g5272 ( 
.A1(n_4938),
.A2(n_1137),
.B(n_1131),
.Y(n_5272)
);

NOR2xp33_ASAP7_75t_SL g5273 ( 
.A(n_4767),
.B(n_3237),
.Y(n_5273)
);

BUFx3_ASAP7_75t_L g5274 ( 
.A(n_4775),
.Y(n_5274)
);

O2A1O1Ixp33_ASAP7_75t_L g5275 ( 
.A1(n_4943),
.A2(n_2346),
.B(n_2349),
.C(n_2345),
.Y(n_5275)
);

BUFx2_ASAP7_75t_L g5276 ( 
.A(n_4685),
.Y(n_5276)
);

OAI21x1_ASAP7_75t_L g5277 ( 
.A1(n_4962),
.A2(n_3332),
.B(n_2070),
.Y(n_5277)
);

INVx3_ASAP7_75t_L g5278 ( 
.A(n_4596),
.Y(n_5278)
);

AOI21xp5_ASAP7_75t_L g5279 ( 
.A1(n_4768),
.A2(n_3249),
.B(n_3240),
.Y(n_5279)
);

A2O1A1Ixp33_ASAP7_75t_L g5280 ( 
.A1(n_4920),
.A2(n_1140),
.B(n_1142),
.C(n_1139),
.Y(n_5280)
);

INVx3_ASAP7_75t_L g5281 ( 
.A(n_4599),
.Y(n_5281)
);

AO21x2_ASAP7_75t_L g5282 ( 
.A1(n_4701),
.A2(n_2516),
.B(n_2514),
.Y(n_5282)
);

BUFx2_ASAP7_75t_L g5283 ( 
.A(n_4685),
.Y(n_5283)
);

NOR2xp33_ASAP7_75t_L g5284 ( 
.A(n_4586),
.B(n_61),
.Y(n_5284)
);

CKINVDCx20_ASAP7_75t_R g5285 ( 
.A(n_4753),
.Y(n_5285)
);

NAND2xp5_ASAP7_75t_L g5286 ( 
.A(n_4827),
.B(n_10),
.Y(n_5286)
);

O2A1O1Ixp33_ASAP7_75t_SL g5287 ( 
.A1(n_4781),
.A2(n_63),
.B(n_64),
.C(n_62),
.Y(n_5287)
);

INVx1_ASAP7_75t_L g5288 ( 
.A(n_4772),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_4778),
.Y(n_5289)
);

AND2x4_ASAP7_75t_L g5290 ( 
.A(n_4733),
.B(n_2948),
.Y(n_5290)
);

AOI22xp5_ASAP7_75t_L g5291 ( 
.A1(n_4932),
.A2(n_1143),
.B1(n_1147),
.B2(n_1141),
.Y(n_5291)
);

NOR2xp33_ASAP7_75t_L g5292 ( 
.A(n_4595),
.B(n_62),
.Y(n_5292)
);

INVx2_ASAP7_75t_L g5293 ( 
.A(n_4725),
.Y(n_5293)
);

OAI22xp5_ASAP7_75t_L g5294 ( 
.A1(n_4932),
.A2(n_3249),
.B1(n_3269),
.B2(n_3240),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_4786),
.Y(n_5295)
);

A2O1A1Ixp33_ASAP7_75t_L g5296 ( 
.A1(n_4947),
.A2(n_1151),
.B(n_1155),
.C(n_1150),
.Y(n_5296)
);

OR2x6_ASAP7_75t_L g5297 ( 
.A(n_4575),
.B(n_3240),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4799),
.Y(n_5298)
);

NAND2xp5_ASAP7_75t_L g5299 ( 
.A(n_4754),
.B(n_11),
.Y(n_5299)
);

OA21x2_ASAP7_75t_L g5300 ( 
.A1(n_4864),
.A2(n_2070),
.B(n_2520),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_4803),
.Y(n_5301)
);

INVx4_ASAP7_75t_L g5302 ( 
.A(n_4682),
.Y(n_5302)
);

AOI22xp5_ASAP7_75t_L g5303 ( 
.A1(n_4947),
.A2(n_1160),
.B1(n_1161),
.B2(n_1159),
.Y(n_5303)
);

OAI21x1_ASAP7_75t_L g5304 ( 
.A1(n_4602),
.A2(n_3332),
.B(n_2523),
.Y(n_5304)
);

BUFx10_ASAP7_75t_L g5305 ( 
.A(n_4657),
.Y(n_5305)
);

A2O1A1Ixp33_ASAP7_75t_L g5306 ( 
.A1(n_4763),
.A2(n_1164),
.B(n_1166),
.C(n_1162),
.Y(n_5306)
);

NAND2xp5_ASAP7_75t_L g5307 ( 
.A(n_4754),
.B(n_12),
.Y(n_5307)
);

O2A1O1Ixp33_ASAP7_75t_SL g5308 ( 
.A1(n_4792),
.A2(n_64),
.B(n_65),
.C(n_63),
.Y(n_5308)
);

BUFx6f_ASAP7_75t_L g5309 ( 
.A(n_4657),
.Y(n_5309)
);

CKINVDCx11_ASAP7_75t_R g5310 ( 
.A(n_4826),
.Y(n_5310)
);

AO31x2_ASAP7_75t_L g5311 ( 
.A1(n_4902),
.A2(n_2523),
.A3(n_2533),
.B(n_2520),
.Y(n_5311)
);

OAI21xp5_ASAP7_75t_L g5312 ( 
.A1(n_4949),
.A2(n_1168),
.B(n_1167),
.Y(n_5312)
);

OAI22xp5_ASAP7_75t_L g5313 ( 
.A1(n_4760),
.A2(n_3269),
.B1(n_3280),
.B2(n_3249),
.Y(n_5313)
);

O2A1O1Ixp33_ASAP7_75t_SL g5314 ( 
.A1(n_4792),
.A2(n_4642),
.B(n_4750),
.C(n_4777),
.Y(n_5314)
);

O2A1O1Ixp33_ASAP7_75t_L g5315 ( 
.A1(n_4939),
.A2(n_4642),
.B(n_4864),
.C(n_4902),
.Y(n_5315)
);

NAND2xp5_ASAP7_75t_SL g5316 ( 
.A(n_4851),
.B(n_3249),
.Y(n_5316)
);

INVx1_ASAP7_75t_SL g5317 ( 
.A(n_4782),
.Y(n_5317)
);

AO31x2_ASAP7_75t_L g5318 ( 
.A1(n_4908),
.A2(n_4919),
.A3(n_4868),
.B(n_4731),
.Y(n_5318)
);

OAI21x1_ASAP7_75t_L g5319 ( 
.A1(n_4602),
.A2(n_2537),
.B(n_2533),
.Y(n_5319)
);

AOI221xp5_ASAP7_75t_SL g5320 ( 
.A1(n_4858),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.C(n_16),
.Y(n_5320)
);

NAND2x1_ASAP7_75t_L g5321 ( 
.A(n_4599),
.B(n_3269),
.Y(n_5321)
);

OR2x2_ASAP7_75t_L g5322 ( 
.A(n_4666),
.B(n_13),
.Y(n_5322)
);

OAI21x1_ASAP7_75t_L g5323 ( 
.A1(n_4619),
.A2(n_2540),
.B(n_2537),
.Y(n_5323)
);

AOI21xp5_ASAP7_75t_L g5324 ( 
.A1(n_4957),
.A2(n_3280),
.B(n_3269),
.Y(n_5324)
);

BUFx10_ASAP7_75t_L g5325 ( 
.A(n_4657),
.Y(n_5325)
);

INVx2_ASAP7_75t_SL g5326 ( 
.A(n_4879),
.Y(n_5326)
);

NOR2xp33_ASAP7_75t_L g5327 ( 
.A(n_4595),
.B(n_65),
.Y(n_5327)
);

AO31x2_ASAP7_75t_L g5328 ( 
.A1(n_4868),
.A2(n_2547),
.A3(n_2548),
.B(n_2540),
.Y(n_5328)
);

O2A1O1Ixp33_ASAP7_75t_L g5329 ( 
.A1(n_4858),
.A2(n_2346),
.B(n_2349),
.C(n_2345),
.Y(n_5329)
);

NAND2xp5_ASAP7_75t_L g5330 ( 
.A(n_4759),
.B(n_15),
.Y(n_5330)
);

OAI21x1_ASAP7_75t_L g5331 ( 
.A1(n_4619),
.A2(n_2548),
.B(n_2547),
.Y(n_5331)
);

A2O1A1Ixp33_ASAP7_75t_L g5332 ( 
.A1(n_4867),
.A2(n_4878),
.B(n_4679),
.C(n_4853),
.Y(n_5332)
);

INVx2_ASAP7_75t_L g5333 ( 
.A(n_4730),
.Y(n_5333)
);

AOI21xp5_ASAP7_75t_L g5334 ( 
.A1(n_4957),
.A2(n_3334),
.B(n_3280),
.Y(n_5334)
);

AOI21xp5_ASAP7_75t_L g5335 ( 
.A1(n_4755),
.A2(n_3334),
.B(n_3280),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_4759),
.B(n_16),
.Y(n_5336)
);

AOI21xp33_ASAP7_75t_L g5337 ( 
.A1(n_4878),
.A2(n_1178),
.B(n_1170),
.Y(n_5337)
);

OAI21x1_ASAP7_75t_L g5338 ( 
.A1(n_4718),
.A2(n_2550),
.B(n_2549),
.Y(n_5338)
);

CKINVDCx20_ASAP7_75t_R g5339 ( 
.A(n_4761),
.Y(n_5339)
);

AO22x1_ASAP7_75t_L g5340 ( 
.A1(n_4733),
.A2(n_1183),
.B1(n_1184),
.B2(n_1182),
.Y(n_5340)
);

AOI22xp33_ASAP7_75t_SL g5341 ( 
.A1(n_4747),
.A2(n_1191),
.B1(n_1195),
.B2(n_1185),
.Y(n_5341)
);

AOI21xp5_ASAP7_75t_L g5342 ( 
.A1(n_4575),
.A2(n_3353),
.B(n_3334),
.Y(n_5342)
);

O2A1O1Ixp33_ASAP7_75t_L g5343 ( 
.A1(n_4666),
.A2(n_2355),
.B(n_2358),
.C(n_2353),
.Y(n_5343)
);

AO32x2_ASAP7_75t_L g5344 ( 
.A1(n_4966),
.A2(n_19),
.A3(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_5344)
);

AND2x2_ASAP7_75t_L g5345 ( 
.A(n_4607),
.B(n_17),
.Y(n_5345)
);

AO21x2_ASAP7_75t_L g5346 ( 
.A1(n_4668),
.A2(n_2550),
.B(n_2549),
.Y(n_5346)
);

A2O1A1Ixp33_ASAP7_75t_L g5347 ( 
.A1(n_4847),
.A2(n_1197),
.B(n_1201),
.C(n_1196),
.Y(n_5347)
);

INVxp67_ASAP7_75t_L g5348 ( 
.A(n_4735),
.Y(n_5348)
);

A2O1A1Ixp33_ASAP7_75t_L g5349 ( 
.A1(n_4847),
.A2(n_1205),
.B(n_1208),
.C(n_1204),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_4805),
.Y(n_5350)
);

INVx2_ASAP7_75t_L g5351 ( 
.A(n_4745),
.Y(n_5351)
);

AND2x2_ASAP7_75t_L g5352 ( 
.A(n_4607),
.B(n_17),
.Y(n_5352)
);

O2A1O1Ixp33_ASAP7_75t_SL g5353 ( 
.A1(n_4808),
.A2(n_67),
.B(n_69),
.C(n_66),
.Y(n_5353)
);

AOI22xp5_ASAP7_75t_L g5354 ( 
.A1(n_4976),
.A2(n_1214),
.B1(n_1217),
.B2(n_1211),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_4817),
.Y(n_5355)
);

AO31x2_ASAP7_75t_L g5356 ( 
.A1(n_4774),
.A2(n_2553),
.A3(n_2555),
.B(n_2552),
.Y(n_5356)
);

AOI22xp33_ASAP7_75t_L g5357 ( 
.A1(n_4887),
.A2(n_2552),
.B1(n_2555),
.B2(n_2553),
.Y(n_5357)
);

AOI22xp33_ASAP7_75t_L g5358 ( 
.A1(n_4871),
.A2(n_2560),
.B1(n_2567),
.B2(n_2564),
.Y(n_5358)
);

AO21x2_ASAP7_75t_L g5359 ( 
.A1(n_4668),
.A2(n_2564),
.B(n_2560),
.Y(n_5359)
);

INVx1_ASAP7_75t_L g5360 ( 
.A(n_4822),
.Y(n_5360)
);

O2A1O1Ixp33_ASAP7_75t_SL g5361 ( 
.A1(n_4825),
.A2(n_69),
.B(n_72),
.C(n_67),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4833),
.Y(n_5362)
);

O2A1O1Ixp33_ASAP7_75t_L g5363 ( 
.A1(n_4676),
.A2(n_2355),
.B(n_2358),
.C(n_2353),
.Y(n_5363)
);

NOR2xp33_ASAP7_75t_L g5364 ( 
.A(n_4886),
.B(n_72),
.Y(n_5364)
);

INVx2_ASAP7_75t_SL g5365 ( 
.A(n_4906),
.Y(n_5365)
);

A2O1A1Ixp33_ASAP7_75t_L g5366 ( 
.A1(n_4853),
.A2(n_1223),
.B(n_1225),
.C(n_1219),
.Y(n_5366)
);

AOI22xp33_ASAP7_75t_L g5367 ( 
.A1(n_4871),
.A2(n_2567),
.B1(n_2631),
.B2(n_2629),
.Y(n_5367)
);

AOI22xp5_ASAP7_75t_L g5368 ( 
.A1(n_4841),
.A2(n_1227),
.B1(n_1228),
.B2(n_1226),
.Y(n_5368)
);

BUFx8_ASAP7_75t_SL g5369 ( 
.A(n_4870),
.Y(n_5369)
);

INVx2_ASAP7_75t_L g5370 ( 
.A(n_4784),
.Y(n_5370)
);

OR2x2_ASAP7_75t_L g5371 ( 
.A(n_4676),
.B(n_19),
.Y(n_5371)
);

O2A1O1Ixp33_ASAP7_75t_L g5372 ( 
.A1(n_4686),
.A2(n_4949),
.B(n_4855),
.C(n_4839),
.Y(n_5372)
);

BUFx3_ASAP7_75t_L g5373 ( 
.A(n_4773),
.Y(n_5373)
);

CKINVDCx6p67_ASAP7_75t_R g5374 ( 
.A(n_4795),
.Y(n_5374)
);

BUFx3_ASAP7_75t_L g5375 ( 
.A(n_4859),
.Y(n_5375)
);

OA21x2_ASAP7_75t_L g5376 ( 
.A1(n_4686),
.A2(n_1231),
.B(n_1230),
.Y(n_5376)
);

AOI22xp33_ASAP7_75t_L g5377 ( 
.A1(n_4788),
.A2(n_2631),
.B1(n_2636),
.B2(n_2634),
.Y(n_5377)
);

O2A1O1Ixp33_ASAP7_75t_SL g5378 ( 
.A1(n_4851),
.A2(n_4855),
.B(n_4720),
.C(n_4718),
.Y(n_5378)
);

OAI21xp5_ASAP7_75t_L g5379 ( 
.A1(n_4852),
.A2(n_1234),
.B(n_1232),
.Y(n_5379)
);

NAND3xp33_ASAP7_75t_L g5380 ( 
.A(n_4907),
.B(n_1236),
.C(n_1235),
.Y(n_5380)
);

AOI211x1_ASAP7_75t_L g5381 ( 
.A1(n_4830),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_4793),
.Y(n_5382)
);

O2A1O1Ixp33_ASAP7_75t_L g5383 ( 
.A1(n_4711),
.A2(n_4744),
.B(n_4789),
.C(n_4743),
.Y(n_5383)
);

OAI221xp5_ASAP7_75t_L g5384 ( 
.A1(n_4907),
.A2(n_2378),
.B1(n_2395),
.B2(n_2376),
.C(n_2362),
.Y(n_5384)
);

OAI22xp33_ASAP7_75t_L g5385 ( 
.A1(n_4575),
.A2(n_3334),
.B1(n_3365),
.B2(n_3353),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_4845),
.Y(n_5386)
);

OAI21x1_ASAP7_75t_L g5387 ( 
.A1(n_4720),
.A2(n_2636),
.B(n_2634),
.Y(n_5387)
);

INVx2_ASAP7_75t_L g5388 ( 
.A(n_4796),
.Y(n_5388)
);

CKINVDCx11_ASAP7_75t_R g5389 ( 
.A(n_4870),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_SL g5390 ( 
.A(n_4747),
.B(n_3353),
.Y(n_5390)
);

AO31x2_ASAP7_75t_L g5391 ( 
.A1(n_4797),
.A2(n_4816),
.A3(n_4820),
.B(n_4801),
.Y(n_5391)
);

NAND2x1p5_ASAP7_75t_L g5392 ( 
.A(n_4736),
.B(n_3367),
.Y(n_5392)
);

OAI221xp5_ASAP7_75t_L g5393 ( 
.A1(n_4907),
.A2(n_2378),
.B1(n_2395),
.B2(n_2376),
.C(n_2362),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_4838),
.Y(n_5394)
);

O2A1O1Ixp33_ASAP7_75t_L g5395 ( 
.A1(n_4743),
.A2(n_4789),
.B(n_4798),
.C(n_4744),
.Y(n_5395)
);

INVx2_ASAP7_75t_L g5396 ( 
.A(n_5318),
.Y(n_5396)
);

OAI22xp5_ASAP7_75t_L g5397 ( 
.A1(n_5007),
.A2(n_4798),
.B1(n_4848),
.B2(n_4812),
.Y(n_5397)
);

AOI22xp33_ASAP7_75t_SL g5398 ( 
.A1(n_5376),
.A2(n_4747),
.B1(n_4691),
.B2(n_4733),
.Y(n_5398)
);

OR2x6_ASAP7_75t_L g5399 ( 
.A(n_5020),
.B(n_4632),
.Y(n_5399)
);

AND2x2_ASAP7_75t_L g5400 ( 
.A(n_5111),
.B(n_4812),
.Y(n_5400)
);

INVx2_ASAP7_75t_L g5401 ( 
.A(n_5318),
.Y(n_5401)
);

INVx2_ASAP7_75t_L g5402 ( 
.A(n_5318),
.Y(n_5402)
);

CKINVDCx5p33_ASAP7_75t_R g5403 ( 
.A(n_5025),
.Y(n_5403)
);

BUFx3_ASAP7_75t_L g5404 ( 
.A(n_4994),
.Y(n_5404)
);

AO31x2_ASAP7_75t_L g5405 ( 
.A1(n_5137),
.A2(n_4904),
.A3(n_4915),
.B(n_4901),
.Y(n_5405)
);

BUFx3_ASAP7_75t_L g5406 ( 
.A(n_5014),
.Y(n_5406)
);

AND2x2_ASAP7_75t_L g5407 ( 
.A(n_5145),
.B(n_4848),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5004),
.Y(n_5408)
);

NOR2x1_ASAP7_75t_SL g5409 ( 
.A(n_5297),
.B(n_5183),
.Y(n_5409)
);

INVxp33_ASAP7_75t_L g5410 ( 
.A(n_5028),
.Y(n_5410)
);

INVx2_ASAP7_75t_L g5411 ( 
.A(n_5391),
.Y(n_5411)
);

INVx2_ASAP7_75t_L g5412 ( 
.A(n_5391),
.Y(n_5412)
);

OAI22xp33_ASAP7_75t_L g5413 ( 
.A1(n_5092),
.A2(n_4733),
.B1(n_4717),
.B2(n_4714),
.Y(n_5413)
);

BUFx2_ASAP7_75t_L g5414 ( 
.A(n_5276),
.Y(n_5414)
);

NOR2xp33_ASAP7_75t_L g5415 ( 
.A(n_5031),
.B(n_4674),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_4996),
.Y(n_5416)
);

NAND2xp5_ASAP7_75t_L g5417 ( 
.A(n_5096),
.B(n_4846),
.Y(n_5417)
);

HB1xp67_ASAP7_75t_L g5418 ( 
.A(n_5218),
.Y(n_5418)
);

INVx2_ASAP7_75t_L g5419 ( 
.A(n_5391),
.Y(n_5419)
);

INVx1_ASAP7_75t_L g5420 ( 
.A(n_5001),
.Y(n_5420)
);

INVx3_ASAP7_75t_L g5421 ( 
.A(n_5086),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_5002),
.Y(n_5422)
);

OAI221xp5_ASAP7_75t_L g5423 ( 
.A1(n_5320),
.A2(n_4856),
.B1(n_4865),
.B2(n_4854),
.C(n_4849),
.Y(n_5423)
);

AOI22xp33_ASAP7_75t_L g5424 ( 
.A1(n_4990),
.A2(n_4691),
.B1(n_4888),
.B2(n_4869),
.Y(n_5424)
);

INVx2_ASAP7_75t_L g5425 ( 
.A(n_5029),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_5233),
.Y(n_5426)
);

OAI22xp5_ASAP7_75t_L g5427 ( 
.A1(n_5032),
.A2(n_4714),
.B1(n_4986),
.B2(n_4836),
.Y(n_5427)
);

INVxp67_ASAP7_75t_L g5428 ( 
.A(n_5052),
.Y(n_5428)
);

BUFx8_ASAP7_75t_SL g5429 ( 
.A(n_5149),
.Y(n_5429)
);

INVx2_ASAP7_75t_L g5430 ( 
.A(n_5036),
.Y(n_5430)
);

INVx2_ASAP7_75t_L g5431 ( 
.A(n_5073),
.Y(n_5431)
);

INVx2_ASAP7_75t_SL g5432 ( 
.A(n_5180),
.Y(n_5432)
);

INVx3_ASAP7_75t_L g5433 ( 
.A(n_5278),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_5241),
.Y(n_5434)
);

INVx4_ASAP7_75t_L g5435 ( 
.A(n_5005),
.Y(n_5435)
);

AOI22xp33_ASAP7_75t_L g5436 ( 
.A1(n_5227),
.A2(n_4691),
.B1(n_4894),
.B2(n_4890),
.Y(n_5436)
);

HB1xp67_ASAP7_75t_L g5437 ( 
.A(n_5103),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_5022),
.B(n_4899),
.Y(n_5438)
);

BUFx2_ASAP7_75t_L g5439 ( 
.A(n_5283),
.Y(n_5439)
);

INVx2_ASAP7_75t_L g5440 ( 
.A(n_5085),
.Y(n_5440)
);

BUFx2_ASAP7_75t_L g5441 ( 
.A(n_5060),
.Y(n_5441)
);

BUFx4f_ASAP7_75t_L g5442 ( 
.A(n_5181),
.Y(n_5442)
);

OAI22xp33_ASAP7_75t_L g5443 ( 
.A1(n_5168),
.A2(n_4717),
.B1(n_4714),
.B2(n_4818),
.Y(n_5443)
);

OAI21x1_ASAP7_75t_L g5444 ( 
.A1(n_4999),
.A2(n_4632),
.B(n_4903),
.Y(n_5444)
);

INVx4_ASAP7_75t_L g5445 ( 
.A(n_5017),
.Y(n_5445)
);

AOI21xp33_ASAP7_75t_L g5446 ( 
.A1(n_5200),
.A2(n_4818),
.B(n_4969),
.Y(n_5446)
);

AND2x2_ASAP7_75t_L g5447 ( 
.A(n_5163),
.B(n_4747),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5055),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5068),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5069),
.Y(n_5450)
);

O2A1O1Ixp5_ASAP7_75t_L g5451 ( 
.A1(n_4995),
.A2(n_4592),
.B(n_4574),
.C(n_4892),
.Y(n_5451)
);

INVx1_ASAP7_75t_SL g5452 ( 
.A(n_5030),
.Y(n_5452)
);

CKINVDCx8_ASAP7_75t_R g5453 ( 
.A(n_5115),
.Y(n_5453)
);

INVx2_ASAP7_75t_L g5454 ( 
.A(n_5099),
.Y(n_5454)
);

NAND2xp5_ASAP7_75t_L g5455 ( 
.A(n_5238),
.B(n_4751),
.Y(n_5455)
);

OAI222xp33_ASAP7_75t_L g5456 ( 
.A1(n_5190),
.A2(n_4863),
.B1(n_4818),
.B2(n_4717),
.C1(n_4643),
.C2(n_4592),
.Y(n_5456)
);

AND2x2_ASAP7_75t_L g5457 ( 
.A(n_5065),
.B(n_4747),
.Y(n_5457)
);

AOI22xp33_ASAP7_75t_L g5458 ( 
.A1(n_5376),
.A2(n_4691),
.B1(n_4717),
.B2(n_4924),
.Y(n_5458)
);

OR2x2_ASAP7_75t_L g5459 ( 
.A(n_5072),
.B(n_4970),
.Y(n_5459)
);

INVx1_ASAP7_75t_L g5460 ( 
.A(n_5084),
.Y(n_5460)
);

AOI22xp33_ASAP7_75t_SL g5461 ( 
.A1(n_5205),
.A2(n_4783),
.B1(n_4574),
.B2(n_4967),
.Y(n_5461)
);

INVx2_ASAP7_75t_L g5462 ( 
.A(n_5176),
.Y(n_5462)
);

NAND2xp5_ASAP7_75t_L g5463 ( 
.A(n_4997),
.B(n_4751),
.Y(n_5463)
);

INVx2_ASAP7_75t_L g5464 ( 
.A(n_5191),
.Y(n_5464)
);

AOI22xp33_ASAP7_75t_L g5465 ( 
.A1(n_5034),
.A2(n_4924),
.B1(n_4896),
.B2(n_4905),
.Y(n_5465)
);

OAI22xp33_ASAP7_75t_L g5466 ( 
.A1(n_5171),
.A2(n_4940),
.B1(n_4968),
.B2(n_4967),
.Y(n_5466)
);

AOI22xp33_ASAP7_75t_L g5467 ( 
.A1(n_5164),
.A2(n_4896),
.B1(n_4950),
.B2(n_4623),
.Y(n_5467)
);

OR2x6_ASAP7_75t_L g5468 ( 
.A(n_5297),
.B(n_5075),
.Y(n_5468)
);

OR2x6_ASAP7_75t_L g5469 ( 
.A(n_5297),
.B(n_5075),
.Y(n_5469)
);

AOI21xp33_ASAP7_75t_L g5470 ( 
.A1(n_5130),
.A2(n_4968),
.B(n_4967),
.Y(n_5470)
);

INVx2_ASAP7_75t_L g5471 ( 
.A(n_5207),
.Y(n_5471)
);

AOI22xp33_ASAP7_75t_L g5472 ( 
.A1(n_5197),
.A2(n_4623),
.B1(n_4625),
.B2(n_4598),
.Y(n_5472)
);

AOI22xp33_ASAP7_75t_L g5473 ( 
.A1(n_5015),
.A2(n_4623),
.B1(n_4625),
.B2(n_4598),
.Y(n_5473)
);

AOI22xp33_ASAP7_75t_L g5474 ( 
.A1(n_5155),
.A2(n_4625),
.B1(n_4598),
.B2(n_4922),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_5100),
.Y(n_5475)
);

AOI22xp33_ASAP7_75t_L g5476 ( 
.A1(n_5155),
.A2(n_4922),
.B1(n_4968),
.B2(n_4870),
.Y(n_5476)
);

OAI22xp5_ASAP7_75t_L g5477 ( 
.A1(n_5381),
.A2(n_4760),
.B1(n_4836),
.B2(n_4900),
.Y(n_5477)
);

AOI221xp5_ASAP7_75t_L g5478 ( 
.A1(n_5381),
.A2(n_4891),
.B1(n_4876),
.B2(n_23),
.C(n_21),
.Y(n_5478)
);

INVx3_ASAP7_75t_SL g5479 ( 
.A(n_5175),
.Y(n_5479)
);

AOI22xp33_ASAP7_75t_SL g5480 ( 
.A1(n_5219),
.A2(n_4783),
.B1(n_4940),
.B2(n_4836),
.Y(n_5480)
);

AOI22xp33_ASAP7_75t_L g5481 ( 
.A1(n_5208),
.A2(n_4815),
.B1(n_4790),
.B2(n_4903),
.Y(n_5481)
);

OR2x6_ASAP7_75t_L g5482 ( 
.A(n_5075),
.B(n_4783),
.Y(n_5482)
);

AND2x4_ASAP7_75t_L g5483 ( 
.A(n_5235),
.B(n_4634),
.Y(n_5483)
);

AOI22xp33_ASAP7_75t_L g5484 ( 
.A1(n_5208),
.A2(n_4815),
.B1(n_4790),
.B2(n_2642),
.Y(n_5484)
);

INVx2_ASAP7_75t_SL g5485 ( 
.A(n_5373),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5108),
.Y(n_5486)
);

INVxp67_ASAP7_75t_L g5487 ( 
.A(n_5053),
.Y(n_5487)
);

AOI22xp33_ASAP7_75t_L g5488 ( 
.A1(n_5252),
.A2(n_2642),
.B1(n_2656),
.B2(n_2652),
.Y(n_5488)
);

NAND2x1p5_ASAP7_75t_L g5489 ( 
.A(n_5064),
.B(n_4741),
.Y(n_5489)
);

INVx1_ASAP7_75t_SL g5490 ( 
.A(n_5127),
.Y(n_5490)
);

AOI22xp33_ASAP7_75t_L g5491 ( 
.A1(n_5267),
.A2(n_5272),
.B1(n_5189),
.B2(n_5152),
.Y(n_5491)
);

AOI221xp5_ASAP7_75t_L g5492 ( 
.A1(n_5253),
.A2(n_4891),
.B1(n_4876),
.B2(n_23),
.C(n_21),
.Y(n_5492)
);

AOI22xp33_ASAP7_75t_L g5493 ( 
.A1(n_5024),
.A2(n_2652),
.B1(n_2659),
.B2(n_2656),
.Y(n_5493)
);

NAND2xp5_ASAP7_75t_L g5494 ( 
.A(n_5383),
.B(n_4751),
.Y(n_5494)
);

AND2x2_ASAP7_75t_L g5495 ( 
.A(n_5209),
.B(n_4659),
.Y(n_5495)
);

CKINVDCx20_ASAP7_75t_R g5496 ( 
.A(n_5167),
.Y(n_5496)
);

INVxp67_ASAP7_75t_L g5497 ( 
.A(n_5133),
.Y(n_5497)
);

AND2x2_ASAP7_75t_L g5498 ( 
.A(n_5080),
.B(n_4659),
.Y(n_5498)
);

CKINVDCx5p33_ASAP7_75t_R g5499 ( 
.A(n_5162),
.Y(n_5499)
);

AND2x4_ASAP7_75t_L g5500 ( 
.A(n_5235),
.B(n_4634),
.Y(n_5500)
);

OR2x2_ASAP7_75t_L g5501 ( 
.A(n_5348),
.B(n_4769),
.Y(n_5501)
);

OAI211xp5_ASAP7_75t_L g5502 ( 
.A1(n_5107),
.A2(n_4892),
.B(n_4875),
.C(n_4693),
.Y(n_5502)
);

CKINVDCx11_ASAP7_75t_R g5503 ( 
.A(n_4998),
.Y(n_5503)
);

AND2x4_ASAP7_75t_L g5504 ( 
.A(n_5024),
.B(n_5278),
.Y(n_5504)
);

INVx1_ASAP7_75t_SL g5505 ( 
.A(n_5057),
.Y(n_5505)
);

AND2x4_ASAP7_75t_L g5506 ( 
.A(n_5281),
.B(n_4700),
.Y(n_5506)
);

AND2x2_ASAP7_75t_L g5507 ( 
.A(n_5184),
.B(n_4693),
.Y(n_5507)
);

AO21x2_ASAP7_75t_L g5508 ( 
.A1(n_5109),
.A2(n_4984),
.B(n_4700),
.Y(n_5508)
);

OR2x2_ASAP7_75t_L g5509 ( 
.A(n_5042),
.B(n_5049),
.Y(n_5509)
);

INVx1_ASAP7_75t_SL g5510 ( 
.A(n_5141),
.Y(n_5510)
);

OAI21xp5_ASAP7_75t_L g5511 ( 
.A1(n_5008),
.A2(n_4852),
.B(n_4931),
.Y(n_5511)
);

INVx2_ASAP7_75t_L g5512 ( 
.A(n_5212),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5110),
.Y(n_5513)
);

AOI322xp5_ASAP7_75t_L g5514 ( 
.A1(n_5188),
.A2(n_27),
.A3(n_26),
.B1(n_24),
.B2(n_28),
.C1(n_23),
.C2(n_25),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5116),
.Y(n_5515)
);

A2O1A1Ixp33_ASAP7_75t_L g5516 ( 
.A1(n_4991),
.A2(n_4779),
.B(n_4804),
.C(n_4769),
.Y(n_5516)
);

OAI21xp5_ASAP7_75t_L g5517 ( 
.A1(n_4992),
.A2(n_4954),
.B(n_4931),
.Y(n_5517)
);

AOI22xp33_ASAP7_75t_L g5518 ( 
.A1(n_5220),
.A2(n_2659),
.B1(n_2673),
.B2(n_2660),
.Y(n_5518)
);

AOI22xp33_ASAP7_75t_L g5519 ( 
.A1(n_5011),
.A2(n_2660),
.B1(n_2675),
.B2(n_2673),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5118),
.Y(n_5520)
);

AOI22xp33_ASAP7_75t_L g5521 ( 
.A1(n_5291),
.A2(n_2675),
.B1(n_2684),
.B2(n_2682),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_5213),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5121),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_5214),
.Y(n_5524)
);

CKINVDCx20_ASAP7_75t_R g5525 ( 
.A(n_5285),
.Y(n_5525)
);

INVx2_ASAP7_75t_L g5526 ( 
.A(n_5257),
.Y(n_5526)
);

NAND2x1p5_ASAP7_75t_L g5527 ( 
.A(n_5390),
.B(n_4741),
.Y(n_5527)
);

CKINVDCx6p67_ASAP7_75t_R g5528 ( 
.A(n_5124),
.Y(n_5528)
);

A2O1A1Ixp33_ASAP7_75t_L g5529 ( 
.A1(n_5006),
.A2(n_4804),
.B(n_4779),
.C(n_4866),
.Y(n_5529)
);

INVx1_ASAP7_75t_L g5530 ( 
.A(n_5128),
.Y(n_5530)
);

AOI21xp5_ASAP7_75t_L g5531 ( 
.A1(n_5063),
.A2(n_4984),
.B(n_4954),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_5138),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_5142),
.Y(n_5533)
);

AND2x2_ASAP7_75t_L g5534 ( 
.A(n_5317),
.B(n_4703),
.Y(n_5534)
);

INVx2_ASAP7_75t_L g5535 ( 
.A(n_5269),
.Y(n_5535)
);

OAI22xp5_ASAP7_75t_L g5536 ( 
.A1(n_5193),
.A2(n_4760),
.B1(n_4900),
.B2(n_4875),
.Y(n_5536)
);

CKINVDCx5p33_ASAP7_75t_R g5537 ( 
.A(n_5105),
.Y(n_5537)
);

AOI22xp33_ASAP7_75t_L g5538 ( 
.A1(n_5291),
.A2(n_2682),
.B1(n_2691),
.B2(n_2684),
.Y(n_5538)
);

AOI21xp5_ASAP7_75t_L g5539 ( 
.A1(n_5016),
.A2(n_4900),
.B(n_4756),
.Y(n_5539)
);

OAI21xp5_ASAP7_75t_L g5540 ( 
.A1(n_5171),
.A2(n_4900),
.B(n_4756),
.Y(n_5540)
);

BUFx6f_ASAP7_75t_L g5541 ( 
.A(n_5310),
.Y(n_5541)
);

INVx2_ASAP7_75t_L g5542 ( 
.A(n_5293),
.Y(n_5542)
);

AND2x2_ASAP7_75t_L g5543 ( 
.A(n_5146),
.B(n_4703),
.Y(n_5543)
);

AOI221xp5_ASAP7_75t_L g5544 ( 
.A1(n_5287),
.A2(n_4891),
.B1(n_4876),
.B2(n_29),
.C(n_22),
.Y(n_5544)
);

CKINVDCx11_ASAP7_75t_R g5545 ( 
.A(n_4998),
.Y(n_5545)
);

A2O1A1Ixp33_ASAP7_75t_L g5546 ( 
.A1(n_5107),
.A2(n_4734),
.B(n_4802),
.C(n_4682),
.Y(n_5546)
);

NOR2x1_ASAP7_75t_L g5547 ( 
.A(n_5375),
.B(n_5173),
.Y(n_5547)
);

AOI221xp5_ASAP7_75t_L g5548 ( 
.A1(n_5308),
.A2(n_29),
.B1(n_22),
.B2(n_24),
.C(n_30),
.Y(n_5548)
);

OAI22xp5_ASAP7_75t_L g5549 ( 
.A1(n_5193),
.A2(n_4832),
.B1(n_4756),
.B2(n_4741),
.Y(n_5549)
);

OR2x2_ASAP7_75t_L g5550 ( 
.A(n_5386),
.B(n_4734),
.Y(n_5550)
);

AOI22xp33_ASAP7_75t_L g5551 ( 
.A1(n_5303),
.A2(n_2691),
.B1(n_2699),
.B2(n_2694),
.Y(n_5551)
);

INVx2_ASAP7_75t_L g5552 ( 
.A(n_5333),
.Y(n_5552)
);

BUFx6f_ASAP7_75t_L g5553 ( 
.A(n_5088),
.Y(n_5553)
);

O2A1O1Ixp5_ASAP7_75t_L g5554 ( 
.A1(n_5221),
.A2(n_4832),
.B(n_31),
.C(n_22),
.Y(n_5554)
);

AND2x2_ASAP7_75t_L g5555 ( 
.A(n_5245),
.B(n_4734),
.Y(n_5555)
);

INVx2_ASAP7_75t_L g5556 ( 
.A(n_5351),
.Y(n_5556)
);

INVx3_ASAP7_75t_L g5557 ( 
.A(n_5281),
.Y(n_5557)
);

CKINVDCx5p33_ASAP7_75t_R g5558 ( 
.A(n_5140),
.Y(n_5558)
);

INVx2_ASAP7_75t_SL g5559 ( 
.A(n_5258),
.Y(n_5559)
);

OAI21x1_ASAP7_75t_L g5560 ( 
.A1(n_5009),
.A2(n_4643),
.B(n_4741),
.Y(n_5560)
);

OAI22xp5_ASAP7_75t_L g5561 ( 
.A1(n_5303),
.A2(n_4756),
.B1(n_4806),
.B2(n_4802),
.Y(n_5561)
);

AOI22xp33_ASAP7_75t_L g5562 ( 
.A1(n_5094),
.A2(n_2694),
.B1(n_2703),
.B2(n_2699),
.Y(n_5562)
);

OAI211xp5_ASAP7_75t_SL g5563 ( 
.A1(n_5125),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_5563)
);

AOI21xp5_ASAP7_75t_L g5564 ( 
.A1(n_5098),
.A2(n_4937),
.B(n_4917),
.Y(n_5564)
);

BUFx12f_ASAP7_75t_L g5565 ( 
.A(n_5115),
.Y(n_5565)
);

OR2x2_ASAP7_75t_L g5566 ( 
.A(n_5192),
.B(n_4802),
.Y(n_5566)
);

OAI22xp5_ASAP7_75t_SL g5567 ( 
.A1(n_5339),
.A2(n_4813),
.B1(n_4828),
.B2(n_4806),
.Y(n_5567)
);

BUFx6f_ASAP7_75t_L g5568 ( 
.A(n_5088),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_5216),
.Y(n_5569)
);

AOI221xp5_ASAP7_75t_L g5570 ( 
.A1(n_5337),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.C(n_33),
.Y(n_5570)
);

OAI22xp5_ASAP7_75t_L g5571 ( 
.A1(n_5003),
.A2(n_4813),
.B1(n_4828),
.B2(n_4806),
.Y(n_5571)
);

AOI22xp33_ASAP7_75t_L g5572 ( 
.A1(n_5217),
.A2(n_2703),
.B1(n_2716),
.B2(n_2713),
.Y(n_5572)
);

OR2x2_ASAP7_75t_L g5573 ( 
.A(n_5242),
.B(n_4813),
.Y(n_5573)
);

INVx2_ASAP7_75t_L g5574 ( 
.A(n_5370),
.Y(n_5574)
);

AOI21xp5_ASAP7_75t_L g5575 ( 
.A1(n_5027),
.A2(n_4937),
.B(n_4917),
.Y(n_5575)
);

OAI21xp33_ASAP7_75t_SL g5576 ( 
.A1(n_5326),
.A2(n_4828),
.B(n_32),
.Y(n_5576)
);

OAI21x1_ASAP7_75t_L g5577 ( 
.A1(n_5256),
.A2(n_2716),
.B(n_2713),
.Y(n_5577)
);

INVx1_ASAP7_75t_L g5578 ( 
.A(n_5262),
.Y(n_5578)
);

AND2x4_ASAP7_75t_L g5579 ( 
.A(n_5132),
.B(n_4917),
.Y(n_5579)
);

AO31x2_ASAP7_75t_L g5580 ( 
.A1(n_5234),
.A2(n_2417),
.A3(n_2418),
.B(n_2413),
.Y(n_5580)
);

AND2x2_ASAP7_75t_L g5581 ( 
.A(n_5365),
.B(n_4937),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_5288),
.Y(n_5582)
);

AOI22xp5_ASAP7_75t_L g5583 ( 
.A1(n_5131),
.A2(n_1880),
.B1(n_2961),
.B2(n_2957),
.Y(n_5583)
);

OAI22xp5_ASAP7_75t_L g5584 ( 
.A1(n_5322),
.A2(n_3367),
.B1(n_3370),
.B2(n_3365),
.Y(n_5584)
);

O2A1O1Ixp5_ASAP7_75t_L g5585 ( 
.A1(n_5228),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_L g5586 ( 
.A(n_5395),
.B(n_5372),
.Y(n_5586)
);

AND2x2_ASAP7_75t_L g5587 ( 
.A(n_5056),
.B(n_33),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5289),
.Y(n_5588)
);

OAI21x1_ASAP7_75t_L g5589 ( 
.A1(n_5178),
.A2(n_2725),
.B(n_2721),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5295),
.Y(n_5590)
);

NOR2x1_ASAP7_75t_SL g5591 ( 
.A(n_5088),
.B(n_3365),
.Y(n_5591)
);

NAND2xp33_ASAP7_75t_L g5592 ( 
.A(n_5240),
.B(n_3365),
.Y(n_5592)
);

AOI22xp33_ASAP7_75t_L g5593 ( 
.A1(n_5199),
.A2(n_2721),
.B1(n_2733),
.B2(n_2725),
.Y(n_5593)
);

OAI22xp5_ASAP7_75t_L g5594 ( 
.A1(n_5371),
.A2(n_3370),
.B1(n_3375),
.B2(n_3367),
.Y(n_5594)
);

BUFx3_ASAP7_75t_L g5595 ( 
.A(n_5018),
.Y(n_5595)
);

OAI221xp5_ASAP7_75t_L g5596 ( 
.A1(n_5125),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.C(n_38),
.Y(n_5596)
);

NAND2x1p5_ASAP7_75t_L g5597 ( 
.A(n_5135),
.B(n_3370),
.Y(n_5597)
);

INVx6_ASAP7_75t_L g5598 ( 
.A(n_5097),
.Y(n_5598)
);

OR2x2_ASAP7_75t_L g5599 ( 
.A(n_5298),
.B(n_36),
.Y(n_5599)
);

NAND2xp5_ASAP7_75t_L g5600 ( 
.A(n_5315),
.B(n_36),
.Y(n_5600)
);

OAI22xp33_ASAP7_75t_L g5601 ( 
.A1(n_5165),
.A2(n_3375),
.B1(n_3388),
.B2(n_3381),
.Y(n_5601)
);

AOI22xp33_ASAP7_75t_L g5602 ( 
.A1(n_5210),
.A2(n_2733),
.B1(n_2738),
.B2(n_2737),
.Y(n_5602)
);

OA22x2_ASAP7_75t_L g5603 ( 
.A1(n_5147),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_5603)
);

AOI22xp33_ASAP7_75t_L g5604 ( 
.A1(n_5039),
.A2(n_2737),
.B1(n_2743),
.B2(n_2738),
.Y(n_5604)
);

AOI22xp33_ASAP7_75t_L g5605 ( 
.A1(n_5312),
.A2(n_2743),
.B1(n_2776),
.B2(n_2769),
.Y(n_5605)
);

AND2x2_ASAP7_75t_L g5606 ( 
.A(n_5000),
.B(n_37),
.Y(n_5606)
);

CKINVDCx6p67_ASAP7_75t_R g5607 ( 
.A(n_5274),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_5301),
.Y(n_5608)
);

NAND2xp5_ASAP7_75t_L g5609 ( 
.A(n_5350),
.B(n_5355),
.Y(n_5609)
);

AND2x4_ASAP7_75t_L g5610 ( 
.A(n_5360),
.B(n_2998),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5362),
.Y(n_5611)
);

OAI22xp5_ASAP7_75t_L g5612 ( 
.A1(n_5259),
.A2(n_3388),
.B1(n_3381),
.B2(n_74),
.Y(n_5612)
);

BUFx2_ASAP7_75t_L g5613 ( 
.A(n_5369),
.Y(n_5613)
);

OAI22xp5_ASAP7_75t_L g5614 ( 
.A1(n_5259),
.A2(n_3388),
.B1(n_3381),
.B2(n_75),
.Y(n_5614)
);

INVx2_ASAP7_75t_L g5615 ( 
.A(n_5382),
.Y(n_5615)
);

OAI22xp5_ASAP7_75t_L g5616 ( 
.A1(n_5143),
.A2(n_3388),
.B1(n_3381),
.B2(n_76),
.Y(n_5616)
);

INVxp67_ASAP7_75t_L g5617 ( 
.A(n_5074),
.Y(n_5617)
);

OAI22xp5_ASAP7_75t_L g5618 ( 
.A1(n_5231),
.A2(n_77),
.B1(n_78),
.B2(n_73),
.Y(n_5618)
);

OAI22xp5_ASAP7_75t_L g5619 ( 
.A1(n_5271),
.A2(n_79),
.B1(n_80),
.B2(n_77),
.Y(n_5619)
);

O2A1O1Ixp33_ASAP7_75t_SL g5620 ( 
.A1(n_5071),
.A2(n_5306),
.B(n_5251),
.C(n_5254),
.Y(n_5620)
);

NAND2x1_ASAP7_75t_L g5621 ( 
.A(n_5122),
.B(n_5093),
.Y(n_5621)
);

INVxp67_ASAP7_75t_L g5622 ( 
.A(n_5058),
.Y(n_5622)
);

AOI22xp33_ASAP7_75t_L g5623 ( 
.A1(n_5266),
.A2(n_2789),
.B1(n_2802),
.B2(n_2783),
.Y(n_5623)
);

AND2x2_ASAP7_75t_L g5624 ( 
.A(n_5374),
.B(n_38),
.Y(n_5624)
);

AOI22xp33_ASAP7_75t_L g5625 ( 
.A1(n_5013),
.A2(n_5286),
.B1(n_5394),
.B2(n_5388),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5083),
.Y(n_5626)
);

INVx1_ASAP7_75t_SL g5627 ( 
.A(n_5389),
.Y(n_5627)
);

OAI22xp5_ASAP7_75t_L g5628 ( 
.A1(n_5129),
.A2(n_81),
.B1(n_83),
.B2(n_79),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5114),
.Y(n_5629)
);

INVx2_ASAP7_75t_L g5630 ( 
.A(n_5134),
.Y(n_5630)
);

AOI22xp5_ASAP7_75t_L g5631 ( 
.A1(n_5054),
.A2(n_1880),
.B1(n_3173),
.B2(n_2961),
.Y(n_5631)
);

BUFx2_ASAP7_75t_L g5632 ( 
.A(n_5093),
.Y(n_5632)
);

INVx1_ASAP7_75t_L g5633 ( 
.A(n_5091),
.Y(n_5633)
);

INVx1_ASAP7_75t_SL g5634 ( 
.A(n_5330),
.Y(n_5634)
);

BUFx2_ASAP7_75t_L g5635 ( 
.A(n_5302),
.Y(n_5635)
);

BUFx12f_ASAP7_75t_L g5636 ( 
.A(n_5097),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_SL g5637 ( 
.A(n_5097),
.B(n_2998),
.Y(n_5637)
);

AOI22xp33_ASAP7_75t_L g5638 ( 
.A1(n_5380),
.A2(n_2769),
.B1(n_2777),
.B2(n_2776),
.Y(n_5638)
);

AOI21xp33_ASAP7_75t_L g5639 ( 
.A1(n_5284),
.A2(n_41),
.B(n_40),
.Y(n_5639)
);

AOI22xp33_ASAP7_75t_L g5640 ( 
.A1(n_5136),
.A2(n_2777),
.B1(n_2783),
.B2(n_2778),
.Y(n_5640)
);

AND2x2_ASAP7_75t_L g5641 ( 
.A(n_5106),
.B(n_39),
.Y(n_5641)
);

BUFx12f_ASAP7_75t_L g5642 ( 
.A(n_5179),
.Y(n_5642)
);

OAI222xp33_ASAP7_75t_L g5643 ( 
.A1(n_5344),
.A2(n_2811),
.B1(n_2789),
.B2(n_2802),
.C1(n_2778),
.C2(n_42),
.Y(n_5643)
);

NOR2xp33_ASAP7_75t_L g5644 ( 
.A(n_5148),
.B(n_84),
.Y(n_5644)
);

AOI22xp5_ASAP7_75t_L g5645 ( 
.A1(n_5047),
.A2(n_1880),
.B1(n_3173),
.B2(n_2961),
.Y(n_5645)
);

OAI21xp33_ASAP7_75t_SL g5646 ( 
.A1(n_5292),
.A2(n_40),
.B(n_41),
.Y(n_5646)
);

NOR2xp33_ASAP7_75t_L g5647 ( 
.A(n_5043),
.B(n_85),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_5091),
.Y(n_5648)
);

INVx1_ASAP7_75t_L g5649 ( 
.A(n_5091),
.Y(n_5649)
);

INVx2_ASAP7_75t_L g5650 ( 
.A(n_5134),
.Y(n_5650)
);

AOI221xp5_ASAP7_75t_L g5651 ( 
.A1(n_5126),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.C(n_87),
.Y(n_5651)
);

AND2x2_ASAP7_75t_L g5652 ( 
.A(n_5345),
.B(n_5352),
.Y(n_5652)
);

NAND2xp5_ASAP7_75t_SL g5653 ( 
.A(n_5179),
.B(n_2998),
.Y(n_5653)
);

CKINVDCx6p67_ASAP7_75t_R g5654 ( 
.A(n_5204),
.Y(n_5654)
);

AOI221xp5_ASAP7_75t_L g5655 ( 
.A1(n_5023),
.A2(n_42),
.B1(n_43),
.B2(n_89),
.C(n_90),
.Y(n_5655)
);

INVx2_ASAP7_75t_SL g5656 ( 
.A(n_5179),
.Y(n_5656)
);

OAI22xp5_ASAP7_75t_L g5657 ( 
.A1(n_5299),
.A2(n_93),
.B1(n_89),
.B2(n_92),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_5307),
.Y(n_5658)
);

BUFx3_ASAP7_75t_L g5659 ( 
.A(n_5309),
.Y(n_5659)
);

INVx2_ASAP7_75t_L g5660 ( 
.A(n_5134),
.Y(n_5660)
);

AOI22xp33_ASAP7_75t_L g5661 ( 
.A1(n_5050),
.A2(n_2811),
.B1(n_3173),
.B2(n_2961),
.Y(n_5661)
);

AND2x2_ASAP7_75t_SL g5662 ( 
.A(n_5120),
.B(n_3360),
.Y(n_5662)
);

AOI322xp5_ASAP7_75t_L g5663 ( 
.A1(n_5035),
.A2(n_97),
.A3(n_96),
.B1(n_94),
.B2(n_92),
.C1(n_93),
.C2(n_95),
.Y(n_5663)
);

INVx4_ASAP7_75t_L g5664 ( 
.A(n_5309),
.Y(n_5664)
);

AOI21xp5_ASAP7_75t_L g5665 ( 
.A1(n_5021),
.A2(n_5117),
.B(n_5104),
.Y(n_5665)
);

AOI22xp33_ASAP7_75t_L g5666 ( 
.A1(n_5050),
.A2(n_3173),
.B1(n_3233),
.B2(n_3188),
.Y(n_5666)
);

AOI221xp5_ASAP7_75t_L g5667 ( 
.A1(n_5353),
.A2(n_99),
.B1(n_94),
.B2(n_96),
.C(n_100),
.Y(n_5667)
);

AOI22xp33_ASAP7_75t_L g5668 ( 
.A1(n_5095),
.A2(n_3188),
.B1(n_3294),
.B2(n_3233),
.Y(n_5668)
);

AND2x4_ASAP7_75t_L g5669 ( 
.A(n_5122),
.B(n_3062),
.Y(n_5669)
);

CKINVDCx5p33_ASAP7_75t_R g5670 ( 
.A(n_5204),
.Y(n_5670)
);

AO221x1_ASAP7_75t_L g5671 ( 
.A1(n_5161),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.C(n_102),
.Y(n_5671)
);

AOI22xp5_ASAP7_75t_SL g5672 ( 
.A1(n_5122),
.A2(n_3233),
.B1(n_3294),
.B2(n_3188),
.Y(n_5672)
);

AOI22xp33_ASAP7_75t_SL g5673 ( 
.A1(n_5344),
.A2(n_3188),
.B1(n_3294),
.B2(n_3233),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_5222),
.Y(n_5674)
);

AOI22xp33_ASAP7_75t_L g5675 ( 
.A1(n_5095),
.A2(n_3188),
.B1(n_3294),
.B2(n_3233),
.Y(n_5675)
);

AND2x2_ASAP7_75t_L g5676 ( 
.A(n_5302),
.B(n_101),
.Y(n_5676)
);

INVx2_ASAP7_75t_L g5677 ( 
.A(n_5346),
.Y(n_5677)
);

AOI22xp33_ASAP7_75t_L g5678 ( 
.A1(n_5268),
.A2(n_3188),
.B1(n_3294),
.B2(n_2403),
.Y(n_5678)
);

OAI21xp5_ASAP7_75t_SL g5679 ( 
.A1(n_5174),
.A2(n_103),
.B(n_104),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5222),
.Y(n_5680)
);

INVx1_ASAP7_75t_L g5681 ( 
.A(n_5222),
.Y(n_5681)
);

AOI22xp33_ASAP7_75t_L g5682 ( 
.A1(n_5357),
.A2(n_3294),
.B1(n_2403),
.B2(n_2341),
.Y(n_5682)
);

BUFx2_ASAP7_75t_L g5683 ( 
.A(n_5336),
.Y(n_5683)
);

OAI22xp5_ASAP7_75t_L g5684 ( 
.A1(n_5170),
.A2(n_107),
.B1(n_104),
.B2(n_106),
.Y(n_5684)
);

INVxp67_ASAP7_75t_L g5685 ( 
.A(n_5327),
.Y(n_5685)
);

AOI221xp5_ASAP7_75t_L g5686 ( 
.A1(n_5361),
.A2(n_5263),
.B1(n_5203),
.B2(n_5153),
.C(n_5250),
.Y(n_5686)
);

OAI221xp5_ASAP7_75t_L g5687 ( 
.A1(n_5139),
.A2(n_2406),
.B1(n_2407),
.B2(n_2404),
.C(n_2399),
.Y(n_5687)
);

OAI22xp5_ASAP7_75t_L g5688 ( 
.A1(n_5154),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_5688)
);

AOI22xp33_ASAP7_75t_SL g5689 ( 
.A1(n_5344),
.A2(n_3360),
.B1(n_3062),
.B2(n_113),
.Y(n_5689)
);

AOI22xp33_ASAP7_75t_SL g5690 ( 
.A1(n_5232),
.A2(n_3360),
.B1(n_3062),
.B2(n_113),
.Y(n_5690)
);

INVx2_ASAP7_75t_L g5691 ( 
.A(n_5346),
.Y(n_5691)
);

AOI22xp33_ASAP7_75t_L g5692 ( 
.A1(n_5354),
.A2(n_2403),
.B1(n_2341),
.B2(n_2348),
.Y(n_5692)
);

OR2x2_ASAP7_75t_L g5693 ( 
.A(n_5119),
.B(n_5311),
.Y(n_5693)
);

OAI21x1_ASAP7_75t_L g5694 ( 
.A1(n_5045),
.A2(n_2403),
.B(n_2413),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_L g5695 ( 
.A(n_5010),
.B(n_109),
.Y(n_5695)
);

OAI22xp5_ASAP7_75t_L g5696 ( 
.A1(n_5159),
.A2(n_114),
.B1(n_109),
.B2(n_110),
.Y(n_5696)
);

OR2x2_ASAP7_75t_L g5697 ( 
.A(n_5311),
.B(n_110),
.Y(n_5697)
);

AND2x4_ASAP7_75t_L g5698 ( 
.A(n_5122),
.B(n_114),
.Y(n_5698)
);

AOI22xp33_ASAP7_75t_L g5699 ( 
.A1(n_5354),
.A2(n_2348),
.B1(n_2369),
.B2(n_2336),
.Y(n_5699)
);

OAI22xp33_ASAP7_75t_L g5700 ( 
.A1(n_5160),
.A2(n_3138),
.B1(n_2404),
.B2(n_2406),
.Y(n_5700)
);

BUFx12f_ASAP7_75t_L g5701 ( 
.A(n_5182),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5314),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5311),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5261),
.Y(n_5704)
);

BUFx8_ASAP7_75t_L g5705 ( 
.A(n_5232),
.Y(n_5705)
);

NAND2xp5_ASAP7_75t_L g5706 ( 
.A(n_5010),
.B(n_116),
.Y(n_5706)
);

INVx1_ASAP7_75t_SL g5707 ( 
.A(n_5316),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5261),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_5010),
.B(n_116),
.Y(n_5709)
);

OAI22xp5_ASAP7_75t_L g5710 ( 
.A1(n_5206),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5261),
.Y(n_5711)
);

OAI22xp5_ASAP7_75t_L g5712 ( 
.A1(n_5255),
.A2(n_120),
.B1(n_117),
.B2(n_119),
.Y(n_5712)
);

O2A1O1Ixp33_ASAP7_75t_SL g5713 ( 
.A1(n_5347),
.A2(n_5366),
.B(n_5349),
.C(n_5364),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_5309),
.B(n_120),
.Y(n_5714)
);

AOI21xp33_ASAP7_75t_L g5715 ( 
.A1(n_5343),
.A2(n_5363),
.B(n_5264),
.Y(n_5715)
);

INVx2_ASAP7_75t_L g5716 ( 
.A(n_5359),
.Y(n_5716)
);

OAI211xp5_ASAP7_75t_L g5717 ( 
.A1(n_5280),
.A2(n_124),
.B(n_121),
.C(n_123),
.Y(n_5717)
);

INVx2_ASAP7_75t_L g5718 ( 
.A(n_5359),
.Y(n_5718)
);

AOI22xp33_ASAP7_75t_L g5719 ( 
.A1(n_5377),
.A2(n_2369),
.B1(n_2336),
.B2(n_2417),
.Y(n_5719)
);

BUFx12f_ASAP7_75t_L g5720 ( 
.A(n_5182),
.Y(n_5720)
);

OAI21x1_ASAP7_75t_L g5721 ( 
.A1(n_5342),
.A2(n_2420),
.B(n_2418),
.Y(n_5721)
);

INVx1_ASAP7_75t_SL g5722 ( 
.A(n_5321),
.Y(n_5722)
);

AND2x2_ASAP7_75t_L g5723 ( 
.A(n_5033),
.B(n_121),
.Y(n_5723)
);

AOI21xp5_ASAP7_75t_L g5724 ( 
.A1(n_5051),
.A2(n_3138),
.B(n_2407),
.Y(n_5724)
);

CKINVDCx20_ASAP7_75t_R g5725 ( 
.A(n_5305),
.Y(n_5725)
);

AOI22xp33_ASAP7_75t_L g5726 ( 
.A1(n_5067),
.A2(n_2420),
.B1(n_2441),
.B2(n_2426),
.Y(n_5726)
);

OAI22xp5_ASAP7_75t_L g5727 ( 
.A1(n_5296),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_5727)
);

INVx3_ASAP7_75t_L g5728 ( 
.A(n_5305),
.Y(n_5728)
);

OAI22xp5_ASAP7_75t_L g5729 ( 
.A1(n_5239),
.A2(n_128),
.B1(n_125),
.B2(n_126),
.Y(n_5729)
);

OAI21xp5_ASAP7_75t_L g5730 ( 
.A1(n_5332),
.A2(n_2399),
.B(n_2426),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5248),
.Y(n_5731)
);

O2A1O1Ixp33_ASAP7_75t_L g5732 ( 
.A1(n_5187),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_5732)
);

AND2x2_ASAP7_75t_L g5733 ( 
.A(n_5033),
.B(n_129),
.Y(n_5733)
);

OAI22xp5_ASAP7_75t_L g5734 ( 
.A1(n_5225),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_5734)
);

AOI22xp33_ASAP7_75t_L g5735 ( 
.A1(n_5067),
.A2(n_2446),
.B1(n_2453),
.B2(n_2441),
.Y(n_5735)
);

AOI21xp33_ASAP7_75t_L g5736 ( 
.A1(n_5329),
.A2(n_131),
.B(n_133),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_5248),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_5378),
.Y(n_5738)
);

AOI21xp5_ASAP7_75t_L g5739 ( 
.A1(n_5101),
.A2(n_3138),
.B(n_2428),
.Y(n_5739)
);

INVx2_ASAP7_75t_L g5740 ( 
.A(n_5328),
.Y(n_5740)
);

NAND2xp5_ASAP7_75t_L g5741 ( 
.A(n_5033),
.B(n_133),
.Y(n_5741)
);

NAND2xp5_ASAP7_75t_L g5742 ( 
.A(n_5041),
.B(n_134),
.Y(n_5742)
);

AOI22xp33_ASAP7_75t_L g5743 ( 
.A1(n_5368),
.A2(n_2453),
.B1(n_2456),
.B2(n_2446),
.Y(n_5743)
);

NOR2xp33_ASAP7_75t_L g5744 ( 
.A(n_5685),
.B(n_5040),
.Y(n_5744)
);

AOI21x1_ASAP7_75t_L g5745 ( 
.A1(n_5600),
.A2(n_5340),
.B(n_5211),
.Y(n_5745)
);

HB1xp67_ASAP7_75t_L g5746 ( 
.A(n_5418),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5426),
.Y(n_5747)
);

INVx2_ASAP7_75t_L g5748 ( 
.A(n_5411),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5434),
.Y(n_5749)
);

OR2x2_ASAP7_75t_L g5750 ( 
.A(n_5490),
.B(n_5195),
.Y(n_5750)
);

OAI21x1_ASAP7_75t_SL g5751 ( 
.A1(n_5435),
.A2(n_5185),
.B(n_5198),
.Y(n_5751)
);

INVx4_ASAP7_75t_L g5752 ( 
.A(n_5541),
.Y(n_5752)
);

INVx2_ASAP7_75t_SL g5753 ( 
.A(n_5541),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5412),
.Y(n_5754)
);

AOI221xp5_ASAP7_75t_L g5755 ( 
.A1(n_5639),
.A2(n_5177),
.B1(n_5082),
.B2(n_5186),
.C(n_5150),
.Y(n_5755)
);

OA21x2_ASAP7_75t_L g5756 ( 
.A1(n_5396),
.A2(n_5037),
.B(n_5026),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5419),
.Y(n_5757)
);

BUFx2_ASAP7_75t_L g5758 ( 
.A(n_5435),
.Y(n_5758)
);

INVx2_ASAP7_75t_L g5759 ( 
.A(n_5401),
.Y(n_5759)
);

AO21x1_ASAP7_75t_SL g5760 ( 
.A1(n_5738),
.A2(n_5379),
.B(n_5368),
.Y(n_5760)
);

BUFx4f_ASAP7_75t_SL g5761 ( 
.A(n_5496),
.Y(n_5761)
);

INVx1_ASAP7_75t_L g5762 ( 
.A(n_5609),
.Y(n_5762)
);

HB1xp67_ASAP7_75t_L g5763 ( 
.A(n_5417),
.Y(n_5763)
);

INVx2_ASAP7_75t_L g5764 ( 
.A(n_5402),
.Y(n_5764)
);

OA21x2_ASAP7_75t_L g5765 ( 
.A1(n_5494),
.A2(n_5237),
.B(n_5215),
.Y(n_5765)
);

INVx2_ASAP7_75t_L g5766 ( 
.A(n_5630),
.Y(n_5766)
);

INVx2_ASAP7_75t_L g5767 ( 
.A(n_5650),
.Y(n_5767)
);

INVx2_ASAP7_75t_L g5768 ( 
.A(n_5660),
.Y(n_5768)
);

OR2x2_ASAP7_75t_L g5769 ( 
.A(n_5490),
.B(n_5294),
.Y(n_5769)
);

INVx2_ASAP7_75t_L g5770 ( 
.A(n_5505),
.Y(n_5770)
);

AND2x2_ASAP7_75t_L g5771 ( 
.A(n_5414),
.B(n_5325),
.Y(n_5771)
);

HB1xp67_ASAP7_75t_L g5772 ( 
.A(n_5417),
.Y(n_5772)
);

INVx1_ASAP7_75t_L g5773 ( 
.A(n_5609),
.Y(n_5773)
);

BUFx3_ASAP7_75t_L g5774 ( 
.A(n_5541),
.Y(n_5774)
);

INVx2_ASAP7_75t_L g5775 ( 
.A(n_5505),
.Y(n_5775)
);

INVx2_ASAP7_75t_L g5776 ( 
.A(n_5405),
.Y(n_5776)
);

BUFx10_ASAP7_75t_L g5777 ( 
.A(n_5499),
.Y(n_5777)
);

INVx2_ASAP7_75t_L g5778 ( 
.A(n_5405),
.Y(n_5778)
);

INVx2_ASAP7_75t_SL g5779 ( 
.A(n_5613),
.Y(n_5779)
);

INVx3_ASAP7_75t_L g5780 ( 
.A(n_5421),
.Y(n_5780)
);

INVx3_ASAP7_75t_L g5781 ( 
.A(n_5421),
.Y(n_5781)
);

INVx4_ASAP7_75t_L g5782 ( 
.A(n_5503),
.Y(n_5782)
);

AO21x2_ASAP7_75t_L g5783 ( 
.A1(n_5741),
.A2(n_5260),
.B(n_5282),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_5438),
.Y(n_5784)
);

INVxp67_ASAP7_75t_SL g5785 ( 
.A(n_5586),
.Y(n_5785)
);

AND2x4_ASAP7_75t_L g5786 ( 
.A(n_5399),
.B(n_5041),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_5438),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5408),
.Y(n_5788)
);

BUFx3_ASAP7_75t_L g5789 ( 
.A(n_5429),
.Y(n_5789)
);

HB1xp67_ASAP7_75t_L g5790 ( 
.A(n_5437),
.Y(n_5790)
);

INVx2_ASAP7_75t_L g5791 ( 
.A(n_5405),
.Y(n_5791)
);

AO21x2_ASAP7_75t_L g5792 ( 
.A1(n_5741),
.A2(n_5282),
.B(n_5172),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_5416),
.Y(n_5793)
);

OR2x6_ASAP7_75t_L g5794 ( 
.A(n_5399),
.B(n_5135),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_5420),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5422),
.Y(n_5796)
);

INVx2_ASAP7_75t_L g5797 ( 
.A(n_5723),
.Y(n_5797)
);

INVx2_ASAP7_75t_L g5798 ( 
.A(n_5733),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5448),
.Y(n_5799)
);

CKINVDCx5p33_ASAP7_75t_R g5800 ( 
.A(n_5525),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5731),
.Y(n_5801)
);

INVx2_ASAP7_75t_L g5802 ( 
.A(n_5737),
.Y(n_5802)
);

NAND2x1p5_ASAP7_75t_L g5803 ( 
.A(n_5698),
.B(n_5290),
.Y(n_5803)
);

INVx2_ASAP7_75t_L g5804 ( 
.A(n_5674),
.Y(n_5804)
);

BUFx3_ASAP7_75t_L g5805 ( 
.A(n_5545),
.Y(n_5805)
);

INVx1_ASAP7_75t_L g5806 ( 
.A(n_5449),
.Y(n_5806)
);

INVx2_ASAP7_75t_L g5807 ( 
.A(n_5680),
.Y(n_5807)
);

OAI21x1_ASAP7_75t_L g5808 ( 
.A1(n_5494),
.A2(n_5244),
.B(n_5229),
.Y(n_5808)
);

HB1xp67_ASAP7_75t_L g5809 ( 
.A(n_5428),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5681),
.Y(n_5810)
);

OAI21x1_ASAP7_75t_L g5811 ( 
.A1(n_5665),
.A2(n_5157),
.B(n_4993),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_5450),
.Y(n_5812)
);

NAND2xp5_ASAP7_75t_L g5813 ( 
.A(n_5586),
.B(n_5041),
.Y(n_5813)
);

HB1xp67_ASAP7_75t_L g5814 ( 
.A(n_5455),
.Y(n_5814)
);

AND2x2_ASAP7_75t_L g5815 ( 
.A(n_5439),
.B(n_5325),
.Y(n_5815)
);

INVx3_ASAP7_75t_L g5816 ( 
.A(n_5504),
.Y(n_5816)
);

INVx2_ASAP7_75t_L g5817 ( 
.A(n_5695),
.Y(n_5817)
);

INVx2_ASAP7_75t_SL g5818 ( 
.A(n_5627),
.Y(n_5818)
);

OAI21x1_ASAP7_75t_L g5819 ( 
.A1(n_5451),
.A2(n_5300),
.B(n_5158),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_5460),
.Y(n_5820)
);

CKINVDCx20_ASAP7_75t_R g5821 ( 
.A(n_5406),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5475),
.Y(n_5822)
);

AND2x2_ASAP7_75t_L g5823 ( 
.A(n_5441),
.B(n_5300),
.Y(n_5823)
);

INVx2_ASAP7_75t_L g5824 ( 
.A(n_5695),
.Y(n_5824)
);

INVx2_ASAP7_75t_L g5825 ( 
.A(n_5706),
.Y(n_5825)
);

AOI22xp5_ASAP7_75t_L g5826 ( 
.A1(n_5705),
.A2(n_5341),
.B1(n_5230),
.B2(n_5385),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5486),
.Y(n_5827)
);

OAI21x1_ASAP7_75t_L g5828 ( 
.A1(n_5539),
.A2(n_5304),
.B(n_5319),
.Y(n_5828)
);

INVx2_ASAP7_75t_L g5829 ( 
.A(n_5706),
.Y(n_5829)
);

INVx2_ASAP7_75t_L g5830 ( 
.A(n_5709),
.Y(n_5830)
);

INVx2_ASAP7_75t_L g5831 ( 
.A(n_5709),
.Y(n_5831)
);

INVx2_ASAP7_75t_L g5832 ( 
.A(n_5677),
.Y(n_5832)
);

OR2x2_ASAP7_75t_L g5833 ( 
.A(n_5626),
.B(n_5328),
.Y(n_5833)
);

INVx2_ASAP7_75t_SL g5834 ( 
.A(n_5627),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5513),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5515),
.Y(n_5836)
);

INVx1_ASAP7_75t_L g5837 ( 
.A(n_5520),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5523),
.Y(n_5838)
);

INVx1_ASAP7_75t_L g5839 ( 
.A(n_5530),
.Y(n_5839)
);

OAI21x1_ASAP7_75t_L g5840 ( 
.A1(n_5455),
.A2(n_5331),
.B(n_5323),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5532),
.Y(n_5841)
);

AOI22xp5_ASAP7_75t_L g5842 ( 
.A1(n_5705),
.A2(n_5230),
.B1(n_5046),
.B2(n_5236),
.Y(n_5842)
);

INVx2_ASAP7_75t_L g5843 ( 
.A(n_5691),
.Y(n_5843)
);

INVx2_ASAP7_75t_L g5844 ( 
.A(n_5716),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_5533),
.Y(n_5845)
);

AND2x2_ASAP7_75t_L g5846 ( 
.A(n_5400),
.B(n_5232),
.Y(n_5846)
);

AND2x2_ASAP7_75t_L g5847 ( 
.A(n_5407),
.B(n_5012),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5569),
.Y(n_5848)
);

AND2x2_ASAP7_75t_L g5849 ( 
.A(n_5504),
.B(n_5012),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_5578),
.Y(n_5850)
);

INVx1_ASAP7_75t_L g5851 ( 
.A(n_5582),
.Y(n_5851)
);

INVx1_ASAP7_75t_L g5852 ( 
.A(n_5588),
.Y(n_5852)
);

BUFx2_ASAP7_75t_L g5853 ( 
.A(n_5445),
.Y(n_5853)
);

INVx2_ASAP7_75t_L g5854 ( 
.A(n_5718),
.Y(n_5854)
);

AOI21x1_ASAP7_75t_L g5855 ( 
.A1(n_5600),
.A2(n_5702),
.B(n_5547),
.Y(n_5855)
);

AOI22xp33_ASAP7_75t_L g5856 ( 
.A1(n_5603),
.A2(n_5048),
.B1(n_5102),
.B2(n_5059),
.Y(n_5856)
);

INVx2_ASAP7_75t_L g5857 ( 
.A(n_5590),
.Y(n_5857)
);

INVx2_ASAP7_75t_L g5858 ( 
.A(n_5608),
.Y(n_5858)
);

AND2x2_ASAP7_75t_L g5859 ( 
.A(n_5447),
.B(n_5012),
.Y(n_5859)
);

AND2x2_ASAP7_75t_L g5860 ( 
.A(n_5457),
.B(n_5328),
.Y(n_5860)
);

INVx1_ASAP7_75t_L g5861 ( 
.A(n_5611),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_5509),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5629),
.Y(n_5863)
);

AO21x2_ASAP7_75t_L g5864 ( 
.A1(n_5742),
.A2(n_5279),
.B(n_5270),
.Y(n_5864)
);

INVx2_ASAP7_75t_L g5865 ( 
.A(n_5425),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5622),
.Y(n_5866)
);

INVx3_ASAP7_75t_L g5867 ( 
.A(n_5433),
.Y(n_5867)
);

INVx1_ASAP7_75t_SL g5868 ( 
.A(n_5479),
.Y(n_5868)
);

OR2x6_ASAP7_75t_L g5869 ( 
.A(n_5399),
.B(n_5194),
.Y(n_5869)
);

CKINVDCx14_ASAP7_75t_R g5870 ( 
.A(n_5654),
.Y(n_5870)
);

BUFx3_ASAP7_75t_L g5871 ( 
.A(n_5404),
.Y(n_5871)
);

AND2x4_ASAP7_75t_L g5872 ( 
.A(n_5579),
.B(n_5070),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5658),
.Y(n_5873)
);

INVx2_ASAP7_75t_L g5874 ( 
.A(n_5430),
.Y(n_5874)
);

OR2x2_ASAP7_75t_L g5875 ( 
.A(n_5463),
.B(n_5497),
.Y(n_5875)
);

INVx2_ASAP7_75t_L g5876 ( 
.A(n_5431),
.Y(n_5876)
);

OR2x2_ASAP7_75t_L g5877 ( 
.A(n_5463),
.B(n_5169),
.Y(n_5877)
);

AND2x4_ASAP7_75t_L g5878 ( 
.A(n_5579),
.B(n_5081),
.Y(n_5878)
);

AND2x4_ASAP7_75t_L g5879 ( 
.A(n_5483),
.B(n_5087),
.Y(n_5879)
);

AOI21x1_ASAP7_75t_L g5880 ( 
.A1(n_5683),
.A2(n_5313),
.B(n_5335),
.Y(n_5880)
);

AND2x4_ASAP7_75t_L g5881 ( 
.A(n_5483),
.B(n_5324),
.Y(n_5881)
);

BUFx2_ASAP7_75t_L g5882 ( 
.A(n_5445),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5617),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5566),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5573),
.Y(n_5885)
);

INVx2_ASAP7_75t_L g5886 ( 
.A(n_5440),
.Y(n_5886)
);

AO21x2_ASAP7_75t_L g5887 ( 
.A1(n_5742),
.A2(n_5076),
.B(n_5334),
.Y(n_5887)
);

INVx4_ASAP7_75t_SL g5888 ( 
.A(n_5698),
.Y(n_5888)
);

INVx1_ASAP7_75t_L g5889 ( 
.A(n_5550),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_5459),
.Y(n_5890)
);

INVx2_ASAP7_75t_L g5891 ( 
.A(n_5454),
.Y(n_5891)
);

INVx2_ASAP7_75t_L g5892 ( 
.A(n_5462),
.Y(n_5892)
);

NAND2x1p5_ASAP7_75t_L g5893 ( 
.A(n_5621),
.B(n_5290),
.Y(n_5893)
);

BUFx6f_ASAP7_75t_L g5894 ( 
.A(n_5560),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5501),
.Y(n_5895)
);

AND2x4_ASAP7_75t_L g5896 ( 
.A(n_5500),
.B(n_5338),
.Y(n_5896)
);

NAND2xp5_ASAP7_75t_L g5897 ( 
.A(n_5634),
.B(n_5265),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5599),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5487),
.Y(n_5899)
);

INVx2_ASAP7_75t_L g5900 ( 
.A(n_5464),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5471),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5512),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5522),
.Y(n_5903)
);

INVx1_ASAP7_75t_L g5904 ( 
.A(n_5524),
.Y(n_5904)
);

INVx1_ASAP7_75t_L g5905 ( 
.A(n_5526),
.Y(n_5905)
);

INVx2_ASAP7_75t_L g5906 ( 
.A(n_5535),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5542),
.Y(n_5907)
);

AO21x2_ASAP7_75t_L g5908 ( 
.A1(n_5446),
.A2(n_5196),
.B(n_5201),
.Y(n_5908)
);

AND2x2_ASAP7_75t_L g5909 ( 
.A(n_5432),
.B(n_5169),
.Y(n_5909)
);

INVx5_ASAP7_75t_L g5910 ( 
.A(n_5701),
.Y(n_5910)
);

OR2x2_ASAP7_75t_L g5911 ( 
.A(n_5634),
.B(n_5144),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5552),
.Y(n_5912)
);

INVx2_ASAP7_75t_L g5913 ( 
.A(n_5556),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5574),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_5615),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5693),
.Y(n_5916)
);

INVx2_ASAP7_75t_SL g5917 ( 
.A(n_5670),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5697),
.Y(n_5918)
);

INVx2_ASAP7_75t_SL g5919 ( 
.A(n_5595),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5707),
.Y(n_5920)
);

INVx3_ASAP7_75t_L g5921 ( 
.A(n_5433),
.Y(n_5921)
);

AND2x2_ASAP7_75t_L g5922 ( 
.A(n_5534),
.B(n_5273),
.Y(n_5922)
);

INVx3_ASAP7_75t_L g5923 ( 
.A(n_5557),
.Y(n_5923)
);

BUFx2_ASAP7_75t_L g5924 ( 
.A(n_5557),
.Y(n_5924)
);

INVx1_ASAP7_75t_L g5925 ( 
.A(n_5707),
.Y(n_5925)
);

AND2x2_ASAP7_75t_L g5926 ( 
.A(n_5452),
.B(n_5151),
.Y(n_5926)
);

OA21x2_ASAP7_75t_L g5927 ( 
.A1(n_5446),
.A2(n_5387),
.B(n_5223),
.Y(n_5927)
);

OAI22xp33_ASAP7_75t_L g5928 ( 
.A1(n_5397),
.A2(n_5393),
.B1(n_5384),
.B2(n_5243),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_5633),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5704),
.Y(n_5930)
);

HB1xp67_ASAP7_75t_L g5931 ( 
.A(n_5510),
.Y(n_5931)
);

OA21x2_ASAP7_75t_L g5932 ( 
.A1(n_5424),
.A2(n_5079),
.B(n_5089),
.Y(n_5932)
);

INVx2_ASAP7_75t_L g5933 ( 
.A(n_5708),
.Y(n_5933)
);

OAI21x1_ASAP7_75t_L g5934 ( 
.A1(n_5575),
.A2(n_5531),
.B(n_5444),
.Y(n_5934)
);

CKINVDCx6p67_ASAP7_75t_R g5935 ( 
.A(n_5528),
.Y(n_5935)
);

BUFx3_ASAP7_75t_L g5936 ( 
.A(n_5725),
.Y(n_5936)
);

INVx1_ASAP7_75t_L g5937 ( 
.A(n_5648),
.Y(n_5937)
);

INVx1_ASAP7_75t_L g5938 ( 
.A(n_5649),
.Y(n_5938)
);

OR2x2_ASAP7_75t_L g5939 ( 
.A(n_5510),
.B(n_5356),
.Y(n_5939)
);

INVx1_ASAP7_75t_L g5940 ( 
.A(n_5423),
.Y(n_5940)
);

INVx2_ASAP7_75t_L g5941 ( 
.A(n_5711),
.Y(n_5941)
);

OR2x6_ASAP7_75t_L g5942 ( 
.A(n_5482),
.B(n_5156),
.Y(n_5942)
);

AND2x4_ASAP7_75t_L g5943 ( 
.A(n_5500),
.B(n_5246),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_5397),
.Y(n_5944)
);

AND2x2_ASAP7_75t_L g5945 ( 
.A(n_5452),
.B(n_5392),
.Y(n_5945)
);

INVx2_ASAP7_75t_L g5946 ( 
.A(n_5740),
.Y(n_5946)
);

OAI21x1_ASAP7_75t_L g5947 ( 
.A1(n_5540),
.A2(n_5367),
.B(n_5358),
.Y(n_5947)
);

HB1xp67_ASAP7_75t_L g5948 ( 
.A(n_5508),
.Y(n_5948)
);

HB1xp67_ASAP7_75t_L g5949 ( 
.A(n_5508),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5498),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5632),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5635),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5722),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5722),
.Y(n_5954)
);

HB1xp67_ASAP7_75t_L g5955 ( 
.A(n_5584),
.Y(n_5955)
);

INVx1_ASAP7_75t_L g5956 ( 
.A(n_5495),
.Y(n_5956)
);

AND2x4_ASAP7_75t_L g5957 ( 
.A(n_5506),
.B(n_5066),
.Y(n_5957)
);

INVx2_ASAP7_75t_L g5958 ( 
.A(n_5703),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5694),
.Y(n_5959)
);

NAND2xp5_ASAP7_75t_L g5960 ( 
.A(n_5559),
.B(n_5123),
.Y(n_5960)
);

INVx1_ASAP7_75t_L g5961 ( 
.A(n_5507),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5581),
.Y(n_5962)
);

INVx1_ASAP7_75t_L g5963 ( 
.A(n_5506),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5584),
.Y(n_5964)
);

OAI21x1_ASAP7_75t_L g5965 ( 
.A1(n_5540),
.A2(n_5249),
.B(n_5277),
.Y(n_5965)
);

AND2x2_ASAP7_75t_L g5966 ( 
.A(n_5543),
.B(n_5077),
.Y(n_5966)
);

AND2x2_ASAP7_75t_L g5967 ( 
.A(n_5485),
.B(n_5077),
.Y(n_5967)
);

AND2x2_ASAP7_75t_L g5968 ( 
.A(n_5555),
.B(n_5077),
.Y(n_5968)
);

INVx2_ASAP7_75t_L g5969 ( 
.A(n_5580),
.Y(n_5969)
);

AND2x4_ASAP7_75t_L g5970 ( 
.A(n_5409),
.B(n_5356),
.Y(n_5970)
);

BUFx2_ASAP7_75t_L g5971 ( 
.A(n_5636),
.Y(n_5971)
);

AO21x2_ASAP7_75t_L g5972 ( 
.A1(n_5639),
.A2(n_5112),
.B(n_5078),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5594),
.Y(n_5973)
);

INVx3_ASAP7_75t_L g5974 ( 
.A(n_5642),
.Y(n_5974)
);

INVx1_ASAP7_75t_L g5975 ( 
.A(n_5594),
.Y(n_5975)
);

BUFx3_ASAP7_75t_L g5976 ( 
.A(n_5607),
.Y(n_5976)
);

INVx2_ASAP7_75t_L g5977 ( 
.A(n_5580),
.Y(n_5977)
);

HB1xp67_ASAP7_75t_L g5978 ( 
.A(n_5656),
.Y(n_5978)
);

INVx3_ASAP7_75t_L g5979 ( 
.A(n_5728),
.Y(n_5979)
);

BUFx10_ASAP7_75t_L g5980 ( 
.A(n_5537),
.Y(n_5980)
);

OAI21x1_ASAP7_75t_L g5981 ( 
.A1(n_5564),
.A2(n_5202),
.B(n_5166),
.Y(n_5981)
);

AND2x4_ASAP7_75t_L g5982 ( 
.A(n_5468),
.B(n_5356),
.Y(n_5982)
);

INVx2_ASAP7_75t_L g5983 ( 
.A(n_5580),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5468),
.Y(n_5984)
);

INVx3_ASAP7_75t_L g5985 ( 
.A(n_5728),
.Y(n_5985)
);

INVx3_ASAP7_75t_L g5986 ( 
.A(n_5598),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5468),
.Y(n_5987)
);

CKINVDCx8_ASAP7_75t_R g5988 ( 
.A(n_5403),
.Y(n_5988)
);

INVx6_ASAP7_75t_L g5989 ( 
.A(n_5720),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5469),
.Y(n_5990)
);

BUFx2_ASAP7_75t_L g5991 ( 
.A(n_5659),
.Y(n_5991)
);

INVx2_ASAP7_75t_L g5992 ( 
.A(n_5589),
.Y(n_5992)
);

INVx2_ASAP7_75t_L g5993 ( 
.A(n_5577),
.Y(n_5993)
);

NAND2xp5_ASAP7_75t_L g5994 ( 
.A(n_5511),
.B(n_5090),
.Y(n_5994)
);

INVx2_ASAP7_75t_SL g5995 ( 
.A(n_5598),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5469),
.Y(n_5996)
);

INVx1_ASAP7_75t_L g5997 ( 
.A(n_5469),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5603),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5676),
.Y(n_5999)
);

BUFx6f_ASAP7_75t_L g6000 ( 
.A(n_5442),
.Y(n_6000)
);

NOR2xp33_ASAP7_75t_L g6001 ( 
.A(n_5410),
.B(n_134),
.Y(n_6001)
);

CKINVDCx5p33_ASAP7_75t_R g6002 ( 
.A(n_5558),
.Y(n_6002)
);

INVx3_ASAP7_75t_L g6003 ( 
.A(n_5553),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5567),
.Y(n_6004)
);

NAND2xp5_ASAP7_75t_L g6005 ( 
.A(n_5511),
.B(n_5113),
.Y(n_6005)
);

INVx3_ASAP7_75t_L g6006 ( 
.A(n_5553),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5616),
.Y(n_6007)
);

AND2x2_ASAP7_75t_L g6008 ( 
.A(n_5652),
.B(n_135),
.Y(n_6008)
);

NAND2xp5_ASAP7_75t_L g6009 ( 
.A(n_5616),
.B(n_5019),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5527),
.Y(n_6010)
);

INVx1_ASAP7_75t_L g6011 ( 
.A(n_5527),
.Y(n_6011)
);

AO21x1_ASAP7_75t_L g6012 ( 
.A1(n_5644),
.A2(n_5226),
.B(n_5247),
.Y(n_6012)
);

INVx2_ASAP7_75t_L g6013 ( 
.A(n_5721),
.Y(n_6013)
);

INVx2_ASAP7_75t_L g6014 ( 
.A(n_5553),
.Y(n_6014)
);

INVx1_ASAP7_75t_L g6015 ( 
.A(n_5516),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5568),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5568),
.Y(n_6017)
);

NAND2xp5_ASAP7_75t_L g6018 ( 
.A(n_5436),
.B(n_5038),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5568),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5625),
.Y(n_6020)
);

BUFx3_ASAP7_75t_L g6021 ( 
.A(n_5565),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_5482),
.Y(n_6022)
);

INVx2_ASAP7_75t_L g6023 ( 
.A(n_5610),
.Y(n_6023)
);

INVx1_ASAP7_75t_L g6024 ( 
.A(n_5482),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5610),
.Y(n_6025)
);

INVx3_ASAP7_75t_L g6026 ( 
.A(n_5664),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5664),
.B(n_135),
.Y(n_6027)
);

INVx3_ASAP7_75t_L g6028 ( 
.A(n_5489),
.Y(n_6028)
);

INVx1_ASAP7_75t_L g6029 ( 
.A(n_5857),
.Y(n_6029)
);

INVx2_ASAP7_75t_L g6030 ( 
.A(n_5953),
.Y(n_6030)
);

AOI22xp33_ASAP7_75t_L g6031 ( 
.A1(n_5940),
.A2(n_5689),
.B1(n_5690),
.B2(n_5673),
.Y(n_6031)
);

OAI221xp5_ASAP7_75t_L g6032 ( 
.A1(n_5785),
.A2(n_5453),
.B1(n_5679),
.B2(n_5646),
.C(n_5478),
.Y(n_6032)
);

INVx2_ASAP7_75t_L g6033 ( 
.A(n_5954),
.Y(n_6033)
);

AOI22xp33_ASAP7_75t_L g6034 ( 
.A1(n_5998),
.A2(n_5671),
.B1(n_5548),
.B2(n_5563),
.Y(n_6034)
);

OAI22xp5_ASAP7_75t_L g6035 ( 
.A1(n_6007),
.A2(n_5491),
.B1(n_5473),
.B2(n_5492),
.Y(n_6035)
);

AOI21xp33_ASAP7_75t_L g6036 ( 
.A1(n_5785),
.A2(n_5576),
.B(n_5618),
.Y(n_6036)
);

OAI21x1_ASAP7_75t_L g6037 ( 
.A1(n_5855),
.A2(n_5456),
.B(n_5536),
.Y(n_6037)
);

NAND2xp5_ASAP7_75t_L g6038 ( 
.A(n_5763),
.B(n_5772),
.Y(n_6038)
);

A2O1A1Ixp33_ASAP7_75t_L g6039 ( 
.A1(n_5847),
.A2(n_5585),
.B(n_5647),
.C(n_5554),
.Y(n_6039)
);

INVx3_ASAP7_75t_L g6040 ( 
.A(n_5881),
.Y(n_6040)
);

OAI221xp5_ASAP7_75t_L g6041 ( 
.A1(n_5813),
.A2(n_5944),
.B1(n_5679),
.B2(n_5825),
.C(n_5824),
.Y(n_6041)
);

AOI22xp33_ASAP7_75t_L g6042 ( 
.A1(n_6020),
.A2(n_5651),
.B1(n_5443),
.B2(n_5427),
.Y(n_6042)
);

AND2x4_ASAP7_75t_L g6043 ( 
.A(n_5888),
.B(n_5517),
.Y(n_6043)
);

AO31x2_ASAP7_75t_L g6044 ( 
.A1(n_5776),
.A2(n_5791),
.A3(n_5778),
.B(n_5817),
.Y(n_6044)
);

INVx2_ASAP7_75t_L g6045 ( 
.A(n_5909),
.Y(n_6045)
);

AOI22xp5_ASAP7_75t_L g6046 ( 
.A1(n_6012),
.A2(n_5427),
.B1(n_5571),
.B2(n_5544),
.Y(n_6046)
);

OAI22xp5_ASAP7_75t_L g6047 ( 
.A1(n_5744),
.A2(n_5571),
.B1(n_5536),
.B2(n_5398),
.Y(n_6047)
);

OAI221xp5_ASAP7_75t_L g6048 ( 
.A1(n_5817),
.A2(n_5458),
.B1(n_5514),
.B2(n_5596),
.C(n_5686),
.Y(n_6048)
);

OAI22xp5_ASAP7_75t_L g6049 ( 
.A1(n_5744),
.A2(n_5461),
.B1(n_5480),
.B2(n_5477),
.Y(n_6049)
);

OAI221xp5_ASAP7_75t_L g6050 ( 
.A1(n_5824),
.A2(n_5667),
.B1(n_5570),
.B2(n_5655),
.C(n_5619),
.Y(n_6050)
);

AND2x4_ASAP7_75t_L g6051 ( 
.A(n_5888),
.B(n_5517),
.Y(n_6051)
);

OR2x2_ASAP7_75t_L g6052 ( 
.A(n_5875),
.B(n_5587),
.Y(n_6052)
);

INVx2_ASAP7_75t_L g6053 ( 
.A(n_5857),
.Y(n_6053)
);

OAI221xp5_ASAP7_75t_SL g6054 ( 
.A1(n_5928),
.A2(n_5663),
.B1(n_5717),
.B2(n_5732),
.C(n_5624),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5858),
.Y(n_6055)
);

OR2x2_ASAP7_75t_L g6056 ( 
.A(n_5770),
.B(n_5465),
.Y(n_6056)
);

AOI221xp5_ASAP7_75t_L g6057 ( 
.A1(n_5763),
.A2(n_5618),
.B1(n_5619),
.B2(n_5657),
.C(n_5729),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5858),
.Y(n_6058)
);

AOI22xp33_ASAP7_75t_L g6059 ( 
.A1(n_5797),
.A2(n_5612),
.B1(n_5614),
.B2(n_5413),
.Y(n_6059)
);

AOI22xp33_ASAP7_75t_L g6060 ( 
.A1(n_5797),
.A2(n_5614),
.B1(n_5612),
.B2(n_5518),
.Y(n_6060)
);

BUFx2_ASAP7_75t_L g6061 ( 
.A(n_5936),
.Y(n_6061)
);

OAI22xp5_ASAP7_75t_L g6062 ( 
.A1(n_6009),
.A2(n_5477),
.B1(n_5549),
.B2(n_5546),
.Y(n_6062)
);

BUFx3_ASAP7_75t_L g6063 ( 
.A(n_5789),
.Y(n_6063)
);

INVx2_ASAP7_75t_L g6064 ( 
.A(n_5939),
.Y(n_6064)
);

INVx2_ASAP7_75t_L g6065 ( 
.A(n_5770),
.Y(n_6065)
);

AOI21xp5_ASAP7_75t_L g6066 ( 
.A1(n_5928),
.A2(n_5994),
.B(n_6015),
.Y(n_6066)
);

AOI21xp5_ASAP7_75t_L g6067 ( 
.A1(n_6005),
.A2(n_5592),
.B(n_5549),
.Y(n_6067)
);

AOI22xp33_ASAP7_75t_L g6068 ( 
.A1(n_5798),
.A2(n_5628),
.B1(n_5684),
.B2(n_5710),
.Y(n_6068)
);

OAI211xp5_ASAP7_75t_L g6069 ( 
.A1(n_5955),
.A2(n_5713),
.B(n_5502),
.C(n_5620),
.Y(n_6069)
);

NOR2xp33_ASAP7_75t_L g6070 ( 
.A(n_5782),
.B(n_5415),
.Y(n_6070)
);

INVx3_ASAP7_75t_L g6071 ( 
.A(n_5881),
.Y(n_6071)
);

CKINVDCx20_ASAP7_75t_R g6072 ( 
.A(n_5761),
.Y(n_6072)
);

AOI21x1_ASAP7_75t_L g6073 ( 
.A1(n_5931),
.A2(n_5641),
.B(n_5606),
.Y(n_6073)
);

AOI221xp5_ASAP7_75t_L g6074 ( 
.A1(n_5772),
.A2(n_5657),
.B1(n_5829),
.B2(n_5830),
.C(n_5825),
.Y(n_6074)
);

AOI22xp33_ASAP7_75t_SL g6075 ( 
.A1(n_5846),
.A2(n_5561),
.B1(n_5730),
.B2(n_5672),
.Y(n_6075)
);

AOI21xp5_ASAP7_75t_L g6076 ( 
.A1(n_5869),
.A2(n_5470),
.B(n_5466),
.Y(n_6076)
);

NOR2xp33_ASAP7_75t_L g6077 ( 
.A(n_5782),
.B(n_5442),
.Y(n_6077)
);

OAI22xp5_ASAP7_75t_L g6078 ( 
.A1(n_5856),
.A2(n_5729),
.B1(n_5684),
.B2(n_5712),
.Y(n_6078)
);

AOI22xp33_ASAP7_75t_L g6079 ( 
.A1(n_5798),
.A2(n_5628),
.B1(n_5712),
.B2(n_5710),
.Y(n_6079)
);

NAND2xp5_ASAP7_75t_L g6080 ( 
.A(n_5784),
.B(n_5714),
.Y(n_6080)
);

AOI22xp33_ASAP7_75t_L g6081 ( 
.A1(n_5918),
.A2(n_5727),
.B1(n_5696),
.B2(n_5688),
.Y(n_6081)
);

BUFx6f_ASAP7_75t_L g6082 ( 
.A(n_5789),
.Y(n_6082)
);

AND2x2_ASAP7_75t_L g6083 ( 
.A(n_5816),
.B(n_5489),
.Y(n_6083)
);

AOI22xp33_ASAP7_75t_SL g6084 ( 
.A1(n_5849),
.A2(n_5561),
.B1(n_5730),
.B2(n_5727),
.Y(n_6084)
);

AND2x4_ASAP7_75t_L g6085 ( 
.A(n_5888),
.B(n_5529),
.Y(n_6085)
);

AOI22xp33_ASAP7_75t_L g6086 ( 
.A1(n_5760),
.A2(n_5696),
.B1(n_5734),
.B2(n_5688),
.Y(n_6086)
);

AOI22xp33_ASAP7_75t_L g6087 ( 
.A1(n_6018),
.A2(n_5734),
.B1(n_5470),
.B2(n_5467),
.Y(n_6087)
);

AND2x2_ASAP7_75t_L g6088 ( 
.A(n_5816),
.B(n_5591),
.Y(n_6088)
);

AOI22xp33_ASAP7_75t_SL g6089 ( 
.A1(n_5859),
.A2(n_5643),
.B1(n_5662),
.B2(n_5669),
.Y(n_6089)
);

OAI22xp5_ASAP7_75t_L g6090 ( 
.A1(n_5826),
.A2(n_6004),
.B1(n_5955),
.B2(n_5803),
.Y(n_6090)
);

OAI22xp33_ASAP7_75t_L g6091 ( 
.A1(n_5942),
.A2(n_5583),
.B1(n_5631),
.B2(n_5645),
.Y(n_6091)
);

OR2x2_ASAP7_75t_L g6092 ( 
.A(n_5775),
.B(n_5593),
.Y(n_6092)
);

CKINVDCx5p33_ASAP7_75t_R g6093 ( 
.A(n_5800),
.Y(n_6093)
);

OAI221xp5_ASAP7_75t_L g6094 ( 
.A1(n_5829),
.A2(n_5476),
.B1(n_5474),
.B2(n_5472),
.C(n_5481),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_5762),
.Y(n_6095)
);

NOR2x1_ASAP7_75t_SL g6096 ( 
.A(n_5794),
.B(n_5637),
.Y(n_6096)
);

OAI211xp5_ASAP7_75t_SL g6097 ( 
.A1(n_5951),
.A2(n_5715),
.B(n_5736),
.C(n_5484),
.Y(n_6097)
);

OAI22xp5_ASAP7_75t_L g6098 ( 
.A1(n_5803),
.A2(n_5666),
.B1(n_5675),
.B2(n_5668),
.Y(n_6098)
);

OAI211xp5_ASAP7_75t_L g6099 ( 
.A1(n_5931),
.A2(n_5715),
.B(n_5736),
.C(n_5602),
.Y(n_6099)
);

OAI22xp5_ASAP7_75t_L g6100 ( 
.A1(n_5869),
.A2(n_5597),
.B1(n_5661),
.B2(n_5572),
.Y(n_6100)
);

INVx2_ASAP7_75t_L g6101 ( 
.A(n_5775),
.Y(n_6101)
);

AOI22xp33_ASAP7_75t_L g6102 ( 
.A1(n_5972),
.A2(n_5519),
.B1(n_5493),
.B2(n_5562),
.Y(n_6102)
);

AOI22xp33_ASAP7_75t_L g6103 ( 
.A1(n_5972),
.A2(n_5743),
.B1(n_5687),
.B2(n_5692),
.Y(n_6103)
);

INVx2_ASAP7_75t_L g6104 ( 
.A(n_5865),
.Y(n_6104)
);

OAI211xp5_ASAP7_75t_L g6105 ( 
.A1(n_6001),
.A2(n_5739),
.B(n_5699),
.C(n_5724),
.Y(n_6105)
);

NOR2xp33_ASAP7_75t_L g6106 ( 
.A(n_5752),
.B(n_5597),
.Y(n_6106)
);

OAI221xp5_ASAP7_75t_L g6107 ( 
.A1(n_5830),
.A2(n_5638),
.B1(n_5538),
.B2(n_5551),
.C(n_5521),
.Y(n_6107)
);

OAI22xp33_ASAP7_75t_L g6108 ( 
.A1(n_5942),
.A2(n_5601),
.B1(n_5669),
.B2(n_5653),
.Y(n_6108)
);

INVx2_ASAP7_75t_L g6109 ( 
.A(n_5865),
.Y(n_6109)
);

AOI211xp5_ASAP7_75t_L g6110 ( 
.A1(n_6001),
.A2(n_5755),
.B(n_5842),
.C(n_5964),
.Y(n_6110)
);

OAI22x1_ASAP7_75t_L g6111 ( 
.A1(n_5999),
.A2(n_5700),
.B1(n_5678),
.B2(n_5726),
.Y(n_6111)
);

AOI22xp33_ASAP7_75t_L g6112 ( 
.A1(n_5831),
.A2(n_5605),
.B1(n_5488),
.B2(n_5735),
.Y(n_6112)
);

HB1xp67_ASAP7_75t_L g6113 ( 
.A(n_5790),
.Y(n_6113)
);

OAI211xp5_ASAP7_75t_L g6114 ( 
.A1(n_5809),
.A2(n_5755),
.B(n_5960),
.C(n_5853),
.Y(n_6114)
);

INVx1_ASAP7_75t_L g6115 ( 
.A(n_5773),
.Y(n_6115)
);

INVx2_ASAP7_75t_L g6116 ( 
.A(n_5874),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5790),
.Y(n_6117)
);

AOI22xp33_ASAP7_75t_L g6118 ( 
.A1(n_5831),
.A2(n_5640),
.B1(n_5682),
.B2(n_5623),
.Y(n_6118)
);

AOI22xp33_ASAP7_75t_L g6119 ( 
.A1(n_5856),
.A2(n_5719),
.B1(n_5604),
.B2(n_2461),
.Y(n_6119)
);

AOI211xp5_ASAP7_75t_L g6120 ( 
.A1(n_5973),
.A2(n_5061),
.B(n_5062),
.C(n_5044),
.Y(n_6120)
);

AOI22xp33_ASAP7_75t_L g6121 ( 
.A1(n_5942),
.A2(n_2461),
.B1(n_2463),
.B2(n_2456),
.Y(n_6121)
);

INVx3_ASAP7_75t_L g6122 ( 
.A(n_5881),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5799),
.Y(n_6123)
);

AOI21xp33_ASAP7_75t_L g6124 ( 
.A1(n_5948),
.A2(n_5224),
.B(n_5275),
.Y(n_6124)
);

OAI22xp5_ASAP7_75t_L g6125 ( 
.A1(n_5869),
.A2(n_140),
.B1(n_136),
.B2(n_138),
.Y(n_6125)
);

INVx2_ASAP7_75t_L g6126 ( 
.A(n_5874),
.Y(n_6126)
);

BUFx3_ASAP7_75t_L g6127 ( 
.A(n_5761),
.Y(n_6127)
);

NOR2xp33_ASAP7_75t_L g6128 ( 
.A(n_5752),
.B(n_141),
.Y(n_6128)
);

INVx1_ASAP7_75t_L g6129 ( 
.A(n_5806),
.Y(n_6129)
);

OAI221xp5_ASAP7_75t_L g6130 ( 
.A1(n_5745),
.A2(n_2469),
.B1(n_2474),
.B2(n_2464),
.C(n_2463),
.Y(n_6130)
);

AOI221xp5_ASAP7_75t_L g6131 ( 
.A1(n_5897),
.A2(n_5814),
.B1(n_5916),
.B2(n_5791),
.C(n_5778),
.Y(n_6131)
);

AOI22xp33_ASAP7_75t_L g6132 ( 
.A1(n_5887),
.A2(n_2469),
.B1(n_2474),
.B2(n_2464),
.Y(n_6132)
);

AOI221xp5_ASAP7_75t_L g6133 ( 
.A1(n_5814),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.C(n_144),
.Y(n_6133)
);

OAI22xp5_ASAP7_75t_L g6134 ( 
.A1(n_5975),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_5966),
.B(n_146),
.Y(n_6135)
);

AOI22xp33_ASAP7_75t_L g6136 ( 
.A1(n_5887),
.A2(n_2484),
.B1(n_2478),
.B2(n_2099),
.Y(n_6136)
);

OAI22xp33_ASAP7_75t_L g6137 ( 
.A1(n_5794),
.A2(n_150),
.B1(n_151),
.B2(n_149),
.Y(n_6137)
);

AOI22xp33_ASAP7_75t_L g6138 ( 
.A1(n_5898),
.A2(n_5863),
.B1(n_5890),
.B2(n_5984),
.Y(n_6138)
);

OR2x6_ASAP7_75t_L g6139 ( 
.A(n_5794),
.B(n_2478),
.Y(n_6139)
);

NAND2xp5_ASAP7_75t_L g6140 ( 
.A(n_5787),
.B(n_147),
.Y(n_6140)
);

AND2x2_ASAP7_75t_L g6141 ( 
.A(n_5968),
.B(n_5771),
.Y(n_6141)
);

AOI21xp33_ASAP7_75t_L g6142 ( 
.A1(n_5948),
.A2(n_147),
.B(n_149),
.Y(n_6142)
);

AOI22xp33_ASAP7_75t_L g6143 ( 
.A1(n_5987),
.A2(n_2484),
.B1(n_2099),
.B2(n_2109),
.Y(n_6143)
);

INVx5_ASAP7_75t_SL g6144 ( 
.A(n_5935),
.Y(n_6144)
);

NAND2xp5_ASAP7_75t_L g6145 ( 
.A(n_5746),
.B(n_152),
.Y(n_6145)
);

AOI22xp33_ASAP7_75t_SL g6146 ( 
.A1(n_5908),
.A2(n_161),
.B1(n_169),
.B2(n_152),
.Y(n_6146)
);

AND2x2_ASAP7_75t_L g6147 ( 
.A(n_5815),
.B(n_153),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_5812),
.Y(n_6148)
);

AND2x2_ASAP7_75t_L g6149 ( 
.A(n_5991),
.B(n_154),
.Y(n_6149)
);

OAI22xp33_ASAP7_75t_L g6150 ( 
.A1(n_5911),
.A2(n_156),
.B1(n_157),
.B2(n_155),
.Y(n_6150)
);

INVx2_ASAP7_75t_L g6151 ( 
.A(n_5876),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_5820),
.Y(n_6152)
);

INVx2_ASAP7_75t_L g6153 ( 
.A(n_5876),
.Y(n_6153)
);

HB1xp67_ASAP7_75t_L g6154 ( 
.A(n_5746),
.Y(n_6154)
);

AOI22xp33_ASAP7_75t_L g6155 ( 
.A1(n_5990),
.A2(n_2099),
.B1(n_2109),
.B2(n_2082),
.Y(n_6155)
);

AND2x2_ASAP7_75t_L g6156 ( 
.A(n_5963),
.B(n_154),
.Y(n_6156)
);

OAI21x1_ASAP7_75t_L g6157 ( 
.A1(n_5776),
.A2(n_2587),
.B(n_2428),
.Y(n_6157)
);

AND2x2_ASAP7_75t_L g6158 ( 
.A(n_5986),
.B(n_155),
.Y(n_6158)
);

AOI22xp33_ASAP7_75t_L g6159 ( 
.A1(n_5996),
.A2(n_2099),
.B1(n_2109),
.B2(n_2082),
.Y(n_6159)
);

AOI22xp33_ASAP7_75t_L g6160 ( 
.A1(n_5997),
.A2(n_5883),
.B1(n_6023),
.B2(n_5786),
.Y(n_6160)
);

OR2x2_ASAP7_75t_L g6161 ( 
.A(n_5866),
.B(n_156),
.Y(n_6161)
);

OAI22xp5_ASAP7_75t_L g6162 ( 
.A1(n_5818),
.A2(n_161),
.B1(n_158),
.B2(n_160),
.Y(n_6162)
);

AOI22xp33_ASAP7_75t_L g6163 ( 
.A1(n_6023),
.A2(n_2099),
.B1(n_2109),
.B2(n_2082),
.Y(n_6163)
);

INVx8_ASAP7_75t_L g6164 ( 
.A(n_5910),
.Y(n_6164)
);

HB1xp67_ASAP7_75t_SL g6165 ( 
.A(n_6021),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_5822),
.Y(n_6166)
);

AOI21xp5_ASAP7_75t_L g6167 ( 
.A1(n_5751),
.A2(n_160),
.B(n_162),
.Y(n_6167)
);

OAI21x1_ASAP7_75t_L g6168 ( 
.A1(n_5880),
.A2(n_2587),
.B(n_2429),
.Y(n_6168)
);

OAI22xp5_ASAP7_75t_L g6169 ( 
.A1(n_5834),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_6169)
);

INVx1_ASAP7_75t_L g6170 ( 
.A(n_5827),
.Y(n_6170)
);

AOI22xp33_ASAP7_75t_SL g6171 ( 
.A1(n_5908),
.A2(n_171),
.B1(n_180),
.B2(n_163),
.Y(n_6171)
);

OR2x2_ASAP7_75t_L g6172 ( 
.A(n_5750),
.B(n_164),
.Y(n_6172)
);

A2O1A1Ixp33_ASAP7_75t_L g6173 ( 
.A1(n_6021),
.A2(n_174),
.B(n_183),
.C(n_165),
.Y(n_6173)
);

OAI22xp33_ASAP7_75t_L g6174 ( 
.A1(n_5769),
.A2(n_5894),
.B1(n_5949),
.B2(n_6022),
.Y(n_6174)
);

OAI22xp5_ASAP7_75t_L g6175 ( 
.A1(n_6024),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_6175)
);

AOI21xp5_ASAP7_75t_SL g6176 ( 
.A1(n_5894),
.A2(n_166),
.B(n_168),
.Y(n_6176)
);

INVx3_ASAP7_75t_L g6177 ( 
.A(n_5894),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_5835),
.Y(n_6178)
);

AOI21xp5_ASAP7_75t_L g6179 ( 
.A1(n_5957),
.A2(n_169),
.B(n_170),
.Y(n_6179)
);

OAI221xp5_ASAP7_75t_L g6180 ( 
.A1(n_5877),
.A2(n_2430),
.B1(n_2432),
.B2(n_2429),
.C(n_2422),
.Y(n_6180)
);

NAND2xp5_ASAP7_75t_L g6181 ( 
.A(n_5809),
.B(n_171),
.Y(n_6181)
);

AND2x2_ASAP7_75t_L g6182 ( 
.A(n_5986),
.B(n_173),
.Y(n_6182)
);

AOI22xp33_ASAP7_75t_L g6183 ( 
.A1(n_5786),
.A2(n_2109),
.B1(n_2111),
.B2(n_2082),
.Y(n_6183)
);

AOI22xp33_ASAP7_75t_L g6184 ( 
.A1(n_5786),
.A2(n_2111),
.B1(n_2122),
.B2(n_2082),
.Y(n_6184)
);

NAND2xp33_ASAP7_75t_R g6185 ( 
.A(n_5800),
.B(n_176),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5836),
.Y(n_6186)
);

INVx1_ASAP7_75t_L g6187 ( 
.A(n_5837),
.Y(n_6187)
);

AND2x4_ASAP7_75t_L g6188 ( 
.A(n_5957),
.B(n_175),
.Y(n_6188)
);

OR2x2_ASAP7_75t_L g6189 ( 
.A(n_5862),
.B(n_5895),
.Y(n_6189)
);

OAI211xp5_ASAP7_75t_L g6190 ( 
.A1(n_5758),
.A2(n_178),
.B(n_175),
.C(n_177),
.Y(n_6190)
);

AND2x2_ASAP7_75t_L g6191 ( 
.A(n_5882),
.B(n_177),
.Y(n_6191)
);

OAI211xp5_ASAP7_75t_SL g6192 ( 
.A1(n_5952),
.A2(n_181),
.B(n_178),
.C(n_179),
.Y(n_6192)
);

AOI222xp33_ASAP7_75t_L g6193 ( 
.A1(n_5873),
.A2(n_185),
.B1(n_187),
.B2(n_182),
.C1(n_184),
.C2(n_186),
.Y(n_6193)
);

INVx2_ASAP7_75t_L g6194 ( 
.A(n_5886),
.Y(n_6194)
);

AOI222xp33_ASAP7_75t_L g6195 ( 
.A1(n_6008),
.A2(n_188),
.B1(n_190),
.B2(n_182),
.C1(n_185),
.C2(n_189),
.Y(n_6195)
);

AOI22xp33_ASAP7_75t_L g6196 ( 
.A1(n_5860),
.A2(n_2122),
.B1(n_2124),
.B2(n_2111),
.Y(n_6196)
);

AOI221xp5_ASAP7_75t_L g6197 ( 
.A1(n_5949),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_191),
.Y(n_6197)
);

AOI22xp33_ASAP7_75t_SL g6198 ( 
.A1(n_5932),
.A2(n_194),
.B1(n_191),
.B2(n_193),
.Y(n_6198)
);

INVx2_ASAP7_75t_L g6199 ( 
.A(n_5886),
.Y(n_6199)
);

INVx2_ASAP7_75t_L g6200 ( 
.A(n_5891),
.Y(n_6200)
);

NOR2x1_ASAP7_75t_SL g6201 ( 
.A(n_6000),
.B(n_193),
.Y(n_6201)
);

INVx2_ASAP7_75t_L g6202 ( 
.A(n_5891),
.Y(n_6202)
);

NAND2xp5_ASAP7_75t_L g6203 ( 
.A(n_5920),
.B(n_195),
.Y(n_6203)
);

OAI22xp5_ASAP7_75t_L g6204 ( 
.A1(n_5899),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_6204)
);

AOI211xp5_ASAP7_75t_L g6205 ( 
.A1(n_5934),
.A2(n_6027),
.B(n_5926),
.C(n_5925),
.Y(n_6205)
);

OAI22xp33_ASAP7_75t_L g6206 ( 
.A1(n_5894),
.A2(n_6025),
.B1(n_5885),
.B2(n_5889),
.Y(n_6206)
);

OAI21xp33_ASAP7_75t_SL g6207 ( 
.A1(n_5780),
.A2(n_200),
.B(n_201),
.Y(n_6207)
);

BUFx3_ASAP7_75t_L g6208 ( 
.A(n_5821),
.Y(n_6208)
);

NAND2xp5_ASAP7_75t_L g6209 ( 
.A(n_5747),
.B(n_200),
.Y(n_6209)
);

OAI21x1_ASAP7_75t_L g6210 ( 
.A1(n_5780),
.A2(n_2587),
.B(n_2430),
.Y(n_6210)
);

OAI22xp5_ASAP7_75t_L g6211 ( 
.A1(n_5779),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_6211)
);

AOI22xp33_ASAP7_75t_SL g6212 ( 
.A1(n_5932),
.A2(n_5765),
.B1(n_5864),
.B2(n_5792),
.Y(n_6212)
);

OR2x6_ASAP7_75t_L g6213 ( 
.A(n_5934),
.B(n_2111),
.Y(n_6213)
);

HB1xp67_ASAP7_75t_L g6214 ( 
.A(n_5967),
.Y(n_6214)
);

OAI22xp33_ASAP7_75t_L g6215 ( 
.A1(n_5884),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_6215)
);

AND2x2_ASAP7_75t_L g6216 ( 
.A(n_5879),
.B(n_204),
.Y(n_6216)
);

OAI22xp5_ASAP7_75t_L g6217 ( 
.A1(n_5893),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_6217)
);

INVx3_ASAP7_75t_L g6218 ( 
.A(n_5781),
.Y(n_6218)
);

OAI22xp33_ASAP7_75t_L g6219 ( 
.A1(n_6028),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_6219)
);

HB1xp67_ASAP7_75t_L g6220 ( 
.A(n_5801),
.Y(n_6220)
);

NAND3xp33_ASAP7_75t_L g6221 ( 
.A(n_5765),
.B(n_208),
.C(n_209),
.Y(n_6221)
);

AND2x2_ASAP7_75t_L g6222 ( 
.A(n_5879),
.B(n_208),
.Y(n_6222)
);

INVx4_ASAP7_75t_SL g6223 ( 
.A(n_5989),
.Y(n_6223)
);

AOI22xp33_ASAP7_75t_L g6224 ( 
.A1(n_5962),
.A2(n_2122),
.B1(n_2124),
.B2(n_2111),
.Y(n_6224)
);

AOI22xp33_ASAP7_75t_L g6225 ( 
.A1(n_5970),
.A2(n_2124),
.B1(n_2135),
.B2(n_2122),
.Y(n_6225)
);

AND2x4_ASAP7_75t_L g6226 ( 
.A(n_5957),
.B(n_209),
.Y(n_6226)
);

OAI22xp5_ASAP7_75t_L g6227 ( 
.A1(n_5893),
.A2(n_5821),
.B1(n_5879),
.B2(n_5950),
.Y(n_6227)
);

OAI22xp5_ASAP7_75t_L g6228 ( 
.A1(n_5919),
.A2(n_213),
.B1(n_210),
.B2(n_211),
.Y(n_6228)
);

AOI21xp5_ASAP7_75t_L g6229 ( 
.A1(n_5872),
.A2(n_210),
.B(n_211),
.Y(n_6229)
);

OAI222xp33_ASAP7_75t_L g6230 ( 
.A1(n_5833),
.A2(n_216),
.B1(n_221),
.B2(n_213),
.C1(n_214),
.C2(n_218),
.Y(n_6230)
);

BUFx8_ASAP7_75t_SL g6231 ( 
.A(n_6002),
.Y(n_6231)
);

BUFx2_ASAP7_75t_L g6232 ( 
.A(n_5936),
.Y(n_6232)
);

INVx2_ASAP7_75t_L g6233 ( 
.A(n_5892),
.Y(n_6233)
);

OR2x2_ASAP7_75t_L g6234 ( 
.A(n_5749),
.B(n_214),
.Y(n_6234)
);

OAI221xp5_ASAP7_75t_L g6235 ( 
.A1(n_5801),
.A2(n_2433),
.B1(n_2434),
.B2(n_2432),
.C(n_2422),
.Y(n_6235)
);

INVx2_ASAP7_75t_L g6236 ( 
.A(n_5892),
.Y(n_6236)
);

AOI221xp5_ASAP7_75t_L g6237 ( 
.A1(n_5802),
.A2(n_5823),
.B1(n_5937),
.B2(n_5938),
.C(n_5929),
.Y(n_6237)
);

OAI221xp5_ASAP7_75t_L g6238 ( 
.A1(n_5802),
.A2(n_2435),
.B1(n_2436),
.B2(n_2434),
.C(n_2433),
.Y(n_6238)
);

CKINVDCx9p33_ASAP7_75t_R g6239 ( 
.A(n_5971),
.Y(n_6239)
);

OAI22xp5_ASAP7_75t_L g6240 ( 
.A1(n_5870),
.A2(n_222),
.B1(n_216),
.B2(n_218),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_5838),
.Y(n_6241)
);

INVx2_ASAP7_75t_L g6242 ( 
.A(n_5900),
.Y(n_6242)
);

OR2x2_ASAP7_75t_L g6243 ( 
.A(n_5788),
.B(n_5793),
.Y(n_6243)
);

OAI221xp5_ASAP7_75t_L g6244 ( 
.A1(n_5958),
.A2(n_2437),
.B1(n_2439),
.B2(n_2436),
.C(n_2435),
.Y(n_6244)
);

AOI22xp33_ASAP7_75t_L g6245 ( 
.A1(n_5970),
.A2(n_2124),
.B1(n_2135),
.B2(n_2122),
.Y(n_6245)
);

OAI22xp5_ASAP7_75t_L g6246 ( 
.A1(n_6028),
.A2(n_225),
.B1(n_222),
.B2(n_223),
.Y(n_6246)
);

AOI22xp33_ASAP7_75t_L g6247 ( 
.A1(n_5970),
.A2(n_2135),
.B1(n_2142),
.B2(n_2124),
.Y(n_6247)
);

BUFx6f_ASAP7_75t_L g6248 ( 
.A(n_5774),
.Y(n_6248)
);

OAI22xp33_ASAP7_75t_L g6249 ( 
.A1(n_5932),
.A2(n_228),
.B1(n_223),
.B2(n_225),
.Y(n_6249)
);

AOI22xp33_ASAP7_75t_L g6250 ( 
.A1(n_5947),
.A2(n_2142),
.B1(n_2159),
.B2(n_2135),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_5839),
.Y(n_6251)
);

OAI22xp5_ASAP7_75t_L g6252 ( 
.A1(n_6010),
.A2(n_232),
.B1(n_228),
.B2(n_231),
.Y(n_6252)
);

AOI22xp5_ASAP7_75t_L g6253 ( 
.A1(n_5947),
.A2(n_2439),
.B1(n_2440),
.B2(n_2437),
.Y(n_6253)
);

AOI22xp33_ASAP7_75t_L g6254 ( 
.A1(n_5982),
.A2(n_2142),
.B1(n_2159),
.B2(n_2135),
.Y(n_6254)
);

OAI22xp5_ASAP7_75t_L g6255 ( 
.A1(n_6011),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5841),
.Y(n_6256)
);

NOR2xp33_ASAP7_75t_L g6257 ( 
.A(n_5989),
.B(n_234),
.Y(n_6257)
);

HB1xp67_ASAP7_75t_L g6258 ( 
.A(n_5845),
.Y(n_6258)
);

AOI221xp5_ASAP7_75t_SL g6259 ( 
.A1(n_5848),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.C(n_238),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_L g6260 ( 
.A(n_5795),
.B(n_236),
.Y(n_6260)
);

OAI211xp5_ASAP7_75t_L g6261 ( 
.A1(n_5870),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_6261)
);

AOI221xp5_ASAP7_75t_L g6262 ( 
.A1(n_5850),
.A2(n_243),
.B1(n_240),
.B2(n_241),
.C(n_244),
.Y(n_6262)
);

AOI22xp33_ASAP7_75t_L g6263 ( 
.A1(n_5982),
.A2(n_2159),
.B1(n_2174),
.B2(n_2142),
.Y(n_6263)
);

INVx3_ASAP7_75t_L g6264 ( 
.A(n_5781),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5851),
.Y(n_6265)
);

AOI221x1_ASAP7_75t_SL g6266 ( 
.A1(n_5852),
.A2(n_246),
.B1(n_243),
.B2(n_245),
.C(n_247),
.Y(n_6266)
);

INVx2_ASAP7_75t_SL g6267 ( 
.A(n_5805),
.Y(n_6267)
);

INVx2_ASAP7_75t_SL g6268 ( 
.A(n_5805),
.Y(n_6268)
);

AND2x2_ASAP7_75t_L g6269 ( 
.A(n_5995),
.B(n_248),
.Y(n_6269)
);

OAI221xp5_ASAP7_75t_SL g6270 ( 
.A1(n_5861),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.C(n_252),
.Y(n_6270)
);

AND2x2_ASAP7_75t_L g6271 ( 
.A(n_5979),
.B(n_251),
.Y(n_6271)
);

OAI22xp5_ASAP7_75t_L g6272 ( 
.A1(n_5871),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_6272)
);

AOI22xp5_ASAP7_75t_L g6273 ( 
.A1(n_5864),
.A2(n_2445),
.B1(n_2449),
.B2(n_2440),
.Y(n_6273)
);

OAI21x1_ASAP7_75t_L g6274 ( 
.A1(n_5979),
.A2(n_2449),
.B(n_2445),
.Y(n_6274)
);

AOI222xp33_ASAP7_75t_L g6275 ( 
.A1(n_5774),
.A2(n_257),
.B1(n_259),
.B2(n_254),
.C1(n_256),
.C2(n_258),
.Y(n_6275)
);

AOI22xp33_ASAP7_75t_SL g6276 ( 
.A1(n_5765),
.A2(n_262),
.B1(n_256),
.B2(n_260),
.Y(n_6276)
);

AOI22xp33_ASAP7_75t_SL g6277 ( 
.A1(n_5792),
.A2(n_5878),
.B1(n_5872),
.B2(n_5783),
.Y(n_6277)
);

OAI221xp5_ASAP7_75t_L g6278 ( 
.A1(n_5958),
.A2(n_5810),
.B1(n_5807),
.B2(n_5804),
.C(n_5930),
.Y(n_6278)
);

OAI21xp33_ASAP7_75t_SL g6279 ( 
.A1(n_5945),
.A2(n_260),
.B(n_263),
.Y(n_6279)
);

AOI221xp5_ASAP7_75t_L g6280 ( 
.A1(n_5796),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_266),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_5804),
.Y(n_6281)
);

INVx3_ASAP7_75t_L g6282 ( 
.A(n_6188),
.Y(n_6282)
);

AND2x2_ASAP7_75t_L g6283 ( 
.A(n_6141),
.B(n_5974),
.Y(n_6283)
);

BUFx2_ASAP7_75t_L g6284 ( 
.A(n_6239),
.Y(n_6284)
);

INVx2_ASAP7_75t_SL g6285 ( 
.A(n_6063),
.Y(n_6285)
);

OR2x2_ASAP7_75t_L g6286 ( 
.A(n_6189),
.B(n_5956),
.Y(n_6286)
);

AND2x2_ASAP7_75t_L g6287 ( 
.A(n_6083),
.B(n_6188),
.Y(n_6287)
);

INVx2_ASAP7_75t_L g6288 ( 
.A(n_6044),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_6258),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_6044),
.Y(n_6290)
);

OR2x2_ASAP7_75t_L g6291 ( 
.A(n_6052),
.B(n_6038),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_6243),
.Y(n_6292)
);

INVx1_ASAP7_75t_L g6293 ( 
.A(n_6123),
.Y(n_6293)
);

AND2x2_ASAP7_75t_L g6294 ( 
.A(n_6226),
.B(n_5974),
.Y(n_6294)
);

INVx1_ASAP7_75t_L g6295 ( 
.A(n_6129),
.Y(n_6295)
);

OR2x2_ASAP7_75t_L g6296 ( 
.A(n_6117),
.B(n_5961),
.Y(n_6296)
);

AOI22xp33_ASAP7_75t_SL g6297 ( 
.A1(n_6078),
.A2(n_6032),
.B1(n_6035),
.B2(n_6114),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_6226),
.B(n_5985),
.Y(n_6298)
);

INVx2_ASAP7_75t_L g6299 ( 
.A(n_6044),
.Y(n_6299)
);

INVx2_ASAP7_75t_SL g6300 ( 
.A(n_6164),
.Y(n_6300)
);

HB1xp67_ASAP7_75t_L g6301 ( 
.A(n_6113),
.Y(n_6301)
);

AND2x2_ASAP7_75t_L g6302 ( 
.A(n_6135),
.B(n_5985),
.Y(n_6302)
);

INVx2_ASAP7_75t_L g6303 ( 
.A(n_6053),
.Y(n_6303)
);

INVxp67_ASAP7_75t_SL g6304 ( 
.A(n_6221),
.Y(n_6304)
);

AOI22xp33_ASAP7_75t_L g6305 ( 
.A1(n_6078),
.A2(n_5783),
.B1(n_5981),
.B2(n_6000),
.Y(n_6305)
);

OR2x6_ASAP7_75t_L g6306 ( 
.A(n_6164),
.B(n_6000),
.Y(n_6306)
);

INVx3_ASAP7_75t_L g6307 ( 
.A(n_6164),
.Y(n_6307)
);

OR2x2_ASAP7_75t_L g6308 ( 
.A(n_6172),
.B(n_5978),
.Y(n_6308)
);

NAND2xp5_ASAP7_75t_L g6309 ( 
.A(n_6066),
.B(n_5872),
.Y(n_6309)
);

NOR2x1_ASAP7_75t_L g6310 ( 
.A(n_6061),
.B(n_5976),
.Y(n_6310)
);

AND2x2_ASAP7_75t_L g6311 ( 
.A(n_6088),
.B(n_5978),
.Y(n_6311)
);

AND2x2_ASAP7_75t_L g6312 ( 
.A(n_6040),
.B(n_5924),
.Y(n_6312)
);

HB1xp67_ASAP7_75t_L g6313 ( 
.A(n_6154),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_6148),
.Y(n_6314)
);

OAI221xp5_ASAP7_75t_L g6315 ( 
.A1(n_6086),
.A2(n_6046),
.B1(n_6185),
.B2(n_6205),
.C(n_6041),
.Y(n_6315)
);

AND2x2_ASAP7_75t_L g6316 ( 
.A(n_6040),
.B(n_5910),
.Y(n_6316)
);

INVx2_ASAP7_75t_L g6317 ( 
.A(n_6030),
.Y(n_6317)
);

NAND2xp5_ASAP7_75t_L g6318 ( 
.A(n_6057),
.B(n_5878),
.Y(n_6318)
);

AND2x4_ASAP7_75t_L g6319 ( 
.A(n_6043),
.B(n_5878),
.Y(n_6319)
);

INVx1_ASAP7_75t_L g6320 ( 
.A(n_6152),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_6166),
.Y(n_6321)
);

AND2x2_ASAP7_75t_L g6322 ( 
.A(n_6071),
.B(n_5910),
.Y(n_6322)
);

INVx2_ASAP7_75t_L g6323 ( 
.A(n_6033),
.Y(n_6323)
);

INVx1_ASAP7_75t_SL g6324 ( 
.A(n_6072),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_6170),
.Y(n_6325)
);

INVx2_ASAP7_75t_L g6326 ( 
.A(n_6092),
.Y(n_6326)
);

OAI22xp5_ASAP7_75t_L g6327 ( 
.A1(n_6084),
.A2(n_5871),
.B1(n_5921),
.B2(n_5867),
.Y(n_6327)
);

AND2x2_ASAP7_75t_L g6328 ( 
.A(n_6071),
.B(n_5910),
.Y(n_6328)
);

BUFx6f_ASAP7_75t_L g6329 ( 
.A(n_6082),
.Y(n_6329)
);

AND2x2_ASAP7_75t_L g6330 ( 
.A(n_6122),
.B(n_6248),
.Y(n_6330)
);

INVx2_ASAP7_75t_L g6331 ( 
.A(n_6045),
.Y(n_6331)
);

OR2x2_ASAP7_75t_L g6332 ( 
.A(n_6214),
.B(n_6014),
.Y(n_6332)
);

A2O1A1Ixp33_ASAP7_75t_L g6333 ( 
.A1(n_6266),
.A2(n_5981),
.B(n_6000),
.C(n_5753),
.Y(n_6333)
);

CKINVDCx6p67_ASAP7_75t_R g6334 ( 
.A(n_6082),
.Y(n_6334)
);

OR2x2_ASAP7_75t_L g6335 ( 
.A(n_6056),
.B(n_6014),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_6178),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_6104),
.Y(n_6337)
);

BUFx2_ASAP7_75t_L g6338 ( 
.A(n_6223),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_6186),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_6187),
.Y(n_6340)
);

INVx2_ASAP7_75t_L g6341 ( 
.A(n_6109),
.Y(n_6341)
);

AND2x2_ASAP7_75t_L g6342 ( 
.A(n_6122),
.B(n_5867),
.Y(n_6342)
);

INVx2_ASAP7_75t_SL g6343 ( 
.A(n_6082),
.Y(n_6343)
);

INVx1_ASAP7_75t_L g6344 ( 
.A(n_6241),
.Y(n_6344)
);

BUFx3_ASAP7_75t_L g6345 ( 
.A(n_6231),
.Y(n_6345)
);

AND2x2_ASAP7_75t_L g6346 ( 
.A(n_6248),
.B(n_5921),
.Y(n_6346)
);

AND2x2_ASAP7_75t_L g6347 ( 
.A(n_6248),
.B(n_5923),
.Y(n_6347)
);

INVx2_ASAP7_75t_L g6348 ( 
.A(n_6116),
.Y(n_6348)
);

NAND2xp5_ASAP7_75t_L g6349 ( 
.A(n_6074),
.B(n_5923),
.Y(n_6349)
);

BUFx6f_ASAP7_75t_L g6350 ( 
.A(n_6127),
.Y(n_6350)
);

INVx1_ASAP7_75t_L g6351 ( 
.A(n_6251),
.Y(n_6351)
);

AND2x2_ASAP7_75t_L g6352 ( 
.A(n_6223),
.B(n_6026),
.Y(n_6352)
);

OR2x2_ASAP7_75t_L g6353 ( 
.A(n_6095),
.B(n_6016),
.Y(n_6353)
);

INVx2_ASAP7_75t_L g6354 ( 
.A(n_6126),
.Y(n_6354)
);

INVx2_ASAP7_75t_L g6355 ( 
.A(n_6151),
.Y(n_6355)
);

INVx2_ASAP7_75t_L g6356 ( 
.A(n_6153),
.Y(n_6356)
);

BUFx6f_ASAP7_75t_L g6357 ( 
.A(n_6181),
.Y(n_6357)
);

INVx2_ASAP7_75t_L g6358 ( 
.A(n_6194),
.Y(n_6358)
);

INVx1_ASAP7_75t_L g6359 ( 
.A(n_6256),
.Y(n_6359)
);

INVx2_ASAP7_75t_L g6360 ( 
.A(n_6199),
.Y(n_6360)
);

BUFx3_ASAP7_75t_L g6361 ( 
.A(n_6232),
.Y(n_6361)
);

INVx1_ASAP7_75t_L g6362 ( 
.A(n_6265),
.Y(n_6362)
);

AND2x2_ASAP7_75t_L g6363 ( 
.A(n_6223),
.B(n_6026),
.Y(n_6363)
);

AND2x2_ASAP7_75t_L g6364 ( 
.A(n_6106),
.B(n_5976),
.Y(n_6364)
);

AND2x2_ASAP7_75t_L g6365 ( 
.A(n_6043),
.B(n_5989),
.Y(n_6365)
);

AND2x2_ASAP7_75t_L g6366 ( 
.A(n_6051),
.B(n_5922),
.Y(n_6366)
);

AND2x2_ASAP7_75t_L g6367 ( 
.A(n_6051),
.B(n_6017),
.Y(n_6367)
);

AND2x2_ASAP7_75t_L g6368 ( 
.A(n_6073),
.B(n_6019),
.Y(n_6368)
);

OR2x2_ASAP7_75t_L g6369 ( 
.A(n_6115),
.B(n_5896),
.Y(n_6369)
);

INVx2_ASAP7_75t_L g6370 ( 
.A(n_6200),
.Y(n_6370)
);

INVx2_ASAP7_75t_L g6371 ( 
.A(n_6202),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_6029),
.Y(n_6372)
);

INVx2_ASAP7_75t_SL g6373 ( 
.A(n_6267),
.Y(n_6373)
);

NOR2xp33_ASAP7_75t_L g6374 ( 
.A(n_6165),
.B(n_5868),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_6055),
.Y(n_6375)
);

NAND2xp5_ASAP7_75t_L g6376 ( 
.A(n_6039),
.B(n_5896),
.Y(n_6376)
);

OAI211xp5_ASAP7_75t_L g6377 ( 
.A1(n_6069),
.A2(n_5988),
.B(n_5811),
.C(n_6003),
.Y(n_6377)
);

HB1xp67_ASAP7_75t_L g6378 ( 
.A(n_6065),
.Y(n_6378)
);

HB1xp67_ASAP7_75t_L g6379 ( 
.A(n_6101),
.Y(n_6379)
);

INVx1_ASAP7_75t_L g6380 ( 
.A(n_6058),
.Y(n_6380)
);

NAND2xp5_ASAP7_75t_L g6381 ( 
.A(n_6110),
.B(n_5896),
.Y(n_6381)
);

AND2x2_ASAP7_75t_L g6382 ( 
.A(n_6216),
.B(n_5943),
.Y(n_6382)
);

INVx2_ASAP7_75t_L g6383 ( 
.A(n_6233),
.Y(n_6383)
);

INVx2_ASAP7_75t_L g6384 ( 
.A(n_6236),
.Y(n_6384)
);

AND2x4_ASAP7_75t_L g6385 ( 
.A(n_6085),
.B(n_5943),
.Y(n_6385)
);

AND2x2_ASAP7_75t_L g6386 ( 
.A(n_6222),
.B(n_5943),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_6140),
.Y(n_6387)
);

AND2x2_ASAP7_75t_L g6388 ( 
.A(n_6205),
.B(n_5917),
.Y(n_6388)
);

INVx2_ASAP7_75t_L g6389 ( 
.A(n_6242),
.Y(n_6389)
);

BUFx3_ASAP7_75t_L g6390 ( 
.A(n_6208),
.Y(n_6390)
);

NAND2xp5_ASAP7_75t_L g6391 ( 
.A(n_6110),
.B(n_5959),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6145),
.Y(n_6392)
);

HB1xp67_ASAP7_75t_L g6393 ( 
.A(n_6221),
.Y(n_6393)
);

CKINVDCx14_ASAP7_75t_R g6394 ( 
.A(n_6070),
.Y(n_6394)
);

INVx2_ASAP7_75t_L g6395 ( 
.A(n_6281),
.Y(n_6395)
);

INVxp67_ASAP7_75t_L g6396 ( 
.A(n_6167),
.Y(n_6396)
);

INVxp67_ASAP7_75t_L g6397 ( 
.A(n_6128),
.Y(n_6397)
);

BUFx2_ASAP7_75t_L g6398 ( 
.A(n_6268),
.Y(n_6398)
);

OR2x2_ASAP7_75t_L g6399 ( 
.A(n_6080),
.B(n_6003),
.Y(n_6399)
);

NAND2x1_ASAP7_75t_L g6400 ( 
.A(n_6218),
.B(n_6264),
.Y(n_6400)
);

AND2x2_ASAP7_75t_L g6401 ( 
.A(n_6085),
.B(n_6006),
.Y(n_6401)
);

BUFx3_ASAP7_75t_L g6402 ( 
.A(n_6093),
.Y(n_6402)
);

OR2x2_ASAP7_75t_L g6403 ( 
.A(n_6203),
.B(n_6006),
.Y(n_6403)
);

INVx2_ASAP7_75t_L g6404 ( 
.A(n_6220),
.Y(n_6404)
);

NAND2xp5_ASAP7_75t_L g6405 ( 
.A(n_6067),
.B(n_5959),
.Y(n_6405)
);

OR2x2_ASAP7_75t_L g6406 ( 
.A(n_6234),
.B(n_5811),
.Y(n_6406)
);

NAND2xp5_ASAP7_75t_L g6407 ( 
.A(n_6198),
.B(n_5807),
.Y(n_6407)
);

INVx2_ASAP7_75t_L g6408 ( 
.A(n_6064),
.Y(n_6408)
);

INVx2_ASAP7_75t_L g6409 ( 
.A(n_6177),
.Y(n_6409)
);

BUFx2_ASAP7_75t_L g6410 ( 
.A(n_6207),
.Y(n_6410)
);

AND2x2_ASAP7_75t_L g6411 ( 
.A(n_6227),
.B(n_5777),
.Y(n_6411)
);

HB1xp67_ASAP7_75t_L g6412 ( 
.A(n_6260),
.Y(n_6412)
);

OAI21xp5_ASAP7_75t_L g6413 ( 
.A1(n_6146),
.A2(n_5965),
.B(n_5819),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_6209),
.Y(n_6414)
);

OR2x2_ASAP7_75t_L g6415 ( 
.A(n_6161),
.B(n_5930),
.Y(n_6415)
);

AOI22xp33_ASAP7_75t_L g6416 ( 
.A1(n_6034),
.A2(n_5927),
.B1(n_5992),
.B2(n_5993),
.Y(n_6416)
);

INVx2_ASAP7_75t_L g6417 ( 
.A(n_6177),
.Y(n_6417)
);

INVx2_ASAP7_75t_L g6418 ( 
.A(n_6213),
.Y(n_6418)
);

NOR2xp33_ASAP7_75t_L g6419 ( 
.A(n_6054),
.B(n_6002),
.Y(n_6419)
);

OR2x2_ASAP7_75t_L g6420 ( 
.A(n_6090),
.B(n_5933),
.Y(n_6420)
);

AND2x2_ASAP7_75t_L g6421 ( 
.A(n_6144),
.B(n_5777),
.Y(n_6421)
);

HB1xp67_ASAP7_75t_L g6422 ( 
.A(n_6237),
.Y(n_6422)
);

AND2x4_ASAP7_75t_L g6423 ( 
.A(n_6037),
.B(n_5965),
.Y(n_6423)
);

HB1xp67_ASAP7_75t_L g6424 ( 
.A(n_6213),
.Y(n_6424)
);

AND2x2_ASAP7_75t_L g6425 ( 
.A(n_6144),
.B(n_5980),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6271),
.Y(n_6426)
);

AND2x2_ASAP7_75t_L g6427 ( 
.A(n_6144),
.B(n_5980),
.Y(n_6427)
);

OR2x2_ASAP7_75t_L g6428 ( 
.A(n_6138),
.B(n_5933),
.Y(n_6428)
);

BUFx2_ASAP7_75t_L g6429 ( 
.A(n_6279),
.Y(n_6429)
);

AND2x2_ASAP7_75t_L g6430 ( 
.A(n_6218),
.B(n_5819),
.Y(n_6430)
);

AOI22xp33_ASAP7_75t_L g6431 ( 
.A1(n_6035),
.A2(n_5927),
.B1(n_5992),
.B2(n_5993),
.Y(n_6431)
);

INVx2_ASAP7_75t_L g6432 ( 
.A(n_6213),
.Y(n_6432)
);

AND2x2_ASAP7_75t_L g6433 ( 
.A(n_6264),
.B(n_6147),
.Y(n_6433)
);

HB1xp67_ASAP7_75t_L g6434 ( 
.A(n_6168),
.Y(n_6434)
);

INVx2_ASAP7_75t_L g6435 ( 
.A(n_6111),
.Y(n_6435)
);

INVx2_ASAP7_75t_L g6436 ( 
.A(n_6278),
.Y(n_6436)
);

AND2x2_ASAP7_75t_L g6437 ( 
.A(n_6156),
.B(n_5828),
.Y(n_6437)
);

INVx2_ASAP7_75t_L g6438 ( 
.A(n_6149),
.Y(n_6438)
);

INVx2_ASAP7_75t_L g6439 ( 
.A(n_6158),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_6182),
.Y(n_6440)
);

NAND2x1p5_ASAP7_75t_L g6441 ( 
.A(n_6077),
.B(n_5927),
.Y(n_6441)
);

OR2x2_ASAP7_75t_L g6442 ( 
.A(n_6059),
.B(n_5941),
.Y(n_6442)
);

INVx2_ASAP7_75t_L g6443 ( 
.A(n_6139),
.Y(n_6443)
);

AND2x2_ASAP7_75t_L g6444 ( 
.A(n_6191),
.B(n_5828),
.Y(n_6444)
);

INVx2_ASAP7_75t_L g6445 ( 
.A(n_6139),
.Y(n_6445)
);

NAND3xp33_ASAP7_75t_L g6446 ( 
.A(n_6171),
.B(n_5756),
.C(n_6013),
.Y(n_6446)
);

AND2x2_ASAP7_75t_L g6447 ( 
.A(n_6062),
.B(n_5756),
.Y(n_6447)
);

AND2x2_ASAP7_75t_L g6448 ( 
.A(n_6047),
.B(n_5756),
.Y(n_6448)
);

HB1xp67_ASAP7_75t_L g6449 ( 
.A(n_6273),
.Y(n_6449)
);

NAND2xp5_ASAP7_75t_L g6450 ( 
.A(n_6036),
.B(n_5810),
.Y(n_6450)
);

INVx1_ASAP7_75t_L g6451 ( 
.A(n_6253),
.Y(n_6451)
);

AOI22xp33_ASAP7_75t_L g6452 ( 
.A1(n_6050),
.A2(n_6013),
.B1(n_5941),
.B2(n_5982),
.Y(n_6452)
);

INVx2_ASAP7_75t_L g6453 ( 
.A(n_6139),
.Y(n_6453)
);

INVx2_ASAP7_75t_L g6454 ( 
.A(n_6269),
.Y(n_6454)
);

CKINVDCx14_ASAP7_75t_R g6455 ( 
.A(n_6240),
.Y(n_6455)
);

HB1xp67_ASAP7_75t_L g6456 ( 
.A(n_6049),
.Y(n_6456)
);

AOI22xp33_ASAP7_75t_L g6457 ( 
.A1(n_6048),
.A2(n_5832),
.B1(n_5844),
.B2(n_5843),
.Y(n_6457)
);

AND2x4_ASAP7_75t_L g6458 ( 
.A(n_6096),
.B(n_5840),
.Y(n_6458)
);

AOI22xp33_ASAP7_75t_L g6459 ( 
.A1(n_6089),
.A2(n_5832),
.B1(n_5844),
.B2(n_5843),
.Y(n_6459)
);

INVx2_ASAP7_75t_L g6460 ( 
.A(n_6157),
.Y(n_6460)
);

INVx1_ASAP7_75t_L g6461 ( 
.A(n_6094),
.Y(n_6461)
);

INVx1_ASAP7_75t_L g6462 ( 
.A(n_6099),
.Y(n_6462)
);

AND2x2_ASAP7_75t_L g6463 ( 
.A(n_6075),
.B(n_5840),
.Y(n_6463)
);

BUFx3_ASAP7_75t_L g6464 ( 
.A(n_6257),
.Y(n_6464)
);

HB1xp67_ASAP7_75t_L g6465 ( 
.A(n_6125),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6249),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_6097),
.Y(n_6467)
);

AND2x2_ASAP7_75t_L g6468 ( 
.A(n_6160),
.B(n_5902),
.Y(n_6468)
);

AND2x2_ASAP7_75t_L g6469 ( 
.A(n_6277),
.B(n_5903),
.Y(n_6469)
);

INVx1_ASAP7_75t_L g6470 ( 
.A(n_6180),
.Y(n_6470)
);

BUFx6f_ASAP7_75t_L g6471 ( 
.A(n_6274),
.Y(n_6471)
);

INVx1_ASAP7_75t_L g6472 ( 
.A(n_6229),
.Y(n_6472)
);

INVx2_ASAP7_75t_L g6473 ( 
.A(n_6201),
.Y(n_6473)
);

OR2x2_ASAP7_75t_L g6474 ( 
.A(n_6068),
.B(n_5904),
.Y(n_6474)
);

AND2x2_ASAP7_75t_L g6475 ( 
.A(n_6179),
.B(n_5905),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_6134),
.Y(n_6476)
);

INVx2_ASAP7_75t_L g6477 ( 
.A(n_6176),
.Y(n_6477)
);

INVx1_ASAP7_75t_L g6478 ( 
.A(n_6134),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_6235),
.Y(n_6479)
);

INVxp67_ASAP7_75t_SL g6480 ( 
.A(n_6212),
.Y(n_6480)
);

AND2x4_ASAP7_75t_L g6481 ( 
.A(n_6076),
.B(n_5808),
.Y(n_6481)
);

AND2x4_ASAP7_75t_L g6482 ( 
.A(n_6079),
.B(n_5808),
.Y(n_6482)
);

NAND2xp5_ASAP7_75t_L g6483 ( 
.A(n_6276),
.B(n_5907),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_6238),
.Y(n_6484)
);

OR2x2_ASAP7_75t_L g6485 ( 
.A(n_6042),
.B(n_5912),
.Y(n_6485)
);

INVx2_ASAP7_75t_L g6486 ( 
.A(n_6210),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6204),
.Y(n_6487)
);

AND2x4_ASAP7_75t_L g6488 ( 
.A(n_6081),
.B(n_5969),
.Y(n_6488)
);

AND2x2_ASAP7_75t_L g6489 ( 
.A(n_6060),
.B(n_5914),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_6204),
.Y(n_6490)
);

AND2x2_ASAP7_75t_L g6491 ( 
.A(n_6131),
.B(n_5900),
.Y(n_6491)
);

INVx2_ASAP7_75t_L g6492 ( 
.A(n_6130),
.Y(n_6492)
);

AOI22xp33_ASAP7_75t_L g6493 ( 
.A1(n_6087),
.A2(n_5854),
.B1(n_5764),
.B2(n_5759),
.Y(n_6493)
);

HB1xp67_ASAP7_75t_L g6494 ( 
.A(n_6266),
.Y(n_6494)
);

INVx2_ASAP7_75t_L g6495 ( 
.A(n_6240),
.Y(n_6495)
);

AND2x2_ASAP7_75t_L g6496 ( 
.A(n_6259),
.B(n_5901),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_6244),
.Y(n_6497)
);

AND2x2_ASAP7_75t_L g6498 ( 
.A(n_6259),
.B(n_5901),
.Y(n_6498)
);

INVx1_ASAP7_75t_L g6499 ( 
.A(n_6108),
.Y(n_6499)
);

INVx2_ASAP7_75t_L g6500 ( 
.A(n_6217),
.Y(n_6500)
);

INVx2_ASAP7_75t_L g6501 ( 
.A(n_6246),
.Y(n_6501)
);

INVx2_ASAP7_75t_L g6502 ( 
.A(n_6211),
.Y(n_6502)
);

INVx2_ASAP7_75t_SL g6503 ( 
.A(n_6211),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6206),
.Y(n_6504)
);

INVx2_ASAP7_75t_L g6505 ( 
.A(n_6252),
.Y(n_6505)
);

NAND2xp5_ASAP7_75t_L g6506 ( 
.A(n_6142),
.B(n_6133),
.Y(n_6506)
);

INVx1_ASAP7_75t_L g6507 ( 
.A(n_6098),
.Y(n_6507)
);

AND2x2_ASAP7_75t_L g6508 ( 
.A(n_6124),
.B(n_5906),
.Y(n_6508)
);

INVx2_ASAP7_75t_L g6509 ( 
.A(n_6255),
.Y(n_6509)
);

INVx1_ASAP7_75t_SL g6510 ( 
.A(n_6162),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6100),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_6174),
.Y(n_6512)
);

INVx2_ASAP7_75t_L g6513 ( 
.A(n_6175),
.Y(n_6513)
);

AND2x2_ASAP7_75t_L g6514 ( 
.A(n_6031),
.B(n_5906),
.Y(n_6514)
);

AND2x2_ASAP7_75t_L g6515 ( 
.A(n_6250),
.B(n_5913),
.Y(n_6515)
);

INVx1_ASAP7_75t_L g6516 ( 
.A(n_6215),
.Y(n_6516)
);

INVx3_ASAP7_75t_L g6517 ( 
.A(n_6137),
.Y(n_6517)
);

AOI22xp33_ASAP7_75t_L g6518 ( 
.A1(n_6192),
.A2(n_5854),
.B1(n_5764),
.B2(n_5759),
.Y(n_6518)
);

AND2x2_ASAP7_75t_L g6519 ( 
.A(n_6196),
.B(n_5913),
.Y(n_6519)
);

HB1xp67_ASAP7_75t_L g6520 ( 
.A(n_6197),
.Y(n_6520)
);

BUFx6f_ASAP7_75t_L g6521 ( 
.A(n_6275),
.Y(n_6521)
);

HB1xp67_ASAP7_75t_L g6522 ( 
.A(n_6169),
.Y(n_6522)
);

INVx2_ASAP7_75t_L g6523 ( 
.A(n_6107),
.Y(n_6523)
);

OR2x2_ASAP7_75t_L g6524 ( 
.A(n_6150),
.B(n_5915),
.Y(n_6524)
);

BUFx3_ASAP7_75t_L g6525 ( 
.A(n_6228),
.Y(n_6525)
);

BUFx3_ASAP7_75t_L g6526 ( 
.A(n_6272),
.Y(n_6526)
);

AND2x2_ASAP7_75t_L g6527 ( 
.A(n_6284),
.B(n_6121),
.Y(n_6527)
);

AOI22xp5_ASAP7_75t_L g6528 ( 
.A1(n_6521),
.A2(n_6261),
.B1(n_6195),
.B2(n_6275),
.Y(n_6528)
);

INVx1_ASAP7_75t_L g6529 ( 
.A(n_6293),
.Y(n_6529)
);

OAI21xp5_ASAP7_75t_L g6530 ( 
.A1(n_6297),
.A2(n_6230),
.B(n_6173),
.Y(n_6530)
);

INVx1_ASAP7_75t_L g6531 ( 
.A(n_6295),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_6314),
.Y(n_6532)
);

AOI322xp5_ASAP7_75t_L g6533 ( 
.A1(n_6494),
.A2(n_6280),
.A3(n_6262),
.B1(n_6219),
.B2(n_6103),
.C1(n_6091),
.C2(n_6102),
.Y(n_6533)
);

AO21x2_ASAP7_75t_L g6534 ( 
.A1(n_6480),
.A2(n_6190),
.B(n_6105),
.Y(n_6534)
);

OAI211xp5_ASAP7_75t_L g6535 ( 
.A1(n_6297),
.A2(n_6195),
.B(n_6193),
.C(n_6270),
.Y(n_6535)
);

AOI22xp33_ASAP7_75t_L g6536 ( 
.A1(n_6521),
.A2(n_6118),
.B1(n_6132),
.B2(n_6136),
.Y(n_6536)
);

OAI221xp5_ASAP7_75t_L g6537 ( 
.A1(n_6480),
.A2(n_6193),
.B1(n_6120),
.B2(n_6119),
.C(n_6225),
.Y(n_6537)
);

AOI31xp33_ASAP7_75t_L g6538 ( 
.A1(n_6494),
.A2(n_6456),
.A3(n_6304),
.B(n_6394),
.Y(n_6538)
);

INVx2_ASAP7_75t_L g6539 ( 
.A(n_6390),
.Y(n_6539)
);

OAI221xp5_ASAP7_75t_L g6540 ( 
.A1(n_6521),
.A2(n_6120),
.B1(n_6247),
.B2(n_6245),
.C(n_6254),
.Y(n_6540)
);

OA222x2_ASAP7_75t_L g6541 ( 
.A1(n_6381),
.A2(n_5969),
.B1(n_5983),
.B2(n_5977),
.C1(n_5754),
.C2(n_5757),
.Y(n_6541)
);

NAND4xp25_ASAP7_75t_L g6542 ( 
.A(n_6419),
.B(n_6224),
.C(n_6112),
.D(n_6184),
.Y(n_6542)
);

NAND3xp33_ASAP7_75t_L g6543 ( 
.A(n_6521),
.B(n_6159),
.C(n_6155),
.Y(n_6543)
);

AOI22xp33_ASAP7_75t_L g6544 ( 
.A1(n_6435),
.A2(n_6263),
.B1(n_6183),
.B2(n_6143),
.Y(n_6544)
);

AOI21xp33_ASAP7_75t_SL g6545 ( 
.A1(n_6419),
.A2(n_265),
.B(n_267),
.Y(n_6545)
);

OAI211xp5_ASAP7_75t_L g6546 ( 
.A1(n_6377),
.A2(n_6163),
.B(n_5977),
.C(n_5983),
.Y(n_6546)
);

INVx2_ASAP7_75t_L g6547 ( 
.A(n_6390),
.Y(n_6547)
);

OA21x2_ASAP7_75t_L g6548 ( 
.A1(n_6391),
.A2(n_5754),
.B(n_5748),
.Y(n_6548)
);

OAI211xp5_ASAP7_75t_L g6549 ( 
.A1(n_6456),
.A2(n_5946),
.B(n_5757),
.C(n_5748),
.Y(n_6549)
);

OAI221xp5_ASAP7_75t_L g6550 ( 
.A1(n_6304),
.A2(n_6315),
.B1(n_6416),
.B2(n_6431),
.C(n_6429),
.Y(n_6550)
);

INVx1_ASAP7_75t_L g6551 ( 
.A(n_6320),
.Y(n_6551)
);

INVx2_ASAP7_75t_L g6552 ( 
.A(n_6471),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_6321),
.Y(n_6553)
);

AOI33xp33_ASAP7_75t_L g6554 ( 
.A1(n_6462),
.A2(n_5946),
.A3(n_5767),
.B1(n_5768),
.B2(n_5766),
.B3(n_273),
.Y(n_6554)
);

NAND3xp33_ASAP7_75t_SL g6555 ( 
.A(n_6410),
.B(n_5767),
.C(n_5766),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_6325),
.Y(n_6556)
);

OAI22xp5_ASAP7_75t_L g6557 ( 
.A1(n_6455),
.A2(n_5768),
.B1(n_5915),
.B2(n_274),
.Y(n_6557)
);

OR2x2_ASAP7_75t_L g6558 ( 
.A(n_6291),
.B(n_270),
.Y(n_6558)
);

OAI322xp33_ASAP7_75t_L g6559 ( 
.A1(n_6455),
.A2(n_278),
.A3(n_277),
.B1(n_274),
.B2(n_270),
.C1(n_271),
.C2(n_276),
.Y(n_6559)
);

AOI33xp33_ASAP7_75t_L g6560 ( 
.A1(n_6467),
.A2(n_279),
.A3(n_282),
.B1(n_276),
.B2(n_278),
.B3(n_280),
.Y(n_6560)
);

INVx2_ASAP7_75t_L g6561 ( 
.A(n_6471),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_6336),
.Y(n_6562)
);

AOI321xp33_ASAP7_75t_L g6563 ( 
.A1(n_6495),
.A2(n_285),
.A3(n_288),
.B1(n_280),
.B2(n_283),
.C(n_287),
.Y(n_6563)
);

INVx1_ASAP7_75t_L g6564 ( 
.A(n_6339),
.Y(n_6564)
);

OR2x2_ASAP7_75t_L g6565 ( 
.A(n_6476),
.B(n_283),
.Y(n_6565)
);

OAI21xp5_ASAP7_75t_L g6566 ( 
.A1(n_6393),
.A2(n_6333),
.B(n_6422),
.Y(n_6566)
);

NAND2xp5_ASAP7_75t_L g6567 ( 
.A(n_6393),
.B(n_6496),
.Y(n_6567)
);

AOI21xp5_ASAP7_75t_L g6568 ( 
.A1(n_6422),
.A2(n_285),
.B(n_288),
.Y(n_6568)
);

BUFx2_ASAP7_75t_L g6569 ( 
.A(n_6421),
.Y(n_6569)
);

HB1xp67_ASAP7_75t_L g6570 ( 
.A(n_6361),
.Y(n_6570)
);

INVx1_ASAP7_75t_L g6571 ( 
.A(n_6340),
.Y(n_6571)
);

AOI22xp33_ASAP7_75t_L g6572 ( 
.A1(n_6435),
.A2(n_2468),
.B1(n_2473),
.B2(n_2455),
.Y(n_6572)
);

HB1xp67_ASAP7_75t_L g6573 ( 
.A(n_6361),
.Y(n_6573)
);

INVx2_ASAP7_75t_L g6574 ( 
.A(n_6471),
.Y(n_6574)
);

NOR2xp33_ASAP7_75t_L g6575 ( 
.A(n_6345),
.B(n_289),
.Y(n_6575)
);

AND2x2_ASAP7_75t_L g6576 ( 
.A(n_6310),
.B(n_289),
.Y(n_6576)
);

AND2x2_ASAP7_75t_L g6577 ( 
.A(n_6433),
.B(n_291),
.Y(n_6577)
);

OAI22xp5_ASAP7_75t_L g6578 ( 
.A1(n_6327),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_6344),
.Y(n_6579)
);

INVx1_ASAP7_75t_L g6580 ( 
.A(n_6351),
.Y(n_6580)
);

OR2x2_ASAP7_75t_L g6581 ( 
.A(n_6478),
.B(n_292),
.Y(n_6581)
);

OAI22xp33_ASAP7_75t_L g6582 ( 
.A1(n_6376),
.A2(n_296),
.B1(n_293),
.B2(n_295),
.Y(n_6582)
);

AO21x2_ASAP7_75t_L g6583 ( 
.A1(n_6512),
.A2(n_2468),
.B(n_2455),
.Y(n_6583)
);

OAI221xp5_ASAP7_75t_SL g6584 ( 
.A1(n_6333),
.A2(n_298),
.B1(n_295),
.B2(n_297),
.C(n_300),
.Y(n_6584)
);

OR2x2_ASAP7_75t_L g6585 ( 
.A(n_6292),
.B(n_297),
.Y(n_6585)
);

AND2x4_ASAP7_75t_L g6586 ( 
.A(n_6365),
.B(n_301),
.Y(n_6586)
);

AOI221xp5_ASAP7_75t_L g6587 ( 
.A1(n_6416),
.A2(n_309),
.B1(n_304),
.B2(n_307),
.C(n_310),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6359),
.Y(n_6588)
);

AOI22xp33_ASAP7_75t_L g6589 ( 
.A1(n_6523),
.A2(n_2476),
.B1(n_2479),
.B2(n_2473),
.Y(n_6589)
);

AOI22xp33_ASAP7_75t_L g6590 ( 
.A1(n_6523),
.A2(n_2479),
.B1(n_2476),
.B2(n_2159),
.Y(n_6590)
);

OR2x2_ASAP7_75t_L g6591 ( 
.A(n_6487),
.B(n_307),
.Y(n_6591)
);

OAI221xp5_ASAP7_75t_L g6592 ( 
.A1(n_6431),
.A2(n_313),
.B1(n_310),
.B2(n_312),
.C(n_314),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6362),
.Y(n_6593)
);

NAND2xp5_ASAP7_75t_L g6594 ( 
.A(n_6498),
.B(n_312),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_6301),
.Y(n_6595)
);

INVx1_ASAP7_75t_L g6596 ( 
.A(n_6301),
.Y(n_6596)
);

AOI221xp5_ASAP7_75t_L g6597 ( 
.A1(n_6396),
.A2(n_316),
.B1(n_313),
.B2(n_314),
.C(n_317),
.Y(n_6597)
);

INVx2_ASAP7_75t_L g6598 ( 
.A(n_6471),
.Y(n_6598)
);

BUFx3_ASAP7_75t_L g6599 ( 
.A(n_6345),
.Y(n_6599)
);

OAI22xp33_ASAP7_75t_L g6600 ( 
.A1(n_6309),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_6600)
);

AOI22xp33_ASAP7_75t_L g6601 ( 
.A1(n_6461),
.A2(n_2159),
.B1(n_2174),
.B2(n_2142),
.Y(n_6601)
);

BUFx2_ASAP7_75t_L g6602 ( 
.A(n_6425),
.Y(n_6602)
);

AND2x2_ASAP7_75t_L g6603 ( 
.A(n_6283),
.B(n_318),
.Y(n_6603)
);

INVx2_ASAP7_75t_L g6604 ( 
.A(n_6454),
.Y(n_6604)
);

NAND2xp5_ASAP7_75t_L g6605 ( 
.A(n_6412),
.B(n_319),
.Y(n_6605)
);

HB1xp67_ASAP7_75t_L g6606 ( 
.A(n_6313),
.Y(n_6606)
);

OAI221xp5_ASAP7_75t_L g6607 ( 
.A1(n_6459),
.A2(n_6305),
.B1(n_6457),
.B2(n_6396),
.C(n_6413),
.Y(n_6607)
);

AOI22xp33_ASAP7_75t_L g6608 ( 
.A1(n_6459),
.A2(n_2174),
.B1(n_2443),
.B2(n_2431),
.Y(n_6608)
);

AOI22xp33_ASAP7_75t_L g6609 ( 
.A1(n_6448),
.A2(n_2174),
.B1(n_2443),
.B2(n_2431),
.Y(n_6609)
);

INVx1_ASAP7_75t_L g6610 ( 
.A(n_6313),
.Y(n_6610)
);

OAI33xp33_ASAP7_75t_L g6611 ( 
.A1(n_6506),
.A2(n_323),
.A3(n_325),
.B1(n_319),
.B2(n_321),
.B3(n_324),
.Y(n_6611)
);

INVx2_ASAP7_75t_L g6612 ( 
.A(n_6454),
.Y(n_6612)
);

INVx2_ASAP7_75t_L g6613 ( 
.A(n_6439),
.Y(n_6613)
);

AOI22xp33_ASAP7_75t_L g6614 ( 
.A1(n_6520),
.A2(n_2174),
.B1(n_2443),
.B2(n_2431),
.Y(n_6614)
);

OR2x2_ASAP7_75t_L g6615 ( 
.A(n_6490),
.B(n_321),
.Y(n_6615)
);

AND2x2_ASAP7_75t_L g6616 ( 
.A(n_6352),
.B(n_323),
.Y(n_6616)
);

OAI22xp5_ASAP7_75t_L g6617 ( 
.A1(n_6394),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_6617)
);

AND2x2_ASAP7_75t_L g6618 ( 
.A(n_6363),
.B(n_326),
.Y(n_6618)
);

AOI221xp5_ASAP7_75t_L g6619 ( 
.A1(n_6482),
.A2(n_331),
.B1(n_328),
.B2(n_329),
.C(n_332),
.Y(n_6619)
);

AOI22xp33_ASAP7_75t_SL g6620 ( 
.A1(n_6463),
.A2(n_333),
.B1(n_329),
.B2(n_331),
.Y(n_6620)
);

INVx2_ASAP7_75t_SL g6621 ( 
.A(n_6350),
.Y(n_6621)
);

OAI22xp33_ASAP7_75t_L g6622 ( 
.A1(n_6407),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_6622)
);

OR2x2_ASAP7_75t_L g6623 ( 
.A(n_6412),
.B(n_335),
.Y(n_6623)
);

AOI22xp33_ASAP7_75t_SL g6624 ( 
.A1(n_6388),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_6624)
);

INVx2_ASAP7_75t_L g6625 ( 
.A(n_6439),
.Y(n_6625)
);

NAND2xp5_ASAP7_75t_L g6626 ( 
.A(n_6465),
.B(n_339),
.Y(n_6626)
);

AOI21xp5_ASAP7_75t_L g6627 ( 
.A1(n_6520),
.A2(n_339),
.B(n_340),
.Y(n_6627)
);

AOI22xp5_ASAP7_75t_L g6628 ( 
.A1(n_6472),
.A2(n_344),
.B1(n_340),
.B2(n_342),
.Y(n_6628)
);

AND2x2_ASAP7_75t_L g6629 ( 
.A(n_6330),
.B(n_6306),
.Y(n_6629)
);

OAI21xp5_ASAP7_75t_L g6630 ( 
.A1(n_6305),
.A2(n_345),
.B(n_347),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6306),
.B(n_6316),
.Y(n_6631)
);

AOI21xp5_ASAP7_75t_L g6632 ( 
.A1(n_6465),
.A2(n_345),
.B(n_347),
.Y(n_6632)
);

AND2x2_ASAP7_75t_L g6633 ( 
.A(n_6306),
.B(n_349),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_6289),
.Y(n_6634)
);

AO21x2_ASAP7_75t_L g6635 ( 
.A1(n_6504),
.A2(n_349),
.B(n_350),
.Y(n_6635)
);

OAI22xp33_ASAP7_75t_L g6636 ( 
.A1(n_6442),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_6636)
);

NAND3xp33_ASAP7_75t_L g6637 ( 
.A(n_6522),
.B(n_351),
.C(n_352),
.Y(n_6637)
);

NAND3xp33_ASAP7_75t_L g6638 ( 
.A(n_6522),
.B(n_353),
.C(n_354),
.Y(n_6638)
);

CKINVDCx5p33_ASAP7_75t_R g6639 ( 
.A(n_6402),
.Y(n_6639)
);

OAI33xp33_ASAP7_75t_L g6640 ( 
.A1(n_6318),
.A2(n_356),
.A3(n_358),
.B1(n_354),
.B2(n_355),
.B3(n_357),
.Y(n_6640)
);

AOI22xp5_ASAP7_75t_L g6641 ( 
.A1(n_6466),
.A2(n_358),
.B1(n_355),
.B2(n_357),
.Y(n_6641)
);

AND2x2_ASAP7_75t_L g6642 ( 
.A(n_6322),
.B(n_359),
.Y(n_6642)
);

OR2x2_ASAP7_75t_L g6643 ( 
.A(n_6296),
.B(n_6502),
.Y(n_6643)
);

AND2x2_ASAP7_75t_L g6644 ( 
.A(n_6328),
.B(n_359),
.Y(n_6644)
);

NAND2xp5_ASAP7_75t_L g6645 ( 
.A(n_6449),
.B(n_360),
.Y(n_6645)
);

INVx2_ASAP7_75t_L g6646 ( 
.A(n_6440),
.Y(n_6646)
);

AOI22xp33_ASAP7_75t_L g6647 ( 
.A1(n_6436),
.A2(n_2443),
.B1(n_2448),
.B2(n_2431),
.Y(n_6647)
);

AOI22xp5_ASAP7_75t_L g6648 ( 
.A1(n_6495),
.A2(n_6502),
.B1(n_6526),
.B2(n_6517),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6474),
.Y(n_6649)
);

OAI22xp5_ASAP7_75t_L g6650 ( 
.A1(n_6526),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_6650)
);

INVx1_ASAP7_75t_L g6651 ( 
.A(n_6414),
.Y(n_6651)
);

AOI33xp33_ASAP7_75t_L g6652 ( 
.A1(n_6503),
.A2(n_365),
.A3(n_367),
.B1(n_361),
.B2(n_363),
.B3(n_366),
.Y(n_6652)
);

OAI221xp5_ASAP7_75t_L g6653 ( 
.A1(n_6457),
.A2(n_366),
.B1(n_363),
.B2(n_365),
.C(n_367),
.Y(n_6653)
);

AOI221xp5_ASAP7_75t_L g6654 ( 
.A1(n_6482),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.C(n_371),
.Y(n_6654)
);

AOI22xp33_ASAP7_75t_L g6655 ( 
.A1(n_6436),
.A2(n_2443),
.B1(n_2448),
.B2(n_2431),
.Y(n_6655)
);

OAI211xp5_ASAP7_75t_L g6656 ( 
.A1(n_6338),
.A2(n_370),
.B(n_368),
.C(n_369),
.Y(n_6656)
);

INVx2_ASAP7_75t_L g6657 ( 
.A(n_6440),
.Y(n_6657)
);

INVx2_ASAP7_75t_L g6658 ( 
.A(n_6282),
.Y(n_6658)
);

NAND2xp5_ASAP7_75t_L g6659 ( 
.A(n_6449),
.B(n_372),
.Y(n_6659)
);

AND2x2_ASAP7_75t_L g6660 ( 
.A(n_6398),
.B(n_373),
.Y(n_6660)
);

AND2x2_ASAP7_75t_L g6661 ( 
.A(n_6311),
.B(n_373),
.Y(n_6661)
);

OAI33xp33_ASAP7_75t_L g6662 ( 
.A1(n_6507),
.A2(n_6516),
.A3(n_6349),
.B1(n_6450),
.B2(n_6499),
.B3(n_6497),
.Y(n_6662)
);

NOR2x1_ASAP7_75t_SL g6663 ( 
.A(n_6308),
.B(n_375),
.Y(n_6663)
);

BUFx3_ASAP7_75t_L g6664 ( 
.A(n_6402),
.Y(n_6664)
);

INVx4_ASAP7_75t_SL g6665 ( 
.A(n_6350),
.Y(n_6665)
);

BUFx3_ASAP7_75t_L g6666 ( 
.A(n_6350),
.Y(n_6666)
);

AOI221xp5_ASAP7_75t_SL g6667 ( 
.A1(n_6397),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.C(n_379),
.Y(n_6667)
);

AOI22xp33_ASAP7_75t_L g6668 ( 
.A1(n_6514),
.A2(n_2448),
.B1(n_2373),
.B2(n_2379),
.Y(n_6668)
);

OA222x2_ASAP7_75t_L g6669 ( 
.A1(n_6420),
.A2(n_381),
.B1(n_385),
.B2(n_378),
.C1(n_380),
.C2(n_384),
.Y(n_6669)
);

OAI22xp5_ASAP7_75t_L g6670 ( 
.A1(n_6397),
.A2(n_386),
.B1(n_380),
.B2(n_384),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_6387),
.Y(n_6671)
);

OAI221xp5_ASAP7_75t_L g6672 ( 
.A1(n_6518),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.C(n_390),
.Y(n_6672)
);

AOI322xp5_ASAP7_75t_L g6673 ( 
.A1(n_6510),
.A2(n_6517),
.A3(n_6500),
.B1(n_6513),
.B2(n_6482),
.C1(n_6505),
.C2(n_6509),
.Y(n_6673)
);

NAND4xp25_ASAP7_75t_L g6674 ( 
.A(n_6374),
.B(n_391),
.C(n_387),
.D(n_388),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_6372),
.Y(n_6675)
);

AND2x4_ASAP7_75t_L g6676 ( 
.A(n_6373),
.B(n_391),
.Y(n_6676)
);

OAI221xp5_ASAP7_75t_L g6677 ( 
.A1(n_6518),
.A2(n_6452),
.B1(n_6446),
.B2(n_6405),
.C(n_6493),
.Y(n_6677)
);

NAND2x1p5_ASAP7_75t_L g6678 ( 
.A(n_6329),
.B(n_392),
.Y(n_6678)
);

OAI221xp5_ASAP7_75t_SL g6679 ( 
.A1(n_6447),
.A2(n_396),
.B1(n_393),
.B2(n_394),
.C(n_397),
.Y(n_6679)
);

BUFx3_ASAP7_75t_L g6680 ( 
.A(n_6350),
.Y(n_6680)
);

OAI221xp5_ASAP7_75t_L g6681 ( 
.A1(n_6452),
.A2(n_399),
.B1(n_396),
.B2(n_398),
.C(n_400),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_6282),
.Y(n_6682)
);

AND2x2_ASAP7_75t_L g6683 ( 
.A(n_6302),
.B(n_6411),
.Y(n_6683)
);

INVx3_ASAP7_75t_L g6684 ( 
.A(n_6329),
.Y(n_6684)
);

AOI21xp5_ASAP7_75t_L g6685 ( 
.A1(n_6374),
.A2(n_398),
.B(n_399),
.Y(n_6685)
);

AND2x2_ASAP7_75t_L g6686 ( 
.A(n_6346),
.B(n_400),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6375),
.Y(n_6687)
);

INVx2_ASAP7_75t_L g6688 ( 
.A(n_6335),
.Y(n_6688)
);

OA21x2_ASAP7_75t_L g6689 ( 
.A1(n_6288),
.A2(n_401),
.B(n_402),
.Y(n_6689)
);

OAI22xp5_ASAP7_75t_L g6690 ( 
.A1(n_6525),
.A2(n_6501),
.B1(n_6509),
.B2(n_6505),
.Y(n_6690)
);

INVx1_ASAP7_75t_L g6691 ( 
.A(n_6380),
.Y(n_6691)
);

OAI21xp5_ASAP7_75t_L g6692 ( 
.A1(n_6501),
.A2(n_401),
.B(n_403),
.Y(n_6692)
);

INVx2_ASAP7_75t_L g6693 ( 
.A(n_6438),
.Y(n_6693)
);

OR2x2_ASAP7_75t_L g6694 ( 
.A(n_6286),
.B(n_403),
.Y(n_6694)
);

AND2x2_ASAP7_75t_L g6695 ( 
.A(n_6347),
.B(n_404),
.Y(n_6695)
);

AOI22xp33_ASAP7_75t_L g6696 ( 
.A1(n_6326),
.A2(n_6469),
.B1(n_6525),
.B2(n_6492),
.Y(n_6696)
);

AOI22xp33_ASAP7_75t_L g6697 ( 
.A1(n_6326),
.A2(n_2448),
.B1(n_2373),
.B2(n_2379),
.Y(n_6697)
);

OA21x2_ASAP7_75t_L g6698 ( 
.A1(n_6288),
.A2(n_407),
.B(n_408),
.Y(n_6698)
);

NAND4xp25_ASAP7_75t_L g6699 ( 
.A(n_6324),
.B(n_410),
.C(n_408),
.D(n_409),
.Y(n_6699)
);

INVx2_ASAP7_75t_L g6700 ( 
.A(n_6438),
.Y(n_6700)
);

AOI221xp5_ASAP7_75t_L g6701 ( 
.A1(n_6479),
.A2(n_6484),
.B1(n_6511),
.B2(n_6423),
.C(n_6508),
.Y(n_6701)
);

AOI211xp5_ASAP7_75t_SL g6702 ( 
.A1(n_6307),
.A2(n_411),
.B(n_409),
.C(n_410),
.Y(n_6702)
);

AOI221xp5_ASAP7_75t_L g6703 ( 
.A1(n_6423),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.C(n_415),
.Y(n_6703)
);

INVx2_ASAP7_75t_L g6704 ( 
.A(n_6329),
.Y(n_6704)
);

AOI21xp5_ASAP7_75t_L g6705 ( 
.A1(n_6488),
.A2(n_412),
.B(n_413),
.Y(n_6705)
);

NAND4xp25_ASAP7_75t_SL g6706 ( 
.A(n_6500),
.B(n_416),
.C(n_414),
.D(n_415),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6404),
.Y(n_6707)
);

OAI22xp5_ASAP7_75t_L g6708 ( 
.A1(n_6513),
.A2(n_420),
.B1(n_417),
.B2(n_419),
.Y(n_6708)
);

OR2x2_ASAP7_75t_L g6709 ( 
.A(n_6392),
.B(n_420),
.Y(n_6709)
);

AOI33xp33_ASAP7_75t_L g6710 ( 
.A1(n_6423),
.A2(n_421),
.A3(n_422),
.B1(n_423),
.B2(n_425),
.B3(n_427),
.Y(n_6710)
);

OAI21x1_ASAP7_75t_L g6711 ( 
.A1(n_6400),
.A2(n_421),
.B(n_423),
.Y(n_6711)
);

CKINVDCx8_ASAP7_75t_R g6712 ( 
.A(n_6329),
.Y(n_6712)
);

OAI21xp5_ASAP7_75t_L g6713 ( 
.A1(n_6488),
.A2(n_427),
.B(n_428),
.Y(n_6713)
);

NAND2xp5_ASAP7_75t_L g6714 ( 
.A(n_6470),
.B(n_429),
.Y(n_6714)
);

AND2x2_ASAP7_75t_L g6715 ( 
.A(n_6364),
.B(n_429),
.Y(n_6715)
);

OR2x2_ASAP7_75t_L g6716 ( 
.A(n_6404),
.B(n_430),
.Y(n_6716)
);

AND2x2_ASAP7_75t_L g6717 ( 
.A(n_6343),
.B(n_430),
.Y(n_6717)
);

OR2x2_ASAP7_75t_L g6718 ( 
.A(n_6373),
.B(n_6332),
.Y(n_6718)
);

NAND4xp25_ASAP7_75t_L g6719 ( 
.A(n_6427),
.B(n_433),
.C(n_431),
.D(n_432),
.Y(n_6719)
);

AOI22xp33_ASAP7_75t_L g6720 ( 
.A1(n_6492),
.A2(n_6464),
.B1(n_6491),
.B2(n_6485),
.Y(n_6720)
);

OAI22xp33_ASAP7_75t_L g6721 ( 
.A1(n_6524),
.A2(n_441),
.B1(n_431),
.B2(n_439),
.Y(n_6721)
);

AOI22xp5_ASAP7_75t_L g6722 ( 
.A1(n_6451),
.A2(n_442),
.B1(n_439),
.B2(n_441),
.Y(n_6722)
);

NAND2x1p5_ASAP7_75t_L g6723 ( 
.A(n_6473),
.B(n_443),
.Y(n_6723)
);

OA222x2_ASAP7_75t_L g6724 ( 
.A1(n_6428),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.C1(n_449),
.C2(n_450),
.Y(n_6724)
);

INVx2_ASAP7_75t_L g6725 ( 
.A(n_6403),
.Y(n_6725)
);

INVx2_ASAP7_75t_L g6726 ( 
.A(n_6399),
.Y(n_6726)
);

NOR2x1_ASAP7_75t_L g6727 ( 
.A(n_6307),
.B(n_445),
.Y(n_6727)
);

INVx1_ASAP7_75t_L g6728 ( 
.A(n_6395),
.Y(n_6728)
);

OAI221xp5_ASAP7_75t_L g6729 ( 
.A1(n_6493),
.A2(n_6477),
.B1(n_6441),
.B2(n_6483),
.C(n_6406),
.Y(n_6729)
);

INVx1_ASAP7_75t_L g6730 ( 
.A(n_6395),
.Y(n_6730)
);

OA21x2_ASAP7_75t_L g6731 ( 
.A1(n_6290),
.A2(n_446),
.B(n_451),
.Y(n_6731)
);

OAI211xp5_ASAP7_75t_L g6732 ( 
.A1(n_6424),
.A2(n_453),
.B(n_451),
.C(n_452),
.Y(n_6732)
);

AOI221xp5_ASAP7_75t_L g6733 ( 
.A1(n_6488),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.C(n_458),
.Y(n_6733)
);

INVx2_ASAP7_75t_L g6734 ( 
.A(n_6443),
.Y(n_6734)
);

NAND2xp5_ASAP7_75t_L g6735 ( 
.A(n_6357),
.B(n_455),
.Y(n_6735)
);

NAND2xp5_ASAP7_75t_L g6736 ( 
.A(n_6357),
.B(n_456),
.Y(n_6736)
);

AND2x2_ASAP7_75t_L g6737 ( 
.A(n_6298),
.B(n_457),
.Y(n_6737)
);

OR2x2_ASAP7_75t_L g6738 ( 
.A(n_6353),
.B(n_459),
.Y(n_6738)
);

INVx2_ASAP7_75t_L g6739 ( 
.A(n_6443),
.Y(n_6739)
);

AOI21xp33_ASAP7_75t_SL g6740 ( 
.A1(n_6285),
.A2(n_6300),
.B(n_6441),
.Y(n_6740)
);

INVx1_ASAP7_75t_L g6741 ( 
.A(n_6415),
.Y(n_6741)
);

AOI22xp33_ASAP7_75t_L g6742 ( 
.A1(n_6464),
.A2(n_2448),
.B1(n_2373),
.B2(n_2379),
.Y(n_6742)
);

INVx1_ASAP7_75t_L g6743 ( 
.A(n_6317),
.Y(n_6743)
);

OR2x2_ASAP7_75t_L g6744 ( 
.A(n_6357),
.B(n_459),
.Y(n_6744)
);

OAI31xp33_ASAP7_75t_L g6745 ( 
.A1(n_6477),
.A2(n_462),
.A3(n_460),
.B(n_461),
.Y(n_6745)
);

AND2x4_ASAP7_75t_SL g6746 ( 
.A(n_6334),
.B(n_460),
.Y(n_6746)
);

OR2x2_ASAP7_75t_L g6747 ( 
.A(n_6357),
.B(n_462),
.Y(n_6747)
);

INVx2_ASAP7_75t_SL g6748 ( 
.A(n_6294),
.Y(n_6748)
);

OAI22xp5_ASAP7_75t_L g6749 ( 
.A1(n_6385),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_6749)
);

OA21x2_ASAP7_75t_L g6750 ( 
.A1(n_6290),
.A2(n_466),
.B(n_467),
.Y(n_6750)
);

AOI22xp33_ASAP7_75t_L g6751 ( 
.A1(n_6489),
.A2(n_6468),
.B1(n_6437),
.B2(n_6481),
.Y(n_6751)
);

INVx2_ASAP7_75t_L g6752 ( 
.A(n_6445),
.Y(n_6752)
);

AND2x2_ASAP7_75t_L g6753 ( 
.A(n_6287),
.B(n_466),
.Y(n_6753)
);

AND2x2_ASAP7_75t_L g6754 ( 
.A(n_6401),
.B(n_467),
.Y(n_6754)
);

OAI221xp5_ASAP7_75t_L g6755 ( 
.A1(n_6473),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.C(n_472),
.Y(n_6755)
);

INVx2_ASAP7_75t_L g6756 ( 
.A(n_6445),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_L g6757 ( 
.A(n_6538),
.B(n_6317),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6606),
.Y(n_6758)
);

AND2x2_ASAP7_75t_L g6759 ( 
.A(n_6666),
.B(n_6334),
.Y(n_6759)
);

AND2x4_ASAP7_75t_SL g6760 ( 
.A(n_6539),
.B(n_6426),
.Y(n_6760)
);

AND2x2_ASAP7_75t_L g6761 ( 
.A(n_6680),
.B(n_6300),
.Y(n_6761)
);

INVx1_ASAP7_75t_L g6762 ( 
.A(n_6605),
.Y(n_6762)
);

NAND2xp5_ASAP7_75t_L g6763 ( 
.A(n_6538),
.B(n_6323),
.Y(n_6763)
);

INVx1_ASAP7_75t_SL g6764 ( 
.A(n_6599),
.Y(n_6764)
);

NAND2xp5_ASAP7_75t_L g6765 ( 
.A(n_6566),
.B(n_6323),
.Y(n_6765)
);

AND2x2_ASAP7_75t_L g6766 ( 
.A(n_6629),
.B(n_6382),
.Y(n_6766)
);

BUFx3_ASAP7_75t_L g6767 ( 
.A(n_6664),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6689),
.Y(n_6768)
);

NAND2xp5_ASAP7_75t_L g6769 ( 
.A(n_6534),
.B(n_6378),
.Y(n_6769)
);

AND2x2_ASAP7_75t_L g6770 ( 
.A(n_6547),
.B(n_6386),
.Y(n_6770)
);

AND2x4_ASAP7_75t_L g6771 ( 
.A(n_6665),
.B(n_6385),
.Y(n_6771)
);

NOR2xp67_ASAP7_75t_L g6772 ( 
.A(n_6555),
.B(n_6385),
.Y(n_6772)
);

INVx1_ASAP7_75t_L g6773 ( 
.A(n_6707),
.Y(n_6773)
);

HB1xp67_ASAP7_75t_L g6774 ( 
.A(n_6567),
.Y(n_6774)
);

INVx2_ASAP7_75t_L g6775 ( 
.A(n_6689),
.Y(n_6775)
);

NAND2xp5_ASAP7_75t_L g6776 ( 
.A(n_6534),
.B(n_6535),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_6623),
.Y(n_6777)
);

INVx1_ASAP7_75t_L g6778 ( 
.A(n_6595),
.Y(n_6778)
);

AND2x2_ASAP7_75t_L g6779 ( 
.A(n_6631),
.B(n_6444),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_6596),
.Y(n_6780)
);

INVx1_ASAP7_75t_L g6781 ( 
.A(n_6610),
.Y(n_6781)
);

INVx1_ASAP7_75t_L g6782 ( 
.A(n_6651),
.Y(n_6782)
);

AND2x2_ASAP7_75t_L g6783 ( 
.A(n_6569),
.B(n_6312),
.Y(n_6783)
);

OR2x2_ASAP7_75t_L g6784 ( 
.A(n_6643),
.B(n_6369),
.Y(n_6784)
);

AND2x2_ASAP7_75t_L g6785 ( 
.A(n_6602),
.B(n_6683),
.Y(n_6785)
);

HB1xp67_ASAP7_75t_L g6786 ( 
.A(n_6594),
.Y(n_6786)
);

INVx3_ASAP7_75t_L g6787 ( 
.A(n_6712),
.Y(n_6787)
);

INVx2_ASAP7_75t_L g6788 ( 
.A(n_6698),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_6671),
.Y(n_6789)
);

AND2x2_ASAP7_75t_L g6790 ( 
.A(n_6621),
.B(n_6342),
.Y(n_6790)
);

INVx2_ASAP7_75t_SL g6791 ( 
.A(n_6746),
.Y(n_6791)
);

INVx2_ASAP7_75t_L g6792 ( 
.A(n_6698),
.Y(n_6792)
);

AND2x2_ASAP7_75t_L g6793 ( 
.A(n_6665),
.B(n_6368),
.Y(n_6793)
);

INVxp33_ASAP7_75t_L g6794 ( 
.A(n_6570),
.Y(n_6794)
);

AND2x2_ASAP7_75t_L g6795 ( 
.A(n_6748),
.B(n_6367),
.Y(n_6795)
);

AND2x2_ASAP7_75t_L g6796 ( 
.A(n_6661),
.B(n_6319),
.Y(n_6796)
);

INVx2_ASAP7_75t_L g6797 ( 
.A(n_6731),
.Y(n_6797)
);

INVx2_ASAP7_75t_L g6798 ( 
.A(n_6731),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_6529),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_6531),
.Y(n_6800)
);

AND2x2_ASAP7_75t_L g6801 ( 
.A(n_6663),
.B(n_6319),
.Y(n_6801)
);

NAND2xp5_ASAP7_75t_L g6802 ( 
.A(n_6632),
.B(n_6378),
.Y(n_6802)
);

NAND2xp5_ASAP7_75t_L g6803 ( 
.A(n_6528),
.B(n_6379),
.Y(n_6803)
);

INVx2_ASAP7_75t_L g6804 ( 
.A(n_6750),
.Y(n_6804)
);

INVx2_ASAP7_75t_L g6805 ( 
.A(n_6750),
.Y(n_6805)
);

NAND2xp5_ASAP7_75t_L g6806 ( 
.A(n_6528),
.B(n_6379),
.Y(n_6806)
);

AND2x4_ASAP7_75t_L g6807 ( 
.A(n_6573),
.B(n_6319),
.Y(n_6807)
);

AND2x2_ASAP7_75t_L g6808 ( 
.A(n_6658),
.B(n_6409),
.Y(n_6808)
);

NAND2x1p5_ASAP7_75t_L g6809 ( 
.A(n_6727),
.B(n_6458),
.Y(n_6809)
);

HB1xp67_ASAP7_75t_L g6810 ( 
.A(n_6637),
.Y(n_6810)
);

INVx1_ASAP7_75t_SL g6811 ( 
.A(n_6639),
.Y(n_6811)
);

INVx2_ASAP7_75t_L g6812 ( 
.A(n_6676),
.Y(n_6812)
);

NAND2xp5_ASAP7_75t_L g6813 ( 
.A(n_6619),
.B(n_6424),
.Y(n_6813)
);

INVx2_ASAP7_75t_L g6814 ( 
.A(n_6676),
.Y(n_6814)
);

INVx1_ASAP7_75t_L g6815 ( 
.A(n_6532),
.Y(n_6815)
);

INVx1_ASAP7_75t_L g6816 ( 
.A(n_6551),
.Y(n_6816)
);

AND2x2_ASAP7_75t_L g6817 ( 
.A(n_6682),
.B(n_6409),
.Y(n_6817)
);

NAND2xp5_ASAP7_75t_L g6818 ( 
.A(n_6654),
.B(n_6331),
.Y(n_6818)
);

AND2x2_ASAP7_75t_L g6819 ( 
.A(n_6642),
.B(n_6417),
.Y(n_6819)
);

AND2x4_ASAP7_75t_L g6820 ( 
.A(n_6586),
.B(n_6366),
.Y(n_6820)
);

AND2x2_ASAP7_75t_L g6821 ( 
.A(n_6644),
.B(n_6417),
.Y(n_6821)
);

INVx1_ASAP7_75t_SL g6822 ( 
.A(n_6576),
.Y(n_6822)
);

INVx2_ASAP7_75t_L g6823 ( 
.A(n_6586),
.Y(n_6823)
);

NAND2xp5_ASAP7_75t_L g6824 ( 
.A(n_6530),
.B(n_6331),
.Y(n_6824)
);

AND2x2_ASAP7_75t_L g6825 ( 
.A(n_6726),
.B(n_6430),
.Y(n_6825)
);

INVx1_ASAP7_75t_L g6826 ( 
.A(n_6553),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_6744),
.Y(n_6827)
);

AND2x4_ASAP7_75t_L g6828 ( 
.A(n_6725),
.B(n_6486),
.Y(n_6828)
);

INVx2_ASAP7_75t_L g6829 ( 
.A(n_6747),
.Y(n_6829)
);

AND2x2_ASAP7_75t_L g6830 ( 
.A(n_6616),
.B(n_6486),
.Y(n_6830)
);

AND2x4_ASAP7_75t_L g6831 ( 
.A(n_6618),
.B(n_6458),
.Y(n_6831)
);

OR2x2_ASAP7_75t_L g6832 ( 
.A(n_6565),
.B(n_6418),
.Y(n_6832)
);

AND2x2_ASAP7_75t_L g6833 ( 
.A(n_6577),
.B(n_6434),
.Y(n_6833)
);

INVx2_ASAP7_75t_L g6834 ( 
.A(n_6678),
.Y(n_6834)
);

OR2x2_ASAP7_75t_L g6835 ( 
.A(n_6581),
.B(n_6418),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_6684),
.Y(n_6836)
);

AND2x2_ASAP7_75t_L g6837 ( 
.A(n_6686),
.B(n_6434),
.Y(n_6837)
);

INVx2_ASAP7_75t_SL g6838 ( 
.A(n_6715),
.Y(n_6838)
);

AND2x2_ASAP7_75t_L g6839 ( 
.A(n_6695),
.B(n_6481),
.Y(n_6839)
);

AND2x2_ASAP7_75t_L g6840 ( 
.A(n_6660),
.B(n_6481),
.Y(n_6840)
);

AND2x4_ASAP7_75t_SL g6841 ( 
.A(n_6753),
.B(n_6475),
.Y(n_6841)
);

AND2x2_ASAP7_75t_L g6842 ( 
.A(n_6704),
.B(n_6432),
.Y(n_6842)
);

INVx1_ASAP7_75t_L g6843 ( 
.A(n_6556),
.Y(n_6843)
);

AND2x2_ASAP7_75t_L g6844 ( 
.A(n_6603),
.B(n_6432),
.Y(n_6844)
);

OR2x2_ASAP7_75t_L g6845 ( 
.A(n_6591),
.B(n_6615),
.Y(n_6845)
);

NAND2x1_ASAP7_75t_L g6846 ( 
.A(n_6684),
.B(n_6458),
.Y(n_6846)
);

AND2x4_ASAP7_75t_L g6847 ( 
.A(n_6754),
.B(n_6453),
.Y(n_6847)
);

AND2x2_ASAP7_75t_L g6848 ( 
.A(n_6737),
.B(n_6527),
.Y(n_6848)
);

HB1xp67_ASAP7_75t_L g6849 ( 
.A(n_6637),
.Y(n_6849)
);

INVxp67_ASAP7_75t_L g6850 ( 
.A(n_6638),
.Y(n_6850)
);

BUFx2_ASAP7_75t_L g6851 ( 
.A(n_6718),
.Y(n_6851)
);

OR2x2_ASAP7_75t_L g6852 ( 
.A(n_6558),
.B(n_6408),
.Y(n_6852)
);

OAI21xp33_ASAP7_75t_L g6853 ( 
.A1(n_6550),
.A2(n_6460),
.B(n_6299),
.Y(n_6853)
);

INVx2_ASAP7_75t_L g6854 ( 
.A(n_6716),
.Y(n_6854)
);

INVx1_ASAP7_75t_L g6855 ( 
.A(n_6562),
.Y(n_6855)
);

NOR2xp33_ASAP7_75t_R g6856 ( 
.A(n_6575),
.B(n_469),
.Y(n_6856)
);

NAND2xp5_ASAP7_75t_L g6857 ( 
.A(n_6638),
.B(n_6673),
.Y(n_6857)
);

NAND2xp33_ASAP7_75t_SL g6858 ( 
.A(n_6626),
.B(n_6453),
.Y(n_6858)
);

INVx2_ASAP7_75t_L g6859 ( 
.A(n_6723),
.Y(n_6859)
);

HB1xp67_ASAP7_75t_L g6860 ( 
.A(n_6634),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6633),
.B(n_6519),
.Y(n_6861)
);

INVx4_ASAP7_75t_L g6862 ( 
.A(n_6717),
.Y(n_6862)
);

NAND2xp5_ASAP7_75t_L g6863 ( 
.A(n_6673),
.B(n_6533),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_6564),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_6571),
.Y(n_6865)
);

OR2x2_ASAP7_75t_L g6866 ( 
.A(n_6741),
.B(n_6408),
.Y(n_6866)
);

INVx1_ASAP7_75t_L g6867 ( 
.A(n_6579),
.Y(n_6867)
);

INVx1_ASAP7_75t_L g6868 ( 
.A(n_6580),
.Y(n_6868)
);

AND2x4_ASAP7_75t_SL g6869 ( 
.A(n_6648),
.B(n_6303),
.Y(n_6869)
);

NAND2xp5_ASAP7_75t_L g6870 ( 
.A(n_6533),
.B(n_6303),
.Y(n_6870)
);

INVxp67_ASAP7_75t_L g6871 ( 
.A(n_6645),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_6588),
.Y(n_6872)
);

INVx2_ASAP7_75t_L g6873 ( 
.A(n_6711),
.Y(n_6873)
);

HB1xp67_ASAP7_75t_L g6874 ( 
.A(n_6593),
.Y(n_6874)
);

AND2x2_ASAP7_75t_L g6875 ( 
.A(n_6694),
.B(n_6460),
.Y(n_6875)
);

AND2x2_ASAP7_75t_L g6876 ( 
.A(n_6624),
.B(n_6738),
.Y(n_6876)
);

NAND2xp5_ASAP7_75t_L g6877 ( 
.A(n_6667),
.B(n_6337),
.Y(n_6877)
);

AND2x2_ASAP7_75t_L g6878 ( 
.A(n_6578),
.B(n_6515),
.Y(n_6878)
);

AND2x2_ASAP7_75t_L g6879 ( 
.A(n_6740),
.B(n_6648),
.Y(n_6879)
);

AND2x2_ASAP7_75t_L g6880 ( 
.A(n_6740),
.B(n_6337),
.Y(n_6880)
);

NOR2x1_ASAP7_75t_L g6881 ( 
.A(n_6674),
.B(n_6299),
.Y(n_6881)
);

INVx2_ASAP7_75t_L g6882 ( 
.A(n_6548),
.Y(n_6882)
);

INVx1_ASAP7_75t_SL g6883 ( 
.A(n_6709),
.Y(n_6883)
);

BUFx3_ASAP7_75t_L g6884 ( 
.A(n_6659),
.Y(n_6884)
);

INVx1_ASAP7_75t_L g6885 ( 
.A(n_6675),
.Y(n_6885)
);

OR2x2_ASAP7_75t_L g6886 ( 
.A(n_6690),
.B(n_6341),
.Y(n_6886)
);

AND2x2_ASAP7_75t_L g6887 ( 
.A(n_6751),
.B(n_6341),
.Y(n_6887)
);

NAND2xp5_ASAP7_75t_L g6888 ( 
.A(n_6667),
.B(n_6693),
.Y(n_6888)
);

OR2x2_ASAP7_75t_L g6889 ( 
.A(n_6585),
.B(n_6348),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6687),
.Y(n_6890)
);

INVx2_ASAP7_75t_L g6891 ( 
.A(n_6548),
.Y(n_6891)
);

OR2x2_ASAP7_75t_L g6892 ( 
.A(n_6700),
.B(n_6348),
.Y(n_6892)
);

BUFx3_ASAP7_75t_L g6893 ( 
.A(n_6641),
.Y(n_6893)
);

AND2x2_ASAP7_75t_L g6894 ( 
.A(n_6691),
.B(n_6354),
.Y(n_6894)
);

HB1xp67_ASAP7_75t_L g6895 ( 
.A(n_6650),
.Y(n_6895)
);

NAND2xp5_ASAP7_75t_L g6896 ( 
.A(n_6620),
.B(n_6354),
.Y(n_6896)
);

NAND2xp5_ASAP7_75t_L g6897 ( 
.A(n_6554),
.B(n_6389),
.Y(n_6897)
);

AND2x2_ASAP7_75t_L g6898 ( 
.A(n_6669),
.B(n_6355),
.Y(n_6898)
);

INVx1_ASAP7_75t_L g6899 ( 
.A(n_6743),
.Y(n_6899)
);

AOI21xp33_ASAP7_75t_SL g6900 ( 
.A1(n_6607),
.A2(n_470),
.B(n_472),
.Y(n_6900)
);

NOR2xp33_ASAP7_75t_L g6901 ( 
.A(n_6545),
.B(n_6355),
.Y(n_6901)
);

OR2x2_ASAP7_75t_L g6902 ( 
.A(n_6604),
.B(n_6356),
.Y(n_6902)
);

INVx1_ASAP7_75t_L g6903 ( 
.A(n_6728),
.Y(n_6903)
);

INVx2_ASAP7_75t_L g6904 ( 
.A(n_6552),
.Y(n_6904)
);

AND2x2_ASAP7_75t_L g6905 ( 
.A(n_6669),
.B(n_6356),
.Y(n_6905)
);

AND2x2_ASAP7_75t_L g6906 ( 
.A(n_6692),
.B(n_6358),
.Y(n_6906)
);

BUFx2_ASAP7_75t_L g6907 ( 
.A(n_6561),
.Y(n_6907)
);

AND2x4_ASAP7_75t_L g6908 ( 
.A(n_6612),
.B(n_6358),
.Y(n_6908)
);

BUFx2_ASAP7_75t_L g6909 ( 
.A(n_6574),
.Y(n_6909)
);

INVx1_ASAP7_75t_L g6910 ( 
.A(n_6730),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6613),
.Y(n_6911)
);

AND2x4_ASAP7_75t_L g6912 ( 
.A(n_6625),
.B(n_6360),
.Y(n_6912)
);

NAND2xp5_ASAP7_75t_L g6913 ( 
.A(n_6703),
.B(n_6360),
.Y(n_6913)
);

INVxp67_ASAP7_75t_L g6914 ( 
.A(n_6630),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6646),
.Y(n_6915)
);

AND2x2_ASAP7_75t_L g6916 ( 
.A(n_6598),
.B(n_6370),
.Y(n_6916)
);

NAND2xp5_ASAP7_75t_SL g6917 ( 
.A(n_6545),
.B(n_6582),
.Y(n_6917)
);

INVx1_ASAP7_75t_L g6918 ( 
.A(n_6657),
.Y(n_6918)
);

INVx1_ASAP7_75t_L g6919 ( 
.A(n_6714),
.Y(n_6919)
);

BUFx2_ASAP7_75t_L g6920 ( 
.A(n_6719),
.Y(n_6920)
);

INVx1_ASAP7_75t_L g6921 ( 
.A(n_6735),
.Y(n_6921)
);

INVx2_ASAP7_75t_L g6922 ( 
.A(n_6688),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_6736),
.Y(n_6923)
);

NOR2x1p5_ASAP7_75t_L g6924 ( 
.A(n_6719),
.B(n_6370),
.Y(n_6924)
);

INVx1_ASAP7_75t_L g6925 ( 
.A(n_6628),
.Y(n_6925)
);

OR2x2_ASAP7_75t_L g6926 ( 
.A(n_6649),
.B(n_6371),
.Y(n_6926)
);

AND2x2_ASAP7_75t_L g6927 ( 
.A(n_6724),
.B(n_6371),
.Y(n_6927)
);

NAND2xp5_ASAP7_75t_L g6928 ( 
.A(n_6710),
.B(n_6389),
.Y(n_6928)
);

AND2x2_ASAP7_75t_L g6929 ( 
.A(n_6724),
.B(n_6383),
.Y(n_6929)
);

INVx2_ASAP7_75t_L g6930 ( 
.A(n_6734),
.Y(n_6930)
);

OR2x2_ASAP7_75t_L g6931 ( 
.A(n_6542),
.B(n_6383),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_6628),
.Y(n_6932)
);

AND2x4_ASAP7_75t_SL g6933 ( 
.A(n_6641),
.B(n_6384),
.Y(n_6933)
);

HB1xp67_ASAP7_75t_L g6934 ( 
.A(n_6583),
.Y(n_6934)
);

INVx2_ASAP7_75t_L g6935 ( 
.A(n_6739),
.Y(n_6935)
);

OR2x2_ASAP7_75t_L g6936 ( 
.A(n_6542),
.B(n_6384),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_6708),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6635),
.Y(n_6938)
);

NOR2xp67_ASAP7_75t_L g6939 ( 
.A(n_6706),
.B(n_473),
.Y(n_6939)
);

OAI31xp33_ASAP7_75t_L g6940 ( 
.A1(n_6863),
.A2(n_6537),
.A3(n_6699),
.B(n_6674),
.Y(n_6940)
);

INVx2_ASAP7_75t_L g6941 ( 
.A(n_6767),
.Y(n_6941)
);

OAI322xp33_ASAP7_75t_L g6942 ( 
.A1(n_6863),
.A2(n_6729),
.A3(n_6622),
.B1(n_6677),
.B2(n_6600),
.C1(n_6685),
.C2(n_6592),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6874),
.Y(n_6943)
);

AND2x4_ASAP7_75t_L g6944 ( 
.A(n_6767),
.B(n_6713),
.Y(n_6944)
);

INVx2_ASAP7_75t_L g6945 ( 
.A(n_6862),
.Y(n_6945)
);

OAI31xp33_ASAP7_75t_L g6946 ( 
.A1(n_6857),
.A2(n_6699),
.A3(n_6584),
.B(n_6568),
.Y(n_6946)
);

HB1xp67_ASAP7_75t_L g6947 ( 
.A(n_6764),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_6874),
.Y(n_6948)
);

INVx2_ASAP7_75t_SL g6949 ( 
.A(n_6771),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_6860),
.Y(n_6950)
);

BUFx2_ASAP7_75t_L g6951 ( 
.A(n_6771),
.Y(n_6951)
);

NAND2xp5_ASAP7_75t_SL g6952 ( 
.A(n_6820),
.B(n_6563),
.Y(n_6952)
);

AND2x2_ASAP7_75t_L g6953 ( 
.A(n_6785),
.B(n_6702),
.Y(n_6953)
);

NAND2xp5_ASAP7_75t_L g6954 ( 
.A(n_6920),
.B(n_6627),
.Y(n_6954)
);

AOI221xp5_ASAP7_75t_L g6955 ( 
.A1(n_6776),
.A2(n_6662),
.B1(n_6701),
.B2(n_6640),
.C(n_6611),
.Y(n_6955)
);

AND2x4_ASAP7_75t_L g6956 ( 
.A(n_6820),
.B(n_6583),
.Y(n_6956)
);

AND2x2_ASAP7_75t_L g6957 ( 
.A(n_6764),
.B(n_6635),
.Y(n_6957)
);

NAND4xp25_ASAP7_75t_L g6958 ( 
.A(n_6776),
.B(n_6563),
.C(n_6597),
.D(n_6652),
.Y(n_6958)
);

HB1xp67_ASAP7_75t_L g6959 ( 
.A(n_6810),
.Y(n_6959)
);

BUFx3_ASAP7_75t_L g6960 ( 
.A(n_6791),
.Y(n_6960)
);

OAI31xp33_ASAP7_75t_L g6961 ( 
.A1(n_6857),
.A2(n_6679),
.A3(n_6672),
.B(n_6732),
.Y(n_6961)
);

OAI33xp33_ASAP7_75t_L g6962 ( 
.A1(n_6757),
.A2(n_6617),
.A3(n_6636),
.B1(n_6721),
.B2(n_6557),
.B3(n_6670),
.Y(n_6962)
);

INVx1_ASAP7_75t_L g6963 ( 
.A(n_6860),
.Y(n_6963)
);

INVx4_ASAP7_75t_L g6964 ( 
.A(n_6787),
.Y(n_6964)
);

AOI22xp33_ASAP7_75t_L g6965 ( 
.A1(n_6870),
.A2(n_6543),
.B1(n_6696),
.B2(n_6720),
.Y(n_6965)
);

INVx2_ASAP7_75t_L g6966 ( 
.A(n_6862),
.Y(n_6966)
);

OAI211xp5_ASAP7_75t_L g6967 ( 
.A1(n_6879),
.A2(n_6656),
.B(n_6587),
.C(n_6733),
.Y(n_6967)
);

INVx2_ASAP7_75t_L g6968 ( 
.A(n_6841),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_SL g6969 ( 
.A(n_6809),
.B(n_6745),
.Y(n_6969)
);

NAND2xp5_ASAP7_75t_SL g6970 ( 
.A(n_6809),
.B(n_6745),
.Y(n_6970)
);

AND2x2_ASAP7_75t_L g6971 ( 
.A(n_6801),
.B(n_6572),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_6926),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6866),
.Y(n_6973)
);

NAND2xp5_ASAP7_75t_L g6974 ( 
.A(n_6883),
.B(n_6786),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6777),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_6796),
.B(n_6722),
.Y(n_6976)
);

INVx2_ASAP7_75t_L g6977 ( 
.A(n_6869),
.Y(n_6977)
);

NAND3xp33_ASAP7_75t_L g6978 ( 
.A(n_6810),
.B(n_6560),
.C(n_6749),
.Y(n_6978)
);

AND2x2_ASAP7_75t_L g6979 ( 
.A(n_6783),
.B(n_6722),
.Y(n_6979)
);

AND2x2_ASAP7_75t_L g6980 ( 
.A(n_6766),
.B(n_6705),
.Y(n_6980)
);

INVx2_ASAP7_75t_L g6981 ( 
.A(n_6838),
.Y(n_6981)
);

AOI211xp5_ASAP7_75t_L g6982 ( 
.A1(n_6849),
.A2(n_6559),
.B(n_6681),
.C(n_6653),
.Y(n_6982)
);

HB1xp67_ASAP7_75t_L g6983 ( 
.A(n_6849),
.Y(n_6983)
);

INVx1_ASAP7_75t_L g6984 ( 
.A(n_6758),
.Y(n_6984)
);

AOI22xp33_ASAP7_75t_L g6985 ( 
.A1(n_6870),
.A2(n_6543),
.B1(n_6536),
.B2(n_6540),
.Y(n_6985)
);

NAND2xp5_ASAP7_75t_L g6986 ( 
.A(n_6883),
.B(n_6786),
.Y(n_6986)
);

INVx2_ASAP7_75t_L g6987 ( 
.A(n_6807),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_6894),
.Y(n_6988)
);

NAND2xp5_ASAP7_75t_L g6989 ( 
.A(n_6850),
.B(n_6589),
.Y(n_6989)
);

NAND5xp2_ASAP7_75t_L g6990 ( 
.A(n_6793),
.B(n_6755),
.C(n_6546),
.D(n_6549),
.E(n_6609),
.Y(n_6990)
);

AOI21xp5_ASAP7_75t_L g6991 ( 
.A1(n_6917),
.A2(n_6559),
.B(n_6544),
.Y(n_6991)
);

AND2x2_ASAP7_75t_L g6992 ( 
.A(n_6819),
.B(n_6752),
.Y(n_6992)
);

NAND2x1_ASAP7_75t_L g6993 ( 
.A(n_6831),
.B(n_6756),
.Y(n_6993)
);

OR2x2_ASAP7_75t_L g6994 ( 
.A(n_6774),
.B(n_6590),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6851),
.Y(n_6995)
);

NAND2xp5_ASAP7_75t_L g6996 ( 
.A(n_6850),
.B(n_6822),
.Y(n_6996)
);

AOI221xp5_ASAP7_75t_L g6997 ( 
.A1(n_6900),
.A2(n_6655),
.B1(n_6647),
.B2(n_6608),
.C(n_6601),
.Y(n_6997)
);

INVx1_ASAP7_75t_L g6998 ( 
.A(n_6934),
.Y(n_6998)
);

AND2x2_ASAP7_75t_L g6999 ( 
.A(n_6821),
.B(n_6541),
.Y(n_6999)
);

NAND4xp25_ASAP7_75t_L g7000 ( 
.A(n_6757),
.B(n_6742),
.C(n_6668),
.D(n_6614),
.Y(n_7000)
);

INVxp67_ASAP7_75t_L g7001 ( 
.A(n_6774),
.Y(n_7001)
);

AND2x2_ASAP7_75t_L g7002 ( 
.A(n_6787),
.B(n_6541),
.Y(n_7002)
);

INVx2_ASAP7_75t_SL g7003 ( 
.A(n_6831),
.Y(n_7003)
);

INVx3_ASAP7_75t_L g7004 ( 
.A(n_6807),
.Y(n_7004)
);

OR2x2_ASAP7_75t_L g7005 ( 
.A(n_6888),
.B(n_6697),
.Y(n_7005)
);

INVx5_ASAP7_75t_L g7006 ( 
.A(n_6759),
.Y(n_7006)
);

AND2x2_ASAP7_75t_L g7007 ( 
.A(n_6770),
.B(n_474),
.Y(n_7007)
);

NAND2xp5_ASAP7_75t_L g7008 ( 
.A(n_6822),
.B(n_474),
.Y(n_7008)
);

NOR3xp33_ASAP7_75t_SL g7009 ( 
.A(n_6763),
.B(n_475),
.C(n_476),
.Y(n_7009)
);

INVx2_ASAP7_75t_L g7010 ( 
.A(n_6845),
.Y(n_7010)
);

OAI211xp5_ASAP7_75t_L g7011 ( 
.A1(n_6763),
.A2(n_6769),
.B(n_6888),
.C(n_6772),
.Y(n_7011)
);

INVx1_ASAP7_75t_L g7012 ( 
.A(n_6934),
.Y(n_7012)
);

OR2x2_ASAP7_75t_L g7013 ( 
.A(n_6877),
.B(n_475),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6903),
.Y(n_7014)
);

BUFx2_ASAP7_75t_L g7015 ( 
.A(n_6839),
.Y(n_7015)
);

AND2x2_ASAP7_75t_L g7016 ( 
.A(n_6840),
.B(n_479),
.Y(n_7016)
);

INVx1_ASAP7_75t_L g7017 ( 
.A(n_6910),
.Y(n_7017)
);

INVx2_ASAP7_75t_L g7018 ( 
.A(n_6823),
.Y(n_7018)
);

AND2x4_ASAP7_75t_L g7019 ( 
.A(n_6812),
.B(n_479),
.Y(n_7019)
);

NAND2xp5_ASAP7_75t_L g7020 ( 
.A(n_6924),
.B(n_480),
.Y(n_7020)
);

INVx2_ASAP7_75t_SL g7021 ( 
.A(n_6760),
.Y(n_7021)
);

NAND2xp5_ASAP7_75t_L g7022 ( 
.A(n_6895),
.B(n_480),
.Y(n_7022)
);

AOI22xp33_ASAP7_75t_L g7023 ( 
.A1(n_6927),
.A2(n_2373),
.B1(n_2379),
.B2(n_2372),
.Y(n_7023)
);

OAI211xp5_ASAP7_75t_SL g7024 ( 
.A1(n_6769),
.A2(n_6917),
.B(n_6881),
.C(n_6811),
.Y(n_7024)
);

INVx1_ASAP7_75t_L g7025 ( 
.A(n_6773),
.Y(n_7025)
);

NAND2xp5_ASAP7_75t_L g7026 ( 
.A(n_6895),
.B(n_482),
.Y(n_7026)
);

INVx4_ASAP7_75t_L g7027 ( 
.A(n_6761),
.Y(n_7027)
);

INVx1_ASAP7_75t_L g7028 ( 
.A(n_6799),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6800),
.Y(n_7029)
);

AOI33xp33_ASAP7_75t_L g7030 ( 
.A1(n_6925),
.A2(n_6932),
.A3(n_6780),
.B1(n_6778),
.B2(n_6781),
.B3(n_6887),
.Y(n_7030)
);

INVx3_ASAP7_75t_L g7031 ( 
.A(n_6846),
.Y(n_7031)
);

INVx2_ASAP7_75t_L g7032 ( 
.A(n_6852),
.Y(n_7032)
);

HB1xp67_ASAP7_75t_L g7033 ( 
.A(n_6814),
.Y(n_7033)
);

INVx1_ASAP7_75t_L g7034 ( 
.A(n_6815),
.Y(n_7034)
);

AND2x4_ASAP7_75t_L g7035 ( 
.A(n_6795),
.B(n_482),
.Y(n_7035)
);

NAND2xp5_ASAP7_75t_L g7036 ( 
.A(n_6884),
.B(n_484),
.Y(n_7036)
);

INVx2_ASAP7_75t_L g7037 ( 
.A(n_6847),
.Y(n_7037)
);

OAI211xp5_ASAP7_75t_SL g7038 ( 
.A1(n_6811),
.A2(n_6824),
.B(n_6806),
.C(n_6803),
.Y(n_7038)
);

OAI31xp33_ASAP7_75t_L g7039 ( 
.A1(n_6914),
.A2(n_486),
.A3(n_484),
.B(n_485),
.Y(n_7039)
);

OAI221xp5_ASAP7_75t_L g7040 ( 
.A1(n_6914),
.A2(n_485),
.B1(n_487),
.B2(n_489),
.C(n_490),
.Y(n_7040)
);

INVxp67_ASAP7_75t_L g7041 ( 
.A(n_6929),
.Y(n_7041)
);

INVx2_ASAP7_75t_L g7042 ( 
.A(n_6847),
.Y(n_7042)
);

OAI21x1_ASAP7_75t_L g7043 ( 
.A1(n_6765),
.A2(n_489),
.B(n_490),
.Y(n_7043)
);

BUFx3_ASAP7_75t_L g7044 ( 
.A(n_6859),
.Y(n_7044)
);

BUFx2_ASAP7_75t_L g7045 ( 
.A(n_6790),
.Y(n_7045)
);

AND2x2_ASAP7_75t_L g7046 ( 
.A(n_6833),
.B(n_491),
.Y(n_7046)
);

AND2x2_ASAP7_75t_L g7047 ( 
.A(n_6837),
.B(n_491),
.Y(n_7047)
);

AOI22xp33_ASAP7_75t_SL g7048 ( 
.A1(n_6898),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6816),
.Y(n_7049)
);

NAND2xp5_ASAP7_75t_L g7050 ( 
.A(n_6876),
.B(n_495),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_6826),
.Y(n_7051)
);

NAND4xp25_ASAP7_75t_L g7052 ( 
.A(n_6803),
.B(n_499),
.C(n_497),
.D(n_498),
.Y(n_7052)
);

INVx1_ASAP7_75t_L g7053 ( 
.A(n_6843),
.Y(n_7053)
);

INVx1_ASAP7_75t_SL g7054 ( 
.A(n_6856),
.Y(n_7054)
);

NAND3xp33_ASAP7_75t_L g7055 ( 
.A(n_6802),
.B(n_6806),
.C(n_6877),
.Y(n_7055)
);

AOI211xp5_ASAP7_75t_L g7056 ( 
.A1(n_6939),
.A2(n_501),
.B(n_497),
.C(n_498),
.Y(n_7056)
);

NAND2xp5_ASAP7_75t_SL g7057 ( 
.A(n_6848),
.B(n_2240),
.Y(n_7057)
);

OR2x2_ASAP7_75t_L g7058 ( 
.A(n_6784),
.B(n_502),
.Y(n_7058)
);

INVx2_ASAP7_75t_L g7059 ( 
.A(n_6844),
.Y(n_7059)
);

NAND4xp25_ASAP7_75t_L g7060 ( 
.A(n_6824),
.B(n_505),
.C(n_503),
.D(n_504),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_6855),
.Y(n_7061)
);

INVx4_ASAP7_75t_L g7062 ( 
.A(n_6907),
.Y(n_7062)
);

AND2x2_ASAP7_75t_L g7063 ( 
.A(n_6779),
.B(n_503),
.Y(n_7063)
);

INVx2_ASAP7_75t_L g7064 ( 
.A(n_6768),
.Y(n_7064)
);

AOI221xp5_ASAP7_75t_L g7065 ( 
.A1(n_6853),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.C(n_508),
.Y(n_7065)
);

OAI211xp5_ASAP7_75t_SL g7066 ( 
.A1(n_6931),
.A2(n_508),
.B(n_506),
.C(n_507),
.Y(n_7066)
);

INVx1_ASAP7_75t_SL g7067 ( 
.A(n_6856),
.Y(n_7067)
);

AND2x2_ASAP7_75t_L g7068 ( 
.A(n_6825),
.B(n_510),
.Y(n_7068)
);

AND2x2_ASAP7_75t_L g7069 ( 
.A(n_6808),
.B(n_510),
.Y(n_7069)
);

OAI21xp33_ASAP7_75t_L g7070 ( 
.A1(n_6794),
.A2(n_512),
.B(n_514),
.Y(n_7070)
);

OR2x2_ASAP7_75t_L g7071 ( 
.A(n_6928),
.B(n_515),
.Y(n_7071)
);

INVx1_ASAP7_75t_L g7072 ( 
.A(n_6864),
.Y(n_7072)
);

BUFx2_ASAP7_75t_L g7073 ( 
.A(n_6909),
.Y(n_7073)
);

INVx1_ASAP7_75t_L g7074 ( 
.A(n_6865),
.Y(n_7074)
);

INVx2_ASAP7_75t_L g7075 ( 
.A(n_6775),
.Y(n_7075)
);

OR2x2_ASAP7_75t_L g7076 ( 
.A(n_6928),
.B(n_516),
.Y(n_7076)
);

AND2x2_ASAP7_75t_L g7077 ( 
.A(n_6817),
.B(n_518),
.Y(n_7077)
);

AND2x2_ASAP7_75t_L g7078 ( 
.A(n_6794),
.B(n_6836),
.Y(n_7078)
);

AND2x2_ASAP7_75t_L g7079 ( 
.A(n_6880),
.B(n_518),
.Y(n_7079)
);

OR2x2_ASAP7_75t_L g7080 ( 
.A(n_6762),
.B(n_519),
.Y(n_7080)
);

OR2x2_ASAP7_75t_L g7081 ( 
.A(n_6897),
.B(n_520),
.Y(n_7081)
);

NAND3xp33_ASAP7_75t_L g7082 ( 
.A(n_6802),
.B(n_521),
.C(n_524),
.Y(n_7082)
);

AND2x4_ASAP7_75t_L g7083 ( 
.A(n_7004),
.B(n_6873),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6959),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6983),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_6947),
.B(n_6919),
.Y(n_7086)
);

AND2x2_ASAP7_75t_L g7087 ( 
.A(n_7015),
.B(n_6842),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_7013),
.Y(n_7088)
);

INVx2_ASAP7_75t_L g7089 ( 
.A(n_7062),
.Y(n_7089)
);

INVx1_ASAP7_75t_L g7090 ( 
.A(n_6974),
.Y(n_7090)
);

INVx2_ASAP7_75t_L g7091 ( 
.A(n_7062),
.Y(n_7091)
);

AND2x2_ASAP7_75t_L g7092 ( 
.A(n_6953),
.B(n_6830),
.Y(n_7092)
);

INVx1_ASAP7_75t_L g7093 ( 
.A(n_6986),
.Y(n_7093)
);

AND2x2_ASAP7_75t_L g7094 ( 
.A(n_6951),
.B(n_7045),
.Y(n_7094)
);

NAND2xp5_ASAP7_75t_L g7095 ( 
.A(n_7069),
.B(n_6871),
.Y(n_7095)
);

INVx1_ASAP7_75t_L g7096 ( 
.A(n_7073),
.Y(n_7096)
);

AND2x2_ASAP7_75t_L g7097 ( 
.A(n_6964),
.B(n_6904),
.Y(n_7097)
);

NOR2xp33_ASAP7_75t_L g7098 ( 
.A(n_6964),
.B(n_6871),
.Y(n_7098)
);

INVx2_ASAP7_75t_L g7099 ( 
.A(n_7004),
.Y(n_7099)
);

INVxp67_ASAP7_75t_L g7100 ( 
.A(n_6960),
.Y(n_7100)
);

OR2x2_ASAP7_75t_L g7101 ( 
.A(n_6996),
.B(n_6897),
.Y(n_7101)
);

INVx2_ASAP7_75t_L g7102 ( 
.A(n_7054),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_7033),
.Y(n_7103)
);

NAND2xp5_ASAP7_75t_L g7104 ( 
.A(n_7077),
.B(n_6905),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_6998),
.Y(n_7105)
);

NAND2xp5_ASAP7_75t_L g7106 ( 
.A(n_7046),
.B(n_6937),
.Y(n_7106)
);

INVx1_ASAP7_75t_L g7107 ( 
.A(n_7012),
.Y(n_7107)
);

AND2x2_ASAP7_75t_L g7108 ( 
.A(n_7027),
.B(n_6782),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6995),
.Y(n_7109)
);

INVxp67_ASAP7_75t_SL g7110 ( 
.A(n_7055),
.Y(n_7110)
);

A2O1A1Ixp33_ASAP7_75t_L g7111 ( 
.A1(n_6946),
.A2(n_6940),
.B(n_6961),
.C(n_7055),
.Y(n_7111)
);

AND2x4_ASAP7_75t_L g7112 ( 
.A(n_6949),
.B(n_6789),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_7064),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_7075),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_7008),
.Y(n_7115)
);

INVx1_ASAP7_75t_L g7116 ( 
.A(n_7010),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_7058),
.Y(n_7117)
);

AOI22xp33_ASAP7_75t_L g7118 ( 
.A1(n_6955),
.A2(n_6936),
.B1(n_6893),
.B2(n_6891),
.Y(n_7118)
);

AND2x4_ASAP7_75t_L g7119 ( 
.A(n_7006),
.B(n_6861),
.Y(n_7119)
);

BUFx2_ASAP7_75t_L g7120 ( 
.A(n_7027),
.Y(n_7120)
);

AND2x2_ASAP7_75t_L g7121 ( 
.A(n_7063),
.B(n_6867),
.Y(n_7121)
);

OR2x2_ASAP7_75t_L g7122 ( 
.A(n_6952),
.B(n_6813),
.Y(n_7122)
);

INVx1_ASAP7_75t_L g7123 ( 
.A(n_7081),
.Y(n_7123)
);

AND2x2_ASAP7_75t_L g7124 ( 
.A(n_7006),
.B(n_6868),
.Y(n_7124)
);

NAND3xp33_ASAP7_75t_L g7125 ( 
.A(n_6940),
.B(n_6765),
.C(n_6901),
.Y(n_7125)
);

INVx1_ASAP7_75t_L g7126 ( 
.A(n_7071),
.Y(n_7126)
);

AND2x2_ASAP7_75t_L g7127 ( 
.A(n_7006),
.B(n_6872),
.Y(n_7127)
);

INVx1_ASAP7_75t_L g7128 ( 
.A(n_7076),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6943),
.Y(n_7129)
);

AND2x4_ASAP7_75t_L g7130 ( 
.A(n_7021),
.B(n_6885),
.Y(n_7130)
);

AND2x4_ASAP7_75t_L g7131 ( 
.A(n_6941),
.B(n_6890),
.Y(n_7131)
);

INVx2_ASAP7_75t_SL g7132 ( 
.A(n_6993),
.Y(n_7132)
);

INVx1_ASAP7_75t_L g7133 ( 
.A(n_7022),
.Y(n_7133)
);

NAND2xp5_ASAP7_75t_L g7134 ( 
.A(n_7047),
.B(n_6901),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_6948),
.Y(n_7135)
);

INVx1_ASAP7_75t_L g7136 ( 
.A(n_7026),
.Y(n_7136)
);

OR2x6_ASAP7_75t_L g7137 ( 
.A(n_7050),
.B(n_6827),
.Y(n_7137)
);

INVxp67_ASAP7_75t_SL g7138 ( 
.A(n_7082),
.Y(n_7138)
);

AND2x2_ASAP7_75t_L g7139 ( 
.A(n_7003),
.B(n_6834),
.Y(n_7139)
);

INVx1_ASAP7_75t_SL g7140 ( 
.A(n_7054),
.Y(n_7140)
);

NAND3xp33_ASAP7_75t_L g7141 ( 
.A(n_7024),
.B(n_6853),
.C(n_6813),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_7035),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_6950),
.Y(n_7143)
);

AND2x4_ASAP7_75t_SL g7144 ( 
.A(n_6968),
.B(n_6829),
.Y(n_7144)
);

INVx1_ASAP7_75t_L g7145 ( 
.A(n_6963),
.Y(n_7145)
);

NOR2xp33_ASAP7_75t_L g7146 ( 
.A(n_7060),
.B(n_6921),
.Y(n_7146)
);

NAND2xp5_ASAP7_75t_L g7147 ( 
.A(n_7048),
.B(n_6878),
.Y(n_7147)
);

NAND2xp5_ASAP7_75t_L g7148 ( 
.A(n_7009),
.B(n_6923),
.Y(n_7148)
);

NAND2xp5_ASAP7_75t_L g7149 ( 
.A(n_7068),
.B(n_6854),
.Y(n_7149)
);

AND2x2_ASAP7_75t_L g7150 ( 
.A(n_6987),
.B(n_6906),
.Y(n_7150)
);

AND2x4_ASAP7_75t_L g7151 ( 
.A(n_7059),
.B(n_6922),
.Y(n_7151)
);

AND2x2_ASAP7_75t_L g7152 ( 
.A(n_7078),
.B(n_6875),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_7036),
.Y(n_7153)
);

NOR3xp33_ASAP7_75t_L g7154 ( 
.A(n_7038),
.B(n_6858),
.C(n_6938),
.Y(n_7154)
);

INVx2_ASAP7_75t_L g7155 ( 
.A(n_7035),
.Y(n_7155)
);

AND2x2_ASAP7_75t_L g7156 ( 
.A(n_6945),
.B(n_6933),
.Y(n_7156)
);

AND2x2_ASAP7_75t_L g7157 ( 
.A(n_6966),
.B(n_6916),
.Y(n_7157)
);

NAND2xp5_ASAP7_75t_L g7158 ( 
.A(n_7007),
.B(n_6911),
.Y(n_7158)
);

INVx1_ASAP7_75t_L g7159 ( 
.A(n_7080),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_6972),
.Y(n_7160)
);

OAI22xp33_ASAP7_75t_L g7161 ( 
.A1(n_6958),
.A2(n_7041),
.B1(n_6896),
.B2(n_6913),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6973),
.Y(n_7162)
);

INVx1_ASAP7_75t_L g7163 ( 
.A(n_7032),
.Y(n_7163)
);

AND3x2_ASAP7_75t_L g7164 ( 
.A(n_7056),
.B(n_7039),
.C(n_7001),
.Y(n_7164)
);

NAND2xp33_ASAP7_75t_R g7165 ( 
.A(n_7079),
.B(n_6896),
.Y(n_7165)
);

AND2x2_ASAP7_75t_L g7166 ( 
.A(n_7016),
.B(n_6899),
.Y(n_7166)
);

INVx2_ASAP7_75t_L g7167 ( 
.A(n_7067),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6957),
.Y(n_7168)
);

NAND2x1p5_ASAP7_75t_L g7169 ( 
.A(n_7019),
.B(n_6832),
.Y(n_7169)
);

OR2x2_ASAP7_75t_L g7170 ( 
.A(n_6988),
.B(n_6818),
.Y(n_7170)
);

NOR2x1_ASAP7_75t_L g7171 ( 
.A(n_7052),
.B(n_6818),
.Y(n_7171)
);

OR2x2_ASAP7_75t_L g7172 ( 
.A(n_6978),
.B(n_6981),
.Y(n_7172)
);

OR2x2_ASAP7_75t_L g7173 ( 
.A(n_6978),
.B(n_6886),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_7018),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_7082),
.Y(n_7175)
);

INVx1_ASAP7_75t_L g7176 ( 
.A(n_7030),
.Y(n_7176)
);

AND2x2_ASAP7_75t_L g7177 ( 
.A(n_6971),
.B(n_6835),
.Y(n_7177)
);

AOI33xp33_ASAP7_75t_L g7178 ( 
.A1(n_6965),
.A2(n_6882),
.A3(n_6918),
.B1(n_6915),
.B2(n_6828),
.B3(n_6797),
.Y(n_7178)
);

INVx2_ASAP7_75t_L g7179 ( 
.A(n_7019),
.Y(n_7179)
);

HB1xp67_ASAP7_75t_L g7180 ( 
.A(n_7044),
.Y(n_7180)
);

OAI21xp5_ASAP7_75t_L g7181 ( 
.A1(n_6969),
.A2(n_6913),
.B(n_6858),
.Y(n_7181)
);

AND2x2_ASAP7_75t_L g7182 ( 
.A(n_6979),
.B(n_6828),
.Y(n_7182)
);

NAND2xp5_ASAP7_75t_L g7183 ( 
.A(n_6946),
.B(n_6889),
.Y(n_7183)
);

NOR2xp33_ASAP7_75t_L g7184 ( 
.A(n_7060),
.B(n_6788),
.Y(n_7184)
);

INVxp67_ASAP7_75t_SL g7185 ( 
.A(n_7056),
.Y(n_7185)
);

INVx1_ASAP7_75t_L g7186 ( 
.A(n_6975),
.Y(n_7186)
);

INVx1_ASAP7_75t_L g7187 ( 
.A(n_6984),
.Y(n_7187)
);

INVx1_ASAP7_75t_L g7188 ( 
.A(n_7014),
.Y(n_7188)
);

OR2x2_ASAP7_75t_L g7189 ( 
.A(n_6958),
.B(n_6892),
.Y(n_7189)
);

HB1xp67_ASAP7_75t_L g7190 ( 
.A(n_6944),
.Y(n_7190)
);

INVx4_ASAP7_75t_L g7191 ( 
.A(n_6944),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_7017),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_7025),
.Y(n_7193)
);

OAI321xp33_ASAP7_75t_L g7194 ( 
.A1(n_7011),
.A2(n_6792),
.A3(n_6798),
.B1(n_6804),
.B2(n_6805),
.C(n_6935),
.Y(n_7194)
);

INVx3_ASAP7_75t_SL g7195 ( 
.A(n_6977),
.Y(n_7195)
);

NAND2xp5_ASAP7_75t_L g7196 ( 
.A(n_7070),
.B(n_6908),
.Y(n_7196)
);

INVx2_ASAP7_75t_L g7197 ( 
.A(n_6992),
.Y(n_7197)
);

INVx2_ASAP7_75t_SL g7198 ( 
.A(n_7031),
.Y(n_7198)
);

NOR2xp67_ASAP7_75t_L g7199 ( 
.A(n_7031),
.B(n_6902),
.Y(n_7199)
);

OR2x2_ASAP7_75t_L g7200 ( 
.A(n_7052),
.B(n_6954),
.Y(n_7200)
);

AND2x2_ASAP7_75t_L g7201 ( 
.A(n_6980),
.B(n_6908),
.Y(n_7201)
);

AND2x2_ASAP7_75t_L g7202 ( 
.A(n_6976),
.B(n_6912),
.Y(n_7202)
);

INVx1_ASAP7_75t_L g7203 ( 
.A(n_7028),
.Y(n_7203)
);

INVx1_ASAP7_75t_L g7204 ( 
.A(n_7029),
.Y(n_7204)
);

INVx1_ASAP7_75t_L g7205 ( 
.A(n_7034),
.Y(n_7205)
);

OR2x2_ASAP7_75t_L g7206 ( 
.A(n_7020),
.B(n_6930),
.Y(n_7206)
);

NAND2xp5_ASAP7_75t_L g7207 ( 
.A(n_7070),
.B(n_6912),
.Y(n_7207)
);

OR2x2_ASAP7_75t_L g7208 ( 
.A(n_6989),
.B(n_521),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_7049),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_6961),
.B(n_524),
.Y(n_7210)
);

NOR3x1_ASAP7_75t_L g7211 ( 
.A(n_6970),
.B(n_526),
.C(n_527),
.Y(n_7211)
);

AND2x4_ASAP7_75t_SL g7212 ( 
.A(n_7037),
.B(n_527),
.Y(n_7212)
);

NOR3xp33_ASAP7_75t_L g7213 ( 
.A(n_7065),
.B(n_528),
.C(n_529),
.Y(n_7213)
);

INVx1_ASAP7_75t_L g7214 ( 
.A(n_7051),
.Y(n_7214)
);

OR2x2_ASAP7_75t_L g7215 ( 
.A(n_6994),
.B(n_7042),
.Y(n_7215)
);

NOR2xp33_ASAP7_75t_L g7216 ( 
.A(n_6962),
.B(n_529),
.Y(n_7216)
);

AND2x4_ASAP7_75t_L g7217 ( 
.A(n_7053),
.B(n_531),
.Y(n_7217)
);

OR2x2_ASAP7_75t_L g7218 ( 
.A(n_7005),
.B(n_532),
.Y(n_7218)
);

AND2x4_ASAP7_75t_SL g7219 ( 
.A(n_7061),
.B(n_532),
.Y(n_7219)
);

INVx2_ASAP7_75t_L g7220 ( 
.A(n_6956),
.Y(n_7220)
);

AND2x2_ASAP7_75t_L g7221 ( 
.A(n_7087),
.B(n_7094),
.Y(n_7221)
);

NOR3xp33_ASAP7_75t_L g7222 ( 
.A(n_7110),
.B(n_6942),
.C(n_6967),
.Y(n_7222)
);

AND2x2_ASAP7_75t_L g7223 ( 
.A(n_7180),
.B(n_7002),
.Y(n_7223)
);

INVx3_ASAP7_75t_L g7224 ( 
.A(n_7191),
.Y(n_7224)
);

INVx1_ASAP7_75t_L g7225 ( 
.A(n_7190),
.Y(n_7225)
);

INVx1_ASAP7_75t_L g7226 ( 
.A(n_7218),
.Y(n_7226)
);

AND2x2_ASAP7_75t_L g7227 ( 
.A(n_7195),
.B(n_7072),
.Y(n_7227)
);

AND3x2_ASAP7_75t_L g7228 ( 
.A(n_7120),
.B(n_7039),
.C(n_6982),
.Y(n_7228)
);

NAND2xp33_ASAP7_75t_SL g7229 ( 
.A(n_7191),
.B(n_7074),
.Y(n_7229)
);

NAND2xp5_ASAP7_75t_L g7230 ( 
.A(n_7111),
.B(n_6982),
.Y(n_7230)
);

AND2x2_ASAP7_75t_SL g7231 ( 
.A(n_7173),
.B(n_6985),
.Y(n_7231)
);

OR2x2_ASAP7_75t_L g7232 ( 
.A(n_7140),
.B(n_6991),
.Y(n_7232)
);

INVx2_ASAP7_75t_SL g7233 ( 
.A(n_7119),
.Y(n_7233)
);

NAND3xp33_ASAP7_75t_SL g7234 ( 
.A(n_7181),
.B(n_6999),
.C(n_7023),
.Y(n_7234)
);

AOI31xp33_ASAP7_75t_L g7235 ( 
.A1(n_7100),
.A2(n_7172),
.A3(n_7085),
.B(n_7084),
.Y(n_7235)
);

OR2x2_ASAP7_75t_L g7236 ( 
.A(n_7102),
.B(n_7057),
.Y(n_7236)
);

AO221x1_ASAP7_75t_L g7237 ( 
.A1(n_7161),
.A2(n_6942),
.B1(n_6990),
.B2(n_7066),
.C(n_6956),
.Y(n_7237)
);

INVx1_ASAP7_75t_L g7238 ( 
.A(n_7096),
.Y(n_7238)
);

AND2x2_ASAP7_75t_L g7239 ( 
.A(n_7092),
.B(n_7119),
.Y(n_7239)
);

NAND2xp5_ASAP7_75t_L g7240 ( 
.A(n_7166),
.B(n_7043),
.Y(n_7240)
);

AND2x2_ASAP7_75t_L g7241 ( 
.A(n_7121),
.B(n_6997),
.Y(n_7241)
);

OR2x2_ASAP7_75t_L g7242 ( 
.A(n_7103),
.B(n_7000),
.Y(n_7242)
);

INVx2_ASAP7_75t_L g7243 ( 
.A(n_7169),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_7167),
.Y(n_7244)
);

INVx2_ASAP7_75t_L g7245 ( 
.A(n_7202),
.Y(n_7245)
);

AND2x4_ASAP7_75t_L g7246 ( 
.A(n_7112),
.B(n_7099),
.Y(n_7246)
);

NAND2xp5_ASAP7_75t_L g7247 ( 
.A(n_7164),
.B(n_7040),
.Y(n_7247)
);

AND2x2_ASAP7_75t_L g7248 ( 
.A(n_7157),
.B(n_7000),
.Y(n_7248)
);

OAI222xp33_ASAP7_75t_L g7249 ( 
.A1(n_7171),
.A2(n_536),
.B1(n_537),
.B2(n_540),
.C1(n_541),
.C2(n_542),
.Y(n_7249)
);

AO21x2_ASAP7_75t_L g7250 ( 
.A1(n_7154),
.A2(n_536),
.B(n_540),
.Y(n_7250)
);

AND2x2_ASAP7_75t_L g7251 ( 
.A(n_7156),
.B(n_541),
.Y(n_7251)
);

AND2x4_ASAP7_75t_L g7252 ( 
.A(n_7112),
.B(n_543),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_7208),
.Y(n_7253)
);

AND2x2_ASAP7_75t_L g7254 ( 
.A(n_7152),
.B(n_544),
.Y(n_7254)
);

NAND2xp5_ASAP7_75t_L g7255 ( 
.A(n_7177),
.B(n_544),
.Y(n_7255)
);

NAND2xp5_ASAP7_75t_L g7256 ( 
.A(n_7217),
.B(n_7201),
.Y(n_7256)
);

NAND2xp5_ASAP7_75t_SL g7257 ( 
.A(n_7141),
.B(n_2240),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_7095),
.Y(n_7258)
);

OR2x2_ASAP7_75t_L g7259 ( 
.A(n_7086),
.B(n_545),
.Y(n_7259)
);

NAND2xp5_ASAP7_75t_L g7260 ( 
.A(n_7138),
.B(n_545),
.Y(n_7260)
);

NAND2xp5_ASAP7_75t_L g7261 ( 
.A(n_7175),
.B(n_547),
.Y(n_7261)
);

CKINVDCx20_ASAP7_75t_R g7262 ( 
.A(n_7144),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_7215),
.Y(n_7263)
);

INVx2_ASAP7_75t_L g7264 ( 
.A(n_7182),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_7084),
.Y(n_7265)
);

AND2x2_ASAP7_75t_L g7266 ( 
.A(n_7130),
.B(n_548),
.Y(n_7266)
);

AND2x2_ASAP7_75t_L g7267 ( 
.A(n_7130),
.B(n_548),
.Y(n_7267)
);

AND2x2_ASAP7_75t_L g7268 ( 
.A(n_7097),
.B(n_549),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_7085),
.Y(n_7269)
);

HB1xp67_ASAP7_75t_L g7270 ( 
.A(n_7199),
.Y(n_7270)
);

INVx1_ASAP7_75t_L g7271 ( 
.A(n_7088),
.Y(n_7271)
);

NOR2xp33_ASAP7_75t_L g7272 ( 
.A(n_7175),
.B(n_549),
.Y(n_7272)
);

INVx1_ASAP7_75t_L g7273 ( 
.A(n_7088),
.Y(n_7273)
);

INVx1_ASAP7_75t_SL g7274 ( 
.A(n_7122),
.Y(n_7274)
);

NAND4xp25_ASAP7_75t_L g7275 ( 
.A(n_7176),
.B(n_555),
.C(n_552),
.D(n_554),
.Y(n_7275)
);

INVx2_ASAP7_75t_L g7276 ( 
.A(n_7132),
.Y(n_7276)
);

AND2x4_ASAP7_75t_SL g7277 ( 
.A(n_7139),
.B(n_552),
.Y(n_7277)
);

AND2x2_ASAP7_75t_SL g7278 ( 
.A(n_7211),
.B(n_554),
.Y(n_7278)
);

INVx2_ASAP7_75t_L g7279 ( 
.A(n_7137),
.Y(n_7279)
);

NAND4xp25_ASAP7_75t_SL g7280 ( 
.A(n_7176),
.B(n_558),
.C(n_556),
.D(n_557),
.Y(n_7280)
);

AND2x2_ASAP7_75t_L g7281 ( 
.A(n_7108),
.B(n_556),
.Y(n_7281)
);

OAI31xp33_ASAP7_75t_L g7282 ( 
.A1(n_7125),
.A2(n_7185),
.A3(n_7216),
.B(n_7210),
.Y(n_7282)
);

INVx1_ASAP7_75t_SL g7283 ( 
.A(n_7189),
.Y(n_7283)
);

HB1xp67_ASAP7_75t_L g7284 ( 
.A(n_7083),
.Y(n_7284)
);

NOR2xp33_ASAP7_75t_L g7285 ( 
.A(n_7142),
.B(n_557),
.Y(n_7285)
);

INVx1_ASAP7_75t_SL g7286 ( 
.A(n_7212),
.Y(n_7286)
);

AND2x2_ASAP7_75t_L g7287 ( 
.A(n_7198),
.B(n_7089),
.Y(n_7287)
);

AOI21xp5_ASAP7_75t_L g7288 ( 
.A1(n_7194),
.A2(n_7147),
.B(n_7183),
.Y(n_7288)
);

OAI322xp33_ASAP7_75t_L g7289 ( 
.A1(n_7200),
.A2(n_559),
.A3(n_560),
.B1(n_561),
.B2(n_564),
.C1(n_565),
.C2(n_566),
.Y(n_7289)
);

INVxp67_ASAP7_75t_L g7290 ( 
.A(n_7165),
.Y(n_7290)
);

INVx3_ASAP7_75t_L g7291 ( 
.A(n_7083),
.Y(n_7291)
);

INVx2_ASAP7_75t_L g7292 ( 
.A(n_7137),
.Y(n_7292)
);

INVx1_ASAP7_75t_L g7293 ( 
.A(n_7149),
.Y(n_7293)
);

NAND2xp5_ASAP7_75t_L g7294 ( 
.A(n_7217),
.B(n_560),
.Y(n_7294)
);

NAND3xp33_ASAP7_75t_L g7295 ( 
.A(n_7118),
.B(n_567),
.C(n_569),
.Y(n_7295)
);

AND2x2_ASAP7_75t_L g7296 ( 
.A(n_7091),
.B(n_569),
.Y(n_7296)
);

HB1xp67_ASAP7_75t_L g7297 ( 
.A(n_7150),
.Y(n_7297)
);

OR2x2_ASAP7_75t_L g7298 ( 
.A(n_7197),
.B(n_571),
.Y(n_7298)
);

INVx2_ASAP7_75t_L g7299 ( 
.A(n_7179),
.Y(n_7299)
);

NAND4xp25_ASAP7_75t_L g7300 ( 
.A(n_7098),
.B(n_571),
.C(n_574),
.D(n_575),
.Y(n_7300)
);

AND2x2_ASAP7_75t_L g7301 ( 
.A(n_7124),
.B(n_574),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_7117),
.Y(n_7302)
);

NAND2xp5_ASAP7_75t_L g7303 ( 
.A(n_7155),
.B(n_575),
.Y(n_7303)
);

OA21x2_ASAP7_75t_L g7304 ( 
.A1(n_7105),
.A2(n_577),
.B(n_579),
.Y(n_7304)
);

AND2x2_ASAP7_75t_L g7305 ( 
.A(n_7127),
.B(n_579),
.Y(n_7305)
);

AND2x2_ASAP7_75t_L g7306 ( 
.A(n_7090),
.B(n_581),
.Y(n_7306)
);

NOR2xp33_ASAP7_75t_L g7307 ( 
.A(n_7104),
.B(n_582),
.Y(n_7307)
);

AND2x2_ASAP7_75t_L g7308 ( 
.A(n_7093),
.B(n_582),
.Y(n_7308)
);

NAND2x1p5_ASAP7_75t_L g7309 ( 
.A(n_7131),
.B(n_583),
.Y(n_7309)
);

NAND2xp5_ASAP7_75t_L g7310 ( 
.A(n_7151),
.B(n_584),
.Y(n_7310)
);

NAND2xp5_ASAP7_75t_SL g7311 ( 
.A(n_7134),
.B(n_2242),
.Y(n_7311)
);

NAND2xp5_ASAP7_75t_L g7312 ( 
.A(n_7151),
.B(n_585),
.Y(n_7312)
);

NAND2xp5_ASAP7_75t_L g7313 ( 
.A(n_7159),
.B(n_585),
.Y(n_7313)
);

INVx2_ASAP7_75t_L g7314 ( 
.A(n_7219),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_7116),
.Y(n_7315)
);

AND2x2_ASAP7_75t_L g7316 ( 
.A(n_7131),
.B(n_586),
.Y(n_7316)
);

INVx2_ASAP7_75t_L g7317 ( 
.A(n_7206),
.Y(n_7317)
);

AND2x2_ASAP7_75t_L g7318 ( 
.A(n_7109),
.B(n_587),
.Y(n_7318)
);

OR2x2_ASAP7_75t_L g7319 ( 
.A(n_7101),
.B(n_588),
.Y(n_7319)
);

OR2x2_ASAP7_75t_L g7320 ( 
.A(n_7106),
.B(n_588),
.Y(n_7320)
);

NAND2xp5_ASAP7_75t_L g7321 ( 
.A(n_7123),
.B(n_589),
.Y(n_7321)
);

AND2x2_ASAP7_75t_L g7322 ( 
.A(n_7160),
.B(n_590),
.Y(n_7322)
);

INVx1_ASAP7_75t_L g7323 ( 
.A(n_7126),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_7128),
.Y(n_7324)
);

NAND2xp5_ASAP7_75t_L g7325 ( 
.A(n_7184),
.B(n_591),
.Y(n_7325)
);

AND2x2_ASAP7_75t_L g7326 ( 
.A(n_7162),
.B(n_592),
.Y(n_7326)
);

INVx1_ASAP7_75t_L g7327 ( 
.A(n_7133),
.Y(n_7327)
);

OR2x2_ASAP7_75t_L g7328 ( 
.A(n_7170),
.B(n_592),
.Y(n_7328)
);

NOR3xp33_ASAP7_75t_L g7329 ( 
.A(n_7133),
.B(n_593),
.C(n_594),
.Y(n_7329)
);

AND2x2_ASAP7_75t_L g7330 ( 
.A(n_7186),
.B(n_595),
.Y(n_7330)
);

BUFx3_ASAP7_75t_L g7331 ( 
.A(n_7163),
.Y(n_7331)
);

AND2x2_ASAP7_75t_L g7332 ( 
.A(n_7187),
.B(n_596),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_L g7333 ( 
.A(n_7178),
.B(n_596),
.Y(n_7333)
);

OAI31xp33_ASAP7_75t_SL g7334 ( 
.A1(n_7146),
.A2(n_597),
.A3(n_598),
.B(n_599),
.Y(n_7334)
);

AND2x4_ASAP7_75t_L g7335 ( 
.A(n_7220),
.B(n_597),
.Y(n_7335)
);

INVx2_ASAP7_75t_L g7336 ( 
.A(n_7136),
.Y(n_7336)
);

NAND4xp25_ASAP7_75t_L g7337 ( 
.A(n_7107),
.B(n_598),
.C(n_600),
.D(n_602),
.Y(n_7337)
);

AND2x4_ASAP7_75t_L g7338 ( 
.A(n_7113),
.B(n_603),
.Y(n_7338)
);

AND2x2_ASAP7_75t_L g7339 ( 
.A(n_7129),
.B(n_603),
.Y(n_7339)
);

OR2x2_ASAP7_75t_L g7340 ( 
.A(n_7297),
.B(n_7168),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_7235),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_SL g7342 ( 
.A(n_7262),
.B(n_7196),
.Y(n_7342)
);

OR2x2_ASAP7_75t_L g7343 ( 
.A(n_7232),
.B(n_7135),
.Y(n_7343)
);

INVxp67_ASAP7_75t_L g7344 ( 
.A(n_7284),
.Y(n_7344)
);

NAND2x1_ASAP7_75t_L g7345 ( 
.A(n_7291),
.B(n_7143),
.Y(n_7345)
);

OR2x2_ASAP7_75t_L g7346 ( 
.A(n_7274),
.B(n_7145),
.Y(n_7346)
);

NAND2xp5_ASAP7_75t_L g7347 ( 
.A(n_7221),
.B(n_7136),
.Y(n_7347)
);

NOR2xp33_ASAP7_75t_L g7348 ( 
.A(n_7249),
.B(n_7148),
.Y(n_7348)
);

INVx1_ASAP7_75t_L g7349 ( 
.A(n_7304),
.Y(n_7349)
);

NOR2xp33_ASAP7_75t_L g7350 ( 
.A(n_7286),
.B(n_7207),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_L g7351 ( 
.A(n_7334),
.B(n_7115),
.Y(n_7351)
);

OR2x2_ASAP7_75t_L g7352 ( 
.A(n_7274),
.B(n_7158),
.Y(n_7352)
);

INVx2_ASAP7_75t_L g7353 ( 
.A(n_7309),
.Y(n_7353)
);

OR2x2_ASAP7_75t_L g7354 ( 
.A(n_7235),
.B(n_7188),
.Y(n_7354)
);

NAND4xp25_ASAP7_75t_L g7355 ( 
.A(n_7222),
.B(n_7214),
.C(n_7192),
.D(n_7209),
.Y(n_7355)
);

INVx1_ASAP7_75t_L g7356 ( 
.A(n_7304),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_7263),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_7328),
.Y(n_7358)
);

OR2x2_ASAP7_75t_L g7359 ( 
.A(n_7225),
.B(n_7193),
.Y(n_7359)
);

AOI21xp5_ASAP7_75t_L g7360 ( 
.A1(n_7230),
.A2(n_7114),
.B(n_7213),
.Y(n_7360)
);

AND2x2_ASAP7_75t_L g7361 ( 
.A(n_7239),
.B(n_7203),
.Y(n_7361)
);

AND2x2_ASAP7_75t_L g7362 ( 
.A(n_7227),
.B(n_7204),
.Y(n_7362)
);

INVx2_ASAP7_75t_L g7363 ( 
.A(n_7291),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_7255),
.Y(n_7364)
);

OR2x2_ASAP7_75t_L g7365 ( 
.A(n_7283),
.B(n_7205),
.Y(n_7365)
);

INVx1_ASAP7_75t_L g7366 ( 
.A(n_7319),
.Y(n_7366)
);

AND2x2_ASAP7_75t_L g7367 ( 
.A(n_7223),
.B(n_7153),
.Y(n_7367)
);

NOR2x1_ASAP7_75t_L g7368 ( 
.A(n_7275),
.B(n_7174),
.Y(n_7368)
);

INVxp67_ASAP7_75t_SL g7369 ( 
.A(n_7290),
.Y(n_7369)
);

INVxp67_ASAP7_75t_L g7370 ( 
.A(n_7270),
.Y(n_7370)
);

AND2x4_ASAP7_75t_L g7371 ( 
.A(n_7246),
.B(n_604),
.Y(n_7371)
);

OR2x2_ASAP7_75t_L g7372 ( 
.A(n_7283),
.B(n_605),
.Y(n_7372)
);

AND2x2_ASAP7_75t_L g7373 ( 
.A(n_7246),
.B(n_607),
.Y(n_7373)
);

INVx1_ASAP7_75t_L g7374 ( 
.A(n_7254),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_L g7375 ( 
.A(n_7334),
.B(n_609),
.Y(n_7375)
);

NAND2xp5_ASAP7_75t_L g7376 ( 
.A(n_7252),
.B(n_610),
.Y(n_7376)
);

AND2x2_ASAP7_75t_L g7377 ( 
.A(n_7245),
.B(n_610),
.Y(n_7377)
);

NOR2x1p5_ASAP7_75t_SL g7378 ( 
.A(n_7276),
.B(n_611),
.Y(n_7378)
);

AND2x2_ASAP7_75t_L g7379 ( 
.A(n_7264),
.B(n_7266),
.Y(n_7379)
);

INVx1_ASAP7_75t_SL g7380 ( 
.A(n_7278),
.Y(n_7380)
);

NOR2xp67_ASAP7_75t_L g7381 ( 
.A(n_7224),
.B(n_7233),
.Y(n_7381)
);

OR2x2_ASAP7_75t_L g7382 ( 
.A(n_7275),
.B(n_612),
.Y(n_7382)
);

INVx3_ASAP7_75t_L g7383 ( 
.A(n_7252),
.Y(n_7383)
);

INVx1_ASAP7_75t_L g7384 ( 
.A(n_7230),
.Y(n_7384)
);

INVx1_ASAP7_75t_SL g7385 ( 
.A(n_7277),
.Y(n_7385)
);

AND2x2_ASAP7_75t_L g7386 ( 
.A(n_7267),
.B(n_7224),
.Y(n_7386)
);

OR2x2_ASAP7_75t_L g7387 ( 
.A(n_7244),
.B(n_612),
.Y(n_7387)
);

AND2x4_ASAP7_75t_L g7388 ( 
.A(n_7251),
.B(n_613),
.Y(n_7388)
);

NAND2xp5_ASAP7_75t_L g7389 ( 
.A(n_7228),
.B(n_614),
.Y(n_7389)
);

INVx1_ASAP7_75t_L g7390 ( 
.A(n_7260),
.Y(n_7390)
);

OR2x2_ASAP7_75t_L g7391 ( 
.A(n_7259),
.B(n_7331),
.Y(n_7391)
);

OAI21xp5_ASAP7_75t_L g7392 ( 
.A1(n_7288),
.A2(n_614),
.B(n_615),
.Y(n_7392)
);

OR2x2_ASAP7_75t_L g7393 ( 
.A(n_7242),
.B(n_615),
.Y(n_7393)
);

AND2x2_ASAP7_75t_L g7394 ( 
.A(n_7281),
.B(n_616),
.Y(n_7394)
);

INVx1_ASAP7_75t_SL g7395 ( 
.A(n_7286),
.Y(n_7395)
);

AOI211x1_ASAP7_75t_L g7396 ( 
.A1(n_7295),
.A2(n_617),
.B(n_619),
.C(n_621),
.Y(n_7396)
);

INVx1_ASAP7_75t_L g7397 ( 
.A(n_7320),
.Y(n_7397)
);

BUFx2_ASAP7_75t_L g7398 ( 
.A(n_7229),
.Y(n_7398)
);

AND2x2_ASAP7_75t_L g7399 ( 
.A(n_7287),
.B(n_617),
.Y(n_7399)
);

INVxp67_ASAP7_75t_L g7400 ( 
.A(n_7316),
.Y(n_7400)
);

NAND2xp5_ASAP7_75t_L g7401 ( 
.A(n_7335),
.B(n_622),
.Y(n_7401)
);

INVx1_ASAP7_75t_L g7402 ( 
.A(n_7306),
.Y(n_7402)
);

NAND2xp5_ASAP7_75t_L g7403 ( 
.A(n_7335),
.B(n_623),
.Y(n_7403)
);

AND2x2_ASAP7_75t_L g7404 ( 
.A(n_7296),
.B(n_623),
.Y(n_7404)
);

AND2x2_ASAP7_75t_L g7405 ( 
.A(n_7301),
.B(n_626),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_7308),
.Y(n_7406)
);

XOR2xp5_ASAP7_75t_L g7407 ( 
.A(n_7231),
.B(n_626),
.Y(n_7407)
);

OR2x2_ASAP7_75t_L g7408 ( 
.A(n_7293),
.B(n_627),
.Y(n_7408)
);

NAND2xp5_ASAP7_75t_L g7409 ( 
.A(n_7268),
.B(n_627),
.Y(n_7409)
);

INVx2_ASAP7_75t_L g7410 ( 
.A(n_7338),
.Y(n_7410)
);

INVx1_ASAP7_75t_L g7411 ( 
.A(n_7310),
.Y(n_7411)
);

OR2x2_ASAP7_75t_L g7412 ( 
.A(n_7271),
.B(n_7273),
.Y(n_7412)
);

NOR2xp33_ASAP7_75t_L g7413 ( 
.A(n_7300),
.B(n_628),
.Y(n_7413)
);

INVx2_ASAP7_75t_L g7414 ( 
.A(n_7338),
.Y(n_7414)
);

OAI21xp33_ASAP7_75t_L g7415 ( 
.A1(n_7256),
.A2(n_7248),
.B(n_7243),
.Y(n_7415)
);

INVx1_ASAP7_75t_L g7416 ( 
.A(n_7312),
.Y(n_7416)
);

AND2x4_ASAP7_75t_L g7417 ( 
.A(n_7314),
.B(n_629),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_7318),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_7322),
.Y(n_7419)
);

INVx1_ASAP7_75t_SL g7420 ( 
.A(n_7305),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_7326),
.Y(n_7421)
);

NAND2xp5_ASAP7_75t_L g7422 ( 
.A(n_7237),
.B(n_629),
.Y(n_7422)
);

OAI21xp33_ASAP7_75t_L g7423 ( 
.A1(n_7258),
.A2(n_632),
.B(n_633),
.Y(n_7423)
);

INVx1_ASAP7_75t_SL g7424 ( 
.A(n_7298),
.Y(n_7424)
);

INVx1_ASAP7_75t_L g7425 ( 
.A(n_7260),
.Y(n_7425)
);

HB1xp67_ASAP7_75t_L g7426 ( 
.A(n_7250),
.Y(n_7426)
);

HB1xp67_ASAP7_75t_L g7427 ( 
.A(n_7250),
.Y(n_7427)
);

OR2x2_ASAP7_75t_L g7428 ( 
.A(n_7395),
.B(n_7315),
.Y(n_7428)
);

AND2x2_ASAP7_75t_L g7429 ( 
.A(n_7367),
.B(n_7361),
.Y(n_7429)
);

AND2x2_ASAP7_75t_L g7430 ( 
.A(n_7386),
.B(n_7323),
.Y(n_7430)
);

NAND2xp5_ASAP7_75t_L g7431 ( 
.A(n_7388),
.B(n_7253),
.Y(n_7431)
);

AND2x2_ASAP7_75t_L g7432 ( 
.A(n_7362),
.B(n_7324),
.Y(n_7432)
);

BUFx2_ASAP7_75t_L g7433 ( 
.A(n_7398),
.Y(n_7433)
);

INVx1_ASAP7_75t_L g7434 ( 
.A(n_7426),
.Y(n_7434)
);

INVx1_ASAP7_75t_SL g7435 ( 
.A(n_7354),
.Y(n_7435)
);

NAND2xp5_ASAP7_75t_L g7436 ( 
.A(n_7388),
.B(n_7241),
.Y(n_7436)
);

INVx1_ASAP7_75t_L g7437 ( 
.A(n_7427),
.Y(n_7437)
);

INVx1_ASAP7_75t_SL g7438 ( 
.A(n_7352),
.Y(n_7438)
);

INVx1_ASAP7_75t_L g7439 ( 
.A(n_7349),
.Y(n_7439)
);

INVx2_ASAP7_75t_L g7440 ( 
.A(n_7383),
.Y(n_7440)
);

AND2x2_ASAP7_75t_L g7441 ( 
.A(n_7379),
.B(n_7238),
.Y(n_7441)
);

NOR3xp33_ASAP7_75t_L g7442 ( 
.A(n_7389),
.B(n_7333),
.C(n_7295),
.Y(n_7442)
);

INVx1_ASAP7_75t_L g7443 ( 
.A(n_7356),
.Y(n_7443)
);

NAND2xp5_ASAP7_75t_L g7444 ( 
.A(n_7420),
.B(n_7330),
.Y(n_7444)
);

AND2x2_ASAP7_75t_L g7445 ( 
.A(n_7399),
.B(n_7302),
.Y(n_7445)
);

BUFx2_ASAP7_75t_L g7446 ( 
.A(n_7383),
.Y(n_7446)
);

AND2x2_ASAP7_75t_L g7447 ( 
.A(n_7350),
.B(n_7339),
.Y(n_7447)
);

AND2x2_ASAP7_75t_L g7448 ( 
.A(n_7342),
.B(n_7307),
.Y(n_7448)
);

NOR2xp33_ASAP7_75t_L g7449 ( 
.A(n_7380),
.B(n_7280),
.Y(n_7449)
);

INVx2_ASAP7_75t_L g7450 ( 
.A(n_7371),
.Y(n_7450)
);

HB1xp67_ASAP7_75t_L g7451 ( 
.A(n_7381),
.Y(n_7451)
);

INVx1_ASAP7_75t_SL g7452 ( 
.A(n_7346),
.Y(n_7452)
);

INVx1_ASAP7_75t_SL g7453 ( 
.A(n_7341),
.Y(n_7453)
);

INVx1_ASAP7_75t_SL g7454 ( 
.A(n_7341),
.Y(n_7454)
);

NAND4xp25_ASAP7_75t_L g7455 ( 
.A(n_7355),
.B(n_7282),
.C(n_7333),
.D(n_7269),
.Y(n_7455)
);

INVx1_ASAP7_75t_L g7456 ( 
.A(n_7340),
.Y(n_7456)
);

INVx1_ASAP7_75t_SL g7457 ( 
.A(n_7343),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_7347),
.Y(n_7458)
);

HB1xp67_ASAP7_75t_L g7459 ( 
.A(n_7345),
.Y(n_7459)
);

AND2x2_ASAP7_75t_L g7460 ( 
.A(n_7363),
.B(n_7332),
.Y(n_7460)
);

OAI21xp5_ASAP7_75t_L g7461 ( 
.A1(n_7368),
.A2(n_7272),
.B(n_7261),
.Y(n_7461)
);

INVx2_ASAP7_75t_L g7462 ( 
.A(n_7371),
.Y(n_7462)
);

AND2x2_ASAP7_75t_L g7463 ( 
.A(n_7344),
.B(n_7369),
.Y(n_7463)
);

INVx2_ASAP7_75t_L g7464 ( 
.A(n_7405),
.Y(n_7464)
);

NOR2x1_ASAP7_75t_L g7465 ( 
.A(n_7365),
.B(n_7300),
.Y(n_7465)
);

OR2x2_ASAP7_75t_L g7466 ( 
.A(n_7359),
.B(n_7261),
.Y(n_7466)
);

OR2x2_ASAP7_75t_L g7467 ( 
.A(n_7391),
.B(n_7325),
.Y(n_7467)
);

NAND2xp5_ASAP7_75t_L g7468 ( 
.A(n_7384),
.B(n_7285),
.Y(n_7468)
);

INVx1_ASAP7_75t_L g7469 ( 
.A(n_7375),
.Y(n_7469)
);

INVx1_ASAP7_75t_L g7470 ( 
.A(n_7394),
.Y(n_7470)
);

AOI211x1_ASAP7_75t_L g7471 ( 
.A1(n_7392),
.A2(n_7234),
.B(n_7247),
.C(n_7240),
.Y(n_7471)
);

INVx1_ASAP7_75t_SL g7472 ( 
.A(n_7373),
.Y(n_7472)
);

NOR2xp33_ASAP7_75t_L g7473 ( 
.A(n_7384),
.B(n_7337),
.Y(n_7473)
);

INVx2_ASAP7_75t_SL g7474 ( 
.A(n_7385),
.Y(n_7474)
);

INVxp67_ASAP7_75t_SL g7475 ( 
.A(n_7348),
.Y(n_7475)
);

NAND4xp75_ASAP7_75t_L g7476 ( 
.A(n_7360),
.B(n_7282),
.C(n_7279),
.D(n_7292),
.Y(n_7476)
);

OR2x2_ASAP7_75t_L g7477 ( 
.A(n_7370),
.B(n_7357),
.Y(n_7477)
);

OR2x2_ASAP7_75t_L g7478 ( 
.A(n_7412),
.B(n_7317),
.Y(n_7478)
);

NOR2xp33_ASAP7_75t_L g7479 ( 
.A(n_7410),
.B(n_7337),
.Y(n_7479)
);

INVx2_ASAP7_75t_L g7480 ( 
.A(n_7404),
.Y(n_7480)
);

NAND2xp5_ASAP7_75t_L g7481 ( 
.A(n_7374),
.B(n_7329),
.Y(n_7481)
);

OR2x2_ASAP7_75t_L g7482 ( 
.A(n_7422),
.B(n_7321),
.Y(n_7482)
);

NAND2xp5_ASAP7_75t_L g7483 ( 
.A(n_7396),
.B(n_7226),
.Y(n_7483)
);

INVx1_ASAP7_75t_L g7484 ( 
.A(n_7351),
.Y(n_7484)
);

AND2x2_ASAP7_75t_L g7485 ( 
.A(n_7415),
.B(n_7236),
.Y(n_7485)
);

INVx1_ASAP7_75t_L g7486 ( 
.A(n_7372),
.Y(n_7486)
);

AND2x2_ASAP7_75t_L g7487 ( 
.A(n_7377),
.B(n_7265),
.Y(n_7487)
);

INVx2_ASAP7_75t_L g7488 ( 
.A(n_7417),
.Y(n_7488)
);

NAND2x1p5_ASAP7_75t_L g7489 ( 
.A(n_7417),
.B(n_7336),
.Y(n_7489)
);

AND2x2_ASAP7_75t_L g7490 ( 
.A(n_7353),
.B(n_7327),
.Y(n_7490)
);

INVx1_ASAP7_75t_L g7491 ( 
.A(n_7401),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_7403),
.Y(n_7492)
);

INVx2_ASAP7_75t_L g7493 ( 
.A(n_7414),
.Y(n_7493)
);

NAND2xp5_ASAP7_75t_L g7494 ( 
.A(n_7418),
.B(n_7299),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_7409),
.Y(n_7495)
);

AO22x1_ASAP7_75t_L g7496 ( 
.A1(n_7413),
.A2(n_7303),
.B1(n_7313),
.B2(n_7294),
.Y(n_7496)
);

AND2x2_ASAP7_75t_L g7497 ( 
.A(n_7400),
.B(n_7257),
.Y(n_7497)
);

NAND2xp5_ASAP7_75t_L g7498 ( 
.A(n_7366),
.B(n_7311),
.Y(n_7498)
);

INVxp67_ASAP7_75t_L g7499 ( 
.A(n_7407),
.Y(n_7499)
);

NAND3xp33_ASAP7_75t_L g7500 ( 
.A(n_7393),
.B(n_7289),
.C(n_633),
.Y(n_7500)
);

INVx1_ASAP7_75t_L g7501 ( 
.A(n_7382),
.Y(n_7501)
);

INVx1_ASAP7_75t_L g7502 ( 
.A(n_7408),
.Y(n_7502)
);

INVx1_ASAP7_75t_L g7503 ( 
.A(n_7387),
.Y(n_7503)
);

AOI22xp5_ASAP7_75t_L g7504 ( 
.A1(n_7402),
.A2(n_7289),
.B1(n_635),
.B2(n_636),
.Y(n_7504)
);

AOI222xp33_ASAP7_75t_L g7505 ( 
.A1(n_7434),
.A2(n_7425),
.B1(n_7390),
.B2(n_7378),
.C1(n_7424),
.C2(n_7358),
.Y(n_7505)
);

NAND2xp5_ASAP7_75t_L g7506 ( 
.A(n_7429),
.B(n_7438),
.Y(n_7506)
);

OAI21xp5_ASAP7_75t_L g7507 ( 
.A1(n_7465),
.A2(n_7421),
.B(n_7419),
.Y(n_7507)
);

OAI21xp5_ASAP7_75t_L g7508 ( 
.A1(n_7438),
.A2(n_7397),
.B(n_7406),
.Y(n_7508)
);

INVxp67_ASAP7_75t_SL g7509 ( 
.A(n_7459),
.Y(n_7509)
);

OAI221xp5_ASAP7_75t_L g7510 ( 
.A1(n_7455),
.A2(n_7425),
.B1(n_7390),
.B2(n_7364),
.C(n_7411),
.Y(n_7510)
);

INVx1_ASAP7_75t_SL g7511 ( 
.A(n_7452),
.Y(n_7511)
);

OAI221xp5_ASAP7_75t_L g7512 ( 
.A1(n_7455),
.A2(n_7416),
.B1(n_7423),
.B2(n_7376),
.C(n_637),
.Y(n_7512)
);

INVx2_ASAP7_75t_L g7513 ( 
.A(n_7489),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_7446),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_7436),
.Y(n_7515)
);

OAI31xp33_ASAP7_75t_SL g7516 ( 
.A1(n_7452),
.A2(n_634),
.A3(n_635),
.B(n_636),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_7489),
.Y(n_7517)
);

OR2x2_ASAP7_75t_L g7518 ( 
.A(n_7457),
.B(n_634),
.Y(n_7518)
);

NAND2xp5_ASAP7_75t_L g7519 ( 
.A(n_7472),
.B(n_640),
.Y(n_7519)
);

NAND2xp5_ASAP7_75t_L g7520 ( 
.A(n_7472),
.B(n_640),
.Y(n_7520)
);

AOI21xp33_ASAP7_75t_SL g7521 ( 
.A1(n_7478),
.A2(n_641),
.B(n_642),
.Y(n_7521)
);

NAND3xp33_ASAP7_75t_L g7522 ( 
.A(n_7437),
.B(n_641),
.C(n_643),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7433),
.Y(n_7523)
);

AND2x2_ASAP7_75t_L g7524 ( 
.A(n_7441),
.B(n_645),
.Y(n_7524)
);

AOI32xp33_ASAP7_75t_L g7525 ( 
.A1(n_7435),
.A2(n_645),
.A3(n_646),
.B1(n_647),
.B2(n_648),
.Y(n_7525)
);

INVx1_ASAP7_75t_L g7526 ( 
.A(n_7432),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_7445),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_7430),
.Y(n_7528)
);

AOI21xp33_ASAP7_75t_L g7529 ( 
.A1(n_7449),
.A2(n_647),
.B(n_649),
.Y(n_7529)
);

NAND2xp5_ASAP7_75t_L g7530 ( 
.A(n_7447),
.B(n_650),
.Y(n_7530)
);

INVx1_ASAP7_75t_L g7531 ( 
.A(n_7428),
.Y(n_7531)
);

AOI22xp5_ASAP7_75t_L g7532 ( 
.A1(n_7442),
.A2(n_7469),
.B1(n_7484),
.B2(n_7473),
.Y(n_7532)
);

NAND2xp5_ASAP7_75t_L g7533 ( 
.A(n_7457),
.B(n_652),
.Y(n_7533)
);

NAND2xp5_ASAP7_75t_L g7534 ( 
.A(n_7451),
.B(n_653),
.Y(n_7534)
);

OAI22xp5_ASAP7_75t_L g7535 ( 
.A1(n_7435),
.A2(n_653),
.B1(n_654),
.B2(n_655),
.Y(n_7535)
);

OAI21xp33_ASAP7_75t_L g7536 ( 
.A1(n_7448),
.A2(n_654),
.B(n_657),
.Y(n_7536)
);

NAND2xp5_ASAP7_75t_L g7537 ( 
.A(n_7470),
.B(n_658),
.Y(n_7537)
);

OAI22xp5_ASAP7_75t_L g7538 ( 
.A1(n_7456),
.A2(n_658),
.B1(n_659),
.B2(n_660),
.Y(n_7538)
);

AND2x2_ASAP7_75t_L g7539 ( 
.A(n_7485),
.B(n_659),
.Y(n_7539)
);

O2A1O1Ixp33_ASAP7_75t_L g7540 ( 
.A1(n_7461),
.A2(n_661),
.B(n_662),
.C(n_663),
.Y(n_7540)
);

NOR2xp33_ASAP7_75t_L g7541 ( 
.A(n_7450),
.B(n_661),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7466),
.Y(n_7542)
);

INVx1_ASAP7_75t_L g7543 ( 
.A(n_7488),
.Y(n_7543)
);

OAI21xp33_ASAP7_75t_L g7544 ( 
.A1(n_7463),
.A2(n_662),
.B(n_663),
.Y(n_7544)
);

NAND3xp33_ASAP7_75t_SL g7545 ( 
.A(n_7461),
.B(n_665),
.C(n_666),
.Y(n_7545)
);

OAI21xp5_ASAP7_75t_SL g7546 ( 
.A1(n_7439),
.A2(n_667),
.B(n_668),
.Y(n_7546)
);

INVx2_ASAP7_75t_L g7547 ( 
.A(n_7480),
.Y(n_7547)
);

AND2x2_ASAP7_75t_L g7548 ( 
.A(n_7474),
.B(n_667),
.Y(n_7548)
);

INVx2_ASAP7_75t_L g7549 ( 
.A(n_7464),
.Y(n_7549)
);

AND2x2_ASAP7_75t_L g7550 ( 
.A(n_7487),
.B(n_668),
.Y(n_7550)
);

AOI21xp33_ASAP7_75t_SL g7551 ( 
.A1(n_7444),
.A2(n_669),
.B(n_670),
.Y(n_7551)
);

INVx2_ASAP7_75t_SL g7552 ( 
.A(n_7460),
.Y(n_7552)
);

INVx2_ASAP7_75t_L g7553 ( 
.A(n_7462),
.Y(n_7553)
);

NAND2xp5_ASAP7_75t_L g7554 ( 
.A(n_7475),
.B(n_7440),
.Y(n_7554)
);

OAI21xp5_ASAP7_75t_L g7555 ( 
.A1(n_7476),
.A2(n_670),
.B(n_671),
.Y(n_7555)
);

NAND2xp5_ASAP7_75t_L g7556 ( 
.A(n_7496),
.B(n_671),
.Y(n_7556)
);

INVx1_ASAP7_75t_SL g7557 ( 
.A(n_7467),
.Y(n_7557)
);

INVx1_ASAP7_75t_SL g7558 ( 
.A(n_7431),
.Y(n_7558)
);

OAI21xp5_ASAP7_75t_L g7559 ( 
.A1(n_7500),
.A2(n_672),
.B(n_673),
.Y(n_7559)
);

NAND2xp5_ASAP7_75t_L g7560 ( 
.A(n_7486),
.B(n_7502),
.Y(n_7560)
);

NAND2x1_ASAP7_75t_SL g7561 ( 
.A(n_7490),
.B(n_672),
.Y(n_7561)
);

AND2x2_ASAP7_75t_L g7562 ( 
.A(n_7458),
.B(n_673),
.Y(n_7562)
);

AOI22xp33_ASAP7_75t_L g7563 ( 
.A1(n_7482),
.A2(n_2207),
.B1(n_2086),
.B2(n_2372),
.Y(n_7563)
);

INVx2_ASAP7_75t_L g7564 ( 
.A(n_7493),
.Y(n_7564)
);

NAND2xp5_ASAP7_75t_L g7565 ( 
.A(n_7471),
.B(n_674),
.Y(n_7565)
);

INVxp67_ASAP7_75t_L g7566 ( 
.A(n_7479),
.Y(n_7566)
);

INVx1_ASAP7_75t_L g7567 ( 
.A(n_7468),
.Y(n_7567)
);

AOI22xp5_ASAP7_75t_L g7568 ( 
.A1(n_7501),
.A2(n_676),
.B1(n_677),
.B2(n_679),
.Y(n_7568)
);

NAND3xp33_ASAP7_75t_SL g7569 ( 
.A(n_7505),
.B(n_7453),
.C(n_7454),
.Y(n_7569)
);

INVx1_ASAP7_75t_L g7570 ( 
.A(n_7506),
.Y(n_7570)
);

AND2x2_ASAP7_75t_L g7571 ( 
.A(n_7511),
.B(n_7497),
.Y(n_7571)
);

NOR2xp33_ASAP7_75t_L g7572 ( 
.A(n_7557),
.B(n_7500),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_7561),
.Y(n_7573)
);

AND2x2_ASAP7_75t_L g7574 ( 
.A(n_7548),
.B(n_7453),
.Y(n_7574)
);

NAND2xp5_ASAP7_75t_L g7575 ( 
.A(n_7516),
.B(n_7503),
.Y(n_7575)
);

INVxp67_ASAP7_75t_L g7576 ( 
.A(n_7509),
.Y(n_7576)
);

INVx1_ASAP7_75t_L g7577 ( 
.A(n_7539),
.Y(n_7577)
);

NAND2xp5_ASAP7_75t_L g7578 ( 
.A(n_7524),
.B(n_7495),
.Y(n_7578)
);

NOR2xp33_ASAP7_75t_L g7579 ( 
.A(n_7558),
.B(n_7483),
.Y(n_7579)
);

OR2x2_ASAP7_75t_L g7580 ( 
.A(n_7552),
.B(n_7494),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_7550),
.Y(n_7581)
);

NAND2xp5_ASAP7_75t_L g7582 ( 
.A(n_7521),
.B(n_7504),
.Y(n_7582)
);

NOR3xp33_ASAP7_75t_L g7583 ( 
.A(n_7510),
.B(n_7499),
.C(n_7454),
.Y(n_7583)
);

NAND2xp5_ASAP7_75t_SL g7584 ( 
.A(n_7513),
.B(n_7494),
.Y(n_7584)
);

OR2x2_ASAP7_75t_L g7585 ( 
.A(n_7554),
.B(n_7477),
.Y(n_7585)
);

NAND2xp5_ASAP7_75t_L g7586 ( 
.A(n_7546),
.B(n_7491),
.Y(n_7586)
);

AOI32xp33_ASAP7_75t_L g7587 ( 
.A1(n_7517),
.A2(n_7443),
.A3(n_7481),
.B1(n_7492),
.B2(n_7498),
.Y(n_7587)
);

OAI21xp33_ASAP7_75t_SL g7588 ( 
.A1(n_7523),
.A2(n_7481),
.B(n_679),
.Y(n_7588)
);

AOI21xp33_ASAP7_75t_L g7589 ( 
.A1(n_7565),
.A2(n_7556),
.B(n_7555),
.Y(n_7589)
);

NAND2xp5_ASAP7_75t_L g7590 ( 
.A(n_7546),
.B(n_676),
.Y(n_7590)
);

XNOR2x2_ASAP7_75t_L g7591 ( 
.A(n_7522),
.B(n_681),
.Y(n_7591)
);

NOR2xp33_ASAP7_75t_L g7592 ( 
.A(n_7536),
.B(n_682),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_7564),
.Y(n_7593)
);

NOR2x1_ASAP7_75t_L g7594 ( 
.A(n_7522),
.B(n_682),
.Y(n_7594)
);

AND2x2_ASAP7_75t_L g7595 ( 
.A(n_7528),
.B(n_683),
.Y(n_7595)
);

NOR2xp33_ASAP7_75t_L g7596 ( 
.A(n_7536),
.B(n_7544),
.Y(n_7596)
);

INVx1_ASAP7_75t_L g7597 ( 
.A(n_7514),
.Y(n_7597)
);

AOI32xp33_ASAP7_75t_L g7598 ( 
.A1(n_7531),
.A2(n_683),
.A3(n_685),
.B1(n_686),
.B2(n_687),
.Y(n_7598)
);

AND2x4_ASAP7_75t_L g7599 ( 
.A(n_7508),
.B(n_7547),
.Y(n_7599)
);

AND2x4_ASAP7_75t_L g7600 ( 
.A(n_7549),
.B(n_688),
.Y(n_7600)
);

AND2x2_ASAP7_75t_L g7601 ( 
.A(n_7527),
.B(n_688),
.Y(n_7601)
);

AND2x2_ASAP7_75t_L g7602 ( 
.A(n_7526),
.B(n_7542),
.Y(n_7602)
);

NOR2xp33_ASAP7_75t_SL g7603 ( 
.A(n_7544),
.B(n_689),
.Y(n_7603)
);

AND2x2_ASAP7_75t_L g7604 ( 
.A(n_7507),
.B(n_7515),
.Y(n_7604)
);

AND2x2_ASAP7_75t_L g7605 ( 
.A(n_7532),
.B(n_7567),
.Y(n_7605)
);

NAND2x1p5_ASAP7_75t_L g7606 ( 
.A(n_7518),
.B(n_689),
.Y(n_7606)
);

NAND4xp25_ASAP7_75t_L g7607 ( 
.A(n_7560),
.B(n_690),
.C(n_692),
.D(n_693),
.Y(n_7607)
);

INVx2_ASAP7_75t_L g7608 ( 
.A(n_7562),
.Y(n_7608)
);

INVx1_ASAP7_75t_L g7609 ( 
.A(n_7530),
.Y(n_7609)
);

O2A1O1Ixp33_ASAP7_75t_L g7610 ( 
.A1(n_7559),
.A2(n_692),
.B(n_694),
.C(n_695),
.Y(n_7610)
);

INVx1_ASAP7_75t_L g7611 ( 
.A(n_7553),
.Y(n_7611)
);

AND2x2_ASAP7_75t_L g7612 ( 
.A(n_7534),
.B(n_694),
.Y(n_7612)
);

INVxp67_ASAP7_75t_SL g7613 ( 
.A(n_7533),
.Y(n_7613)
);

INVx1_ASAP7_75t_L g7614 ( 
.A(n_7519),
.Y(n_7614)
);

INVx1_ASAP7_75t_L g7615 ( 
.A(n_7520),
.Y(n_7615)
);

OR2x2_ASAP7_75t_L g7616 ( 
.A(n_7545),
.B(n_696),
.Y(n_7616)
);

NAND2xp5_ASAP7_75t_L g7617 ( 
.A(n_7599),
.B(n_7551),
.Y(n_7617)
);

HB1xp67_ASAP7_75t_L g7618 ( 
.A(n_7599),
.Y(n_7618)
);

NAND2xp5_ASAP7_75t_L g7619 ( 
.A(n_7600),
.B(n_7525),
.Y(n_7619)
);

NAND2xp5_ASAP7_75t_L g7620 ( 
.A(n_7600),
.B(n_7541),
.Y(n_7620)
);

NAND2xp33_ASAP7_75t_SL g7621 ( 
.A(n_7580),
.B(n_7535),
.Y(n_7621)
);

INVx2_ASAP7_75t_L g7622 ( 
.A(n_7606),
.Y(n_7622)
);

NAND2xp5_ASAP7_75t_L g7623 ( 
.A(n_7574),
.B(n_7543),
.Y(n_7623)
);

OAI221xp5_ASAP7_75t_L g7624 ( 
.A1(n_7579),
.A2(n_7512),
.B1(n_7566),
.B2(n_7537),
.C(n_7540),
.Y(n_7624)
);

OAI221xp5_ASAP7_75t_L g7625 ( 
.A1(n_7572),
.A2(n_7568),
.B1(n_7529),
.B2(n_7563),
.C(n_7538),
.Y(n_7625)
);

NOR2xp33_ASAP7_75t_L g7626 ( 
.A(n_7588),
.B(n_698),
.Y(n_7626)
);

OAI322xp33_ASAP7_75t_L g7627 ( 
.A1(n_7576),
.A2(n_698),
.A3(n_700),
.B1(n_701),
.B2(n_702),
.C1(n_703),
.C2(n_705),
.Y(n_7627)
);

NAND2xp5_ASAP7_75t_L g7628 ( 
.A(n_7573),
.B(n_700),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_7571),
.Y(n_7629)
);

INVx2_ASAP7_75t_L g7630 ( 
.A(n_7591),
.Y(n_7630)
);

AOI311xp33_ASAP7_75t_L g7631 ( 
.A1(n_7583),
.A2(n_7597),
.A3(n_7570),
.B(n_7593),
.C(n_7611),
.Y(n_7631)
);

INVxp67_ASAP7_75t_L g7632 ( 
.A(n_7603),
.Y(n_7632)
);

HB1xp67_ASAP7_75t_L g7633 ( 
.A(n_7594),
.Y(n_7633)
);

NAND2xp5_ASAP7_75t_L g7634 ( 
.A(n_7581),
.B(n_701),
.Y(n_7634)
);

INVx1_ASAP7_75t_L g7635 ( 
.A(n_7585),
.Y(n_7635)
);

NAND2xp5_ASAP7_75t_SL g7636 ( 
.A(n_7604),
.B(n_702),
.Y(n_7636)
);

NAND2xp5_ASAP7_75t_SL g7637 ( 
.A(n_7605),
.B(n_705),
.Y(n_7637)
);

NAND2xp5_ASAP7_75t_L g7638 ( 
.A(n_7595),
.B(n_7601),
.Y(n_7638)
);

OR2x2_ASAP7_75t_L g7639 ( 
.A(n_7569),
.B(n_1703),
.Y(n_7639)
);

INVxp67_ASAP7_75t_SL g7640 ( 
.A(n_7575),
.Y(n_7640)
);

OR2x2_ASAP7_75t_L g7641 ( 
.A(n_7584),
.B(n_1703),
.Y(n_7641)
);

NAND2xp5_ASAP7_75t_L g7642 ( 
.A(n_7577),
.B(n_1703),
.Y(n_7642)
);

OAI21xp5_ASAP7_75t_L g7643 ( 
.A1(n_7602),
.A2(n_2184),
.B(n_2685),
.Y(n_7643)
);

NAND2xp5_ASAP7_75t_L g7644 ( 
.A(n_7598),
.B(n_1703),
.Y(n_7644)
);

AOI32xp33_ASAP7_75t_L g7645 ( 
.A1(n_7596),
.A2(n_2618),
.A3(n_2685),
.B1(n_2663),
.B2(n_2639),
.Y(n_7645)
);

INVx1_ASAP7_75t_L g7646 ( 
.A(n_7578),
.Y(n_7646)
);

INVx1_ASAP7_75t_L g7647 ( 
.A(n_7590),
.Y(n_7647)
);

OR2x2_ASAP7_75t_L g7648 ( 
.A(n_7618),
.B(n_7586),
.Y(n_7648)
);

NOR3xp33_ASAP7_75t_L g7649 ( 
.A(n_7640),
.B(n_7613),
.C(n_7587),
.Y(n_7649)
);

INVx2_ASAP7_75t_L g7650 ( 
.A(n_7635),
.Y(n_7650)
);

AOI22xp5_ASAP7_75t_L g7651 ( 
.A1(n_7626),
.A2(n_7592),
.B1(n_7615),
.B2(n_7614),
.Y(n_7651)
);

XNOR2x1_ASAP7_75t_L g7652 ( 
.A(n_7630),
.B(n_7616),
.Y(n_7652)
);

NAND2xp5_ASAP7_75t_L g7653 ( 
.A(n_7629),
.B(n_7608),
.Y(n_7653)
);

INVx1_ASAP7_75t_L g7654 ( 
.A(n_7623),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_7633),
.Y(n_7655)
);

XNOR2xp5_ASAP7_75t_L g7656 ( 
.A(n_7638),
.B(n_7607),
.Y(n_7656)
);

AO22x1_ASAP7_75t_L g7657 ( 
.A1(n_7646),
.A2(n_7617),
.B1(n_7612),
.B2(n_7628),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7619),
.Y(n_7658)
);

OAI211xp5_ASAP7_75t_L g7659 ( 
.A1(n_7631),
.A2(n_7587),
.B(n_7598),
.C(n_7589),
.Y(n_7659)
);

INVxp67_ASAP7_75t_L g7660 ( 
.A(n_7621),
.Y(n_7660)
);

NOR2xp33_ASAP7_75t_L g7661 ( 
.A(n_7622),
.B(n_7637),
.Y(n_7661)
);

NAND2xp5_ASAP7_75t_SL g7662 ( 
.A(n_7632),
.B(n_7610),
.Y(n_7662)
);

NAND2xp5_ASAP7_75t_L g7663 ( 
.A(n_7636),
.B(n_7609),
.Y(n_7663)
);

INVx1_ASAP7_75t_L g7664 ( 
.A(n_7620),
.Y(n_7664)
);

INVxp67_ASAP7_75t_L g7665 ( 
.A(n_7634),
.Y(n_7665)
);

INVx1_ASAP7_75t_L g7666 ( 
.A(n_7641),
.Y(n_7666)
);

OAI22xp5_ASAP7_75t_SL g7667 ( 
.A1(n_7624),
.A2(n_7625),
.B1(n_7582),
.B2(n_7647),
.Y(n_7667)
);

AOI21xp33_ASAP7_75t_L g7668 ( 
.A1(n_7644),
.A2(n_2242),
.B(n_2248),
.Y(n_7668)
);

OAI21xp5_ASAP7_75t_L g7669 ( 
.A1(n_7639),
.A2(n_2618),
.B(n_2685),
.Y(n_7669)
);

OAI31xp33_ASAP7_75t_L g7670 ( 
.A1(n_7642),
.A2(n_1851),
.A3(n_1901),
.B(n_1846),
.Y(n_7670)
);

INVx1_ASAP7_75t_L g7671 ( 
.A(n_7627),
.Y(n_7671)
);

XOR2xp5_ASAP7_75t_L g7672 ( 
.A(n_7643),
.B(n_1703),
.Y(n_7672)
);

AOI322xp5_ASAP7_75t_L g7673 ( 
.A1(n_7643),
.A2(n_1888),
.A3(n_1896),
.B1(n_2758),
.B2(n_2605),
.C1(n_2359),
.C2(n_2304),
.Y(n_7673)
);

INVx1_ASAP7_75t_L g7674 ( 
.A(n_7645),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_7618),
.Y(n_7675)
);

NOR3x1_ASAP7_75t_L g7676 ( 
.A(n_7659),
.B(n_7653),
.C(n_7655),
.Y(n_7676)
);

AOI22xp33_ASAP7_75t_L g7677 ( 
.A1(n_7675),
.A2(n_2086),
.B1(n_2207),
.B2(n_2386),
.Y(n_7677)
);

XNOR2x1_ASAP7_75t_SL g7678 ( 
.A(n_7652),
.B(n_1888),
.Y(n_7678)
);

NAND4xp75_ASAP7_75t_L g7679 ( 
.A(n_7651),
.B(n_2184),
.C(n_2207),
.D(n_2086),
.Y(n_7679)
);

AOI22xp33_ASAP7_75t_L g7680 ( 
.A1(n_7665),
.A2(n_2207),
.B1(n_2386),
.B2(n_2372),
.Y(n_7680)
);

INVxp33_ASAP7_75t_L g7681 ( 
.A(n_7649),
.Y(n_7681)
);

NOR3x1_ASAP7_75t_L g7682 ( 
.A(n_7654),
.B(n_2184),
.C(n_2297),
.Y(n_7682)
);

NOR3xp33_ASAP7_75t_L g7683 ( 
.A(n_7657),
.B(n_1896),
.C(n_1888),
.Y(n_7683)
);

NAND3xp33_ASAP7_75t_L g7684 ( 
.A(n_7648),
.B(n_2242),
.C(n_2248),
.Y(n_7684)
);

NOR2x1_ASAP7_75t_L g7685 ( 
.A(n_7650),
.B(n_2184),
.Y(n_7685)
);

NOR3xp33_ASAP7_75t_L g7686 ( 
.A(n_7660),
.B(n_1896),
.C(n_2685),
.Y(n_7686)
);

NAND4xp75_ASAP7_75t_L g7687 ( 
.A(n_7651),
.B(n_2758),
.C(n_2605),
.D(n_2639),
.Y(n_7687)
);

HB1xp67_ASAP7_75t_L g7688 ( 
.A(n_7656),
.Y(n_7688)
);

NOR2x1p5_ASAP7_75t_L g7689 ( 
.A(n_7671),
.B(n_2242),
.Y(n_7689)
);

NOR3x1_ASAP7_75t_L g7690 ( 
.A(n_7662),
.B(n_2299),
.C(n_2248),
.Y(n_7690)
);

NAND3xp33_ASAP7_75t_SL g7691 ( 
.A(n_7663),
.B(n_2663),
.C(n_2639),
.Y(n_7691)
);

AOI22xp5_ASAP7_75t_L g7692 ( 
.A1(n_7658),
.A2(n_2242),
.B1(n_2360),
.B2(n_2359),
.Y(n_7692)
);

NOR3xp33_ASAP7_75t_L g7693 ( 
.A(n_7667),
.B(n_2663),
.C(n_2639),
.Y(n_7693)
);

AO22x2_ASAP7_75t_SL g7694 ( 
.A1(n_7664),
.A2(n_2294),
.B1(n_2292),
.B2(n_2285),
.Y(n_7694)
);

INVx1_ASAP7_75t_SL g7695 ( 
.A(n_7666),
.Y(n_7695)
);

NOR4xp25_ASAP7_75t_L g7696 ( 
.A(n_7661),
.B(n_7674),
.C(n_7668),
.D(n_7670),
.Y(n_7696)
);

HB1xp67_ASAP7_75t_L g7697 ( 
.A(n_7672),
.Y(n_7697)
);

INVxp67_ASAP7_75t_SL g7698 ( 
.A(n_7669),
.Y(n_7698)
);

XNOR2x1_ASAP7_75t_SL g7699 ( 
.A(n_7673),
.B(n_2248),
.Y(n_7699)
);

NAND4xp25_ASAP7_75t_L g7700 ( 
.A(n_7649),
.B(n_2663),
.C(n_2618),
.D(n_1901),
.Y(n_7700)
);

NOR3xp33_ASAP7_75t_L g7701 ( 
.A(n_7659),
.B(n_2618),
.C(n_1851),
.Y(n_7701)
);

NAND3xp33_ASAP7_75t_L g7702 ( 
.A(n_7649),
.B(n_2758),
.C(n_2605),
.Y(n_7702)
);

OAI211xp5_ASAP7_75t_SL g7703 ( 
.A1(n_7660),
.A2(n_2605),
.B(n_2758),
.C(n_1706),
.Y(n_7703)
);

NOR2xp33_ASAP7_75t_SL g7704 ( 
.A(n_7660),
.B(n_2294),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_7675),
.Y(n_7705)
);

INVxp67_ASAP7_75t_SL g7706 ( 
.A(n_7660),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_7675),
.Y(n_7707)
);

INVxp67_ASAP7_75t_L g7708 ( 
.A(n_7706),
.Y(n_7708)
);

INVx1_ASAP7_75t_L g7709 ( 
.A(n_7705),
.Y(n_7709)
);

OAI21xp5_ASAP7_75t_SL g7710 ( 
.A1(n_7681),
.A2(n_7707),
.B(n_7688),
.Y(n_7710)
);

A2O1A1Ixp33_ASAP7_75t_SL g7711 ( 
.A1(n_7701),
.A2(n_2294),
.B(n_2292),
.C(n_2285),
.Y(n_7711)
);

CKINVDCx20_ASAP7_75t_R g7712 ( 
.A(n_7695),
.Y(n_7712)
);

INVx1_ASAP7_75t_L g7713 ( 
.A(n_7678),
.Y(n_7713)
);

AOI322xp5_ASAP7_75t_L g7714 ( 
.A1(n_7698),
.A2(n_2758),
.A3(n_2605),
.B1(n_2248),
.B2(n_2359),
.C1(n_2285),
.C2(n_2292),
.Y(n_7714)
);

AOI22x1_ASAP7_75t_L g7715 ( 
.A1(n_7689),
.A2(n_2285),
.B1(n_2292),
.B2(n_2294),
.Y(n_7715)
);

AOI222xp33_ASAP7_75t_L g7716 ( 
.A1(n_7691),
.A2(n_2285),
.B1(n_2292),
.B2(n_2294),
.C1(n_2297),
.C2(n_2299),
.Y(n_7716)
);

AOI22xp5_ASAP7_75t_L g7717 ( 
.A1(n_7685),
.A2(n_2297),
.B1(n_2299),
.B2(n_2304),
.Y(n_7717)
);

AND2x2_ASAP7_75t_L g7718 ( 
.A(n_7676),
.B(n_1857),
.Y(n_7718)
);

OAI22xp33_ASAP7_75t_SL g7719 ( 
.A1(n_7704),
.A2(n_2758),
.B1(n_1903),
.B2(n_1870),
.Y(n_7719)
);

INVx1_ASAP7_75t_SL g7720 ( 
.A(n_7687),
.Y(n_7720)
);

NAND3xp33_ASAP7_75t_L g7721 ( 
.A(n_7693),
.B(n_2297),
.C(n_2299),
.Y(n_7721)
);

AOI322xp5_ASAP7_75t_L g7722 ( 
.A1(n_7697),
.A2(n_2297),
.A3(n_2299),
.B1(n_2304),
.B2(n_2335),
.C1(n_2359),
.C2(n_2360),
.Y(n_7722)
);

NOR2xp33_ASAP7_75t_L g7723 ( 
.A(n_7700),
.B(n_2411),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7694),
.Y(n_7724)
);

AND2x4_ASAP7_75t_L g7725 ( 
.A(n_7702),
.B(n_1800),
.Y(n_7725)
);

AOI22xp5_ASAP7_75t_L g7726 ( 
.A1(n_7679),
.A2(n_2360),
.B1(n_2304),
.B2(n_2359),
.Y(n_7726)
);

OA21x2_ASAP7_75t_L g7727 ( 
.A1(n_7684),
.A2(n_2304),
.B(n_2335),
.Y(n_7727)
);

AOI21xp33_ASAP7_75t_SL g7728 ( 
.A1(n_7696),
.A2(n_2335),
.B(n_2360),
.Y(n_7728)
);

INVx1_ASAP7_75t_L g7729 ( 
.A(n_7690),
.Y(n_7729)
);

A2O1A1Ixp33_ASAP7_75t_SL g7730 ( 
.A1(n_7683),
.A2(n_2335),
.B(n_2360),
.C(n_2396),
.Y(n_7730)
);

AOI22xp5_ASAP7_75t_L g7731 ( 
.A1(n_7686),
.A2(n_2335),
.B1(n_2402),
.B2(n_2396),
.Y(n_7731)
);

NAND2x1p5_ASAP7_75t_L g7732 ( 
.A(n_7692),
.B(n_2411),
.Y(n_7732)
);

INVx2_ASAP7_75t_SL g7733 ( 
.A(n_7684),
.Y(n_7733)
);

AOI21xp33_ASAP7_75t_L g7734 ( 
.A1(n_7680),
.A2(n_2411),
.B(n_2372),
.Y(n_7734)
);

OAI21xp5_ASAP7_75t_L g7735 ( 
.A1(n_7703),
.A2(n_1699),
.B(n_1884),
.Y(n_7735)
);

AND3x4_ASAP7_75t_L g7736 ( 
.A(n_7699),
.B(n_2411),
.C(n_2372),
.Y(n_7736)
);

NAND4xp75_ASAP7_75t_L g7737 ( 
.A(n_7682),
.B(n_1783),
.C(n_1706),
.D(n_1875),
.Y(n_7737)
);

OAI21xp5_ASAP7_75t_L g7738 ( 
.A1(n_7677),
.A2(n_1699),
.B(n_1884),
.Y(n_7738)
);

AO221x1_ASAP7_75t_L g7739 ( 
.A1(n_7705),
.A2(n_2411),
.B1(n_2373),
.B2(n_2402),
.C(n_2396),
.Y(n_7739)
);

XNOR2xp5_ASAP7_75t_L g7740 ( 
.A(n_7712),
.B(n_1833),
.Y(n_7740)
);

AOI21xp5_ASAP7_75t_L g7741 ( 
.A1(n_7708),
.A2(n_2402),
.B(n_2396),
.Y(n_7741)
);

BUFx2_ASAP7_75t_L g7742 ( 
.A(n_7709),
.Y(n_7742)
);

NAND2xp5_ASAP7_75t_L g7743 ( 
.A(n_7710),
.B(n_1833),
.Y(n_7743)
);

NAND2x1_ASAP7_75t_L g7744 ( 
.A(n_7729),
.B(n_7713),
.Y(n_7744)
);

AND2x4_ASAP7_75t_L g7745 ( 
.A(n_7720),
.B(n_1833),
.Y(n_7745)
);

NAND2xp5_ASAP7_75t_L g7746 ( 
.A(n_7724),
.B(n_7718),
.Y(n_7746)
);

NOR3xp33_ASAP7_75t_L g7747 ( 
.A(n_7728),
.B(n_1833),
.C(n_1706),
.Y(n_7747)
);

OAI21xp33_ASAP7_75t_L g7748 ( 
.A1(n_7723),
.A2(n_2402),
.B(n_2396),
.Y(n_7748)
);

NOR2x1_ASAP7_75t_L g7749 ( 
.A(n_7738),
.B(n_2402),
.Y(n_7749)
);

AOI211xp5_ASAP7_75t_L g7750 ( 
.A1(n_7719),
.A2(n_2392),
.B(n_2386),
.C(n_2383),
.Y(n_7750)
);

NAND2xp5_ASAP7_75t_L g7751 ( 
.A(n_7739),
.B(n_1815),
.Y(n_7751)
);

NAND5xp2_ASAP7_75t_L g7752 ( 
.A(n_7716),
.B(n_1815),
.C(n_1706),
.D(n_1900),
.E(n_1889),
.Y(n_7752)
);

NOR2xp67_ASAP7_75t_L g7753 ( 
.A(n_7721),
.B(n_1699),
.Y(n_7753)
);

NOR2x1_ASAP7_75t_L g7754 ( 
.A(n_7736),
.B(n_2392),
.Y(n_7754)
);

NOR2x1p5_ASAP7_75t_L g7755 ( 
.A(n_7737),
.B(n_7725),
.Y(n_7755)
);

NAND5xp2_ASAP7_75t_L g7756 ( 
.A(n_7731),
.B(n_1815),
.C(n_1706),
.D(n_1900),
.E(n_1889),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_7733),
.Y(n_7757)
);

NOR3x1_ASAP7_75t_L g7758 ( 
.A(n_7711),
.B(n_1815),
.C(n_1900),
.Y(n_7758)
);

NOR3xp33_ASAP7_75t_L g7759 ( 
.A(n_7735),
.B(n_1815),
.C(n_1900),
.Y(n_7759)
);

AND2x4_ASAP7_75t_L g7760 ( 
.A(n_7717),
.B(n_1833),
.Y(n_7760)
);

AOI211xp5_ASAP7_75t_SL g7761 ( 
.A1(n_7734),
.A2(n_2392),
.B(n_2386),
.C(n_2383),
.Y(n_7761)
);

NOR3x1_ASAP7_75t_L g7762 ( 
.A(n_7730),
.B(n_1814),
.C(n_1900),
.Y(n_7762)
);

NOR3xp33_ASAP7_75t_L g7763 ( 
.A(n_7726),
.B(n_7715),
.C(n_7722),
.Y(n_7763)
);

NOR3xp33_ASAP7_75t_L g7764 ( 
.A(n_7714),
.B(n_1814),
.C(n_1889),
.Y(n_7764)
);

NOR3xp33_ASAP7_75t_L g7765 ( 
.A(n_7732),
.B(n_7727),
.C(n_1814),
.Y(n_7765)
);

NAND2xp5_ASAP7_75t_L g7766 ( 
.A(n_7727),
.B(n_1814),
.Y(n_7766)
);

NOR4xp75_ASAP7_75t_L g7767 ( 
.A(n_7738),
.B(n_1814),
.C(n_1889),
.D(n_1878),
.Y(n_7767)
);

NOR3xp33_ASAP7_75t_L g7768 ( 
.A(n_7710),
.B(n_1889),
.C(n_1878),
.Y(n_7768)
);

AOI211xp5_ASAP7_75t_L g7769 ( 
.A1(n_7757),
.A2(n_2392),
.B(n_2386),
.C(n_2383),
.Y(n_7769)
);

AOI22xp5_ASAP7_75t_L g7770 ( 
.A1(n_7742),
.A2(n_2392),
.B1(n_2383),
.B2(n_2379),
.Y(n_7770)
);

AOI211xp5_ASAP7_75t_L g7771 ( 
.A1(n_7746),
.A2(n_2383),
.B(n_1800),
.C(n_1807),
.Y(n_7771)
);

OAI22xp5_ASAP7_75t_L g7772 ( 
.A1(n_7744),
.A2(n_7740),
.B1(n_7743),
.B2(n_7750),
.Y(n_7772)
);

OAI21xp33_ASAP7_75t_SL g7773 ( 
.A1(n_7754),
.A2(n_1800),
.B(n_1878),
.Y(n_7773)
);

INVx1_ASAP7_75t_SL g7774 ( 
.A(n_7767),
.Y(n_7774)
);

INVx1_ASAP7_75t_L g7775 ( 
.A(n_7751),
.Y(n_7775)
);

NOR2x1p5_ASAP7_75t_L g7776 ( 
.A(n_7766),
.B(n_1800),
.Y(n_7776)
);

NOR2x1_ASAP7_75t_L g7777 ( 
.A(n_7755),
.B(n_1800),
.Y(n_7777)
);

NAND4xp25_ASAP7_75t_L g7778 ( 
.A(n_7762),
.B(n_7752),
.C(n_7758),
.D(n_7761),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7745),
.Y(n_7779)
);

OAI21xp5_ASAP7_75t_SL g7780 ( 
.A1(n_7759),
.A2(n_1878),
.B(n_1875),
.Y(n_7780)
);

NAND4xp75_ASAP7_75t_L g7781 ( 
.A(n_7749),
.B(n_1878),
.C(n_1875),
.D(n_1874),
.Y(n_7781)
);

O2A1O1Ixp33_ASAP7_75t_L g7782 ( 
.A1(n_7768),
.A2(n_1875),
.B(n_1874),
.C(n_1859),
.Y(n_7782)
);

OAI22x1_ASAP7_75t_L g7783 ( 
.A1(n_7745),
.A2(n_7760),
.B1(n_7763),
.B2(n_7753),
.Y(n_7783)
);

NOR2x1_ASAP7_75t_L g7784 ( 
.A(n_7741),
.B(n_1875),
.Y(n_7784)
);

NOR3xp33_ASAP7_75t_L g7785 ( 
.A(n_7748),
.B(n_1787),
.C(n_1874),
.Y(n_7785)
);

NAND4xp25_ASAP7_75t_L g7786 ( 
.A(n_7756),
.B(n_1787),
.C(n_1874),
.D(n_1859),
.Y(n_7786)
);

OAI221xp5_ASAP7_75t_L g7787 ( 
.A1(n_7765),
.A2(n_1787),
.B1(n_1874),
.B2(n_1859),
.C(n_1715),
.Y(n_7787)
);

NAND2xp5_ASAP7_75t_SL g7788 ( 
.A(n_7774),
.B(n_7764),
.Y(n_7788)
);

INVx1_ASAP7_75t_L g7789 ( 
.A(n_7777),
.Y(n_7789)
);

INVx1_ASAP7_75t_L g7790 ( 
.A(n_7776),
.Y(n_7790)
);

INVx2_ASAP7_75t_L g7791 ( 
.A(n_7781),
.Y(n_7791)
);

NOR2x1_ASAP7_75t_SL g7792 ( 
.A(n_7772),
.B(n_7747),
.Y(n_7792)
);

INVx1_ASAP7_75t_L g7793 ( 
.A(n_7778),
.Y(n_7793)
);

NOR3xp33_ASAP7_75t_L g7794 ( 
.A(n_7775),
.B(n_7779),
.C(n_7787),
.Y(n_7794)
);

NOR3xp33_ASAP7_75t_L g7795 ( 
.A(n_7773),
.B(n_7760),
.C(n_1787),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_7783),
.Y(n_7796)
);

AND2x4_ASAP7_75t_L g7797 ( 
.A(n_7770),
.B(n_1787),
.Y(n_7797)
);

NAND2x1p5_ASAP7_75t_L g7798 ( 
.A(n_7784),
.B(n_1783),
.Y(n_7798)
);

NOR3xp33_ASAP7_75t_SL g7799 ( 
.A(n_7780),
.B(n_1783),
.C(n_1859),
.Y(n_7799)
);

AOI22xp5_ASAP7_75t_L g7800 ( 
.A1(n_7786),
.A2(n_1783),
.B1(n_1859),
.B2(n_1857),
.Y(n_7800)
);

NAND3xp33_ASAP7_75t_L g7801 ( 
.A(n_7771),
.B(n_1783),
.C(n_1857),
.Y(n_7801)
);

NAND2xp5_ASAP7_75t_L g7802 ( 
.A(n_7769),
.B(n_1782),
.Y(n_7802)
);

NOR2xp33_ASAP7_75t_R g7803 ( 
.A(n_7785),
.B(n_1782),
.Y(n_7803)
);

NOR3xp33_ASAP7_75t_SL g7804 ( 
.A(n_7782),
.B(n_1782),
.C(n_1857),
.Y(n_7804)
);

NAND5xp2_ASAP7_75t_L g7805 ( 
.A(n_7796),
.B(n_1782),
.C(n_1778),
.D(n_1807),
.E(n_1715),
.Y(n_7805)
);

OAI221xp5_ASAP7_75t_L g7806 ( 
.A1(n_7793),
.A2(n_1782),
.B1(n_1857),
.B2(n_1850),
.C(n_1715),
.Y(n_7806)
);

NAND3xp33_ASAP7_75t_SL g7807 ( 
.A(n_7794),
.B(n_1778),
.C(n_1850),
.Y(n_7807)
);

NAND2xp5_ASAP7_75t_SL g7808 ( 
.A(n_7790),
.B(n_1778),
.Y(n_7808)
);

AO211x2_ASAP7_75t_L g7809 ( 
.A1(n_7789),
.A2(n_1778),
.B(n_1850),
.C(n_1839),
.Y(n_7809)
);

INVx1_ASAP7_75t_L g7810 ( 
.A(n_7798),
.Y(n_7810)
);

NAND5xp2_ASAP7_75t_L g7811 ( 
.A(n_7795),
.B(n_1778),
.C(n_1762),
.D(n_1807),
.E(n_1715),
.Y(n_7811)
);

OAI22xp33_ASAP7_75t_L g7812 ( 
.A1(n_7791),
.A2(n_1850),
.B1(n_1839),
.B2(n_1807),
.Y(n_7812)
);

XNOR2xp5_ASAP7_75t_L g7813 ( 
.A(n_7788),
.B(n_1850),
.Y(n_7813)
);

AOI22xp5_ASAP7_75t_L g7814 ( 
.A1(n_7797),
.A2(n_1839),
.B1(n_1807),
.B2(n_1762),
.Y(n_7814)
);

NAND4xp25_ASAP7_75t_L g7815 ( 
.A(n_7800),
.B(n_1839),
.C(n_1762),
.D(n_1755),
.Y(n_7815)
);

INVx1_ASAP7_75t_L g7816 ( 
.A(n_7792),
.Y(n_7816)
);

O2A1O1Ixp33_ASAP7_75t_L g7817 ( 
.A1(n_7802),
.A2(n_1839),
.B(n_1762),
.C(n_1755),
.Y(n_7817)
);

AND3x1_ASAP7_75t_L g7818 ( 
.A(n_7799),
.B(n_1762),
.C(n_1755),
.Y(n_7818)
);

BUFx2_ASAP7_75t_L g7819 ( 
.A(n_7803),
.Y(n_7819)
);

NOR3xp33_ASAP7_75t_L g7820 ( 
.A(n_7801),
.B(n_1755),
.C(n_1749),
.Y(n_7820)
);

CKINVDCx16_ASAP7_75t_R g7821 ( 
.A(n_7804),
.Y(n_7821)
);

OR3x1_ASAP7_75t_L g7822 ( 
.A(n_7796),
.B(n_1755),
.C(n_1749),
.Y(n_7822)
);

NAND3xp33_ASAP7_75t_SL g7823 ( 
.A(n_7796),
.B(n_1749),
.C(n_1735),
.Y(n_7823)
);

HB1xp67_ASAP7_75t_L g7824 ( 
.A(n_7816),
.Y(n_7824)
);

NAND4xp75_ASAP7_75t_L g7825 ( 
.A(n_7810),
.B(n_1749),
.C(n_1735),
.D(n_1731),
.Y(n_7825)
);

AND2x4_ASAP7_75t_L g7826 ( 
.A(n_7819),
.B(n_1749),
.Y(n_7826)
);

OAI22xp5_ASAP7_75t_SL g7827 ( 
.A1(n_7821),
.A2(n_1735),
.B1(n_1715),
.B2(n_1731),
.Y(n_7827)
);

NAND2xp5_ASAP7_75t_L g7828 ( 
.A(n_7813),
.B(n_7822),
.Y(n_7828)
);

OAI221xp5_ASAP7_75t_SL g7829 ( 
.A1(n_7814),
.A2(n_1735),
.B1(n_1731),
.B2(n_1714),
.C(n_1711),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_7818),
.Y(n_7830)
);

INVx1_ASAP7_75t_L g7831 ( 
.A(n_7805),
.Y(n_7831)
);

NAND2xp5_ASAP7_75t_L g7832 ( 
.A(n_7808),
.B(n_7809),
.Y(n_7832)
);

AOI22xp5_ASAP7_75t_L g7833 ( 
.A1(n_7806),
.A2(n_1735),
.B1(n_1731),
.B2(n_1714),
.Y(n_7833)
);

OAI31xp67_ASAP7_75t_L g7834 ( 
.A1(n_7811),
.A2(n_1731),
.A3(n_1711),
.B(n_1714),
.Y(n_7834)
);

NAND2xp5_ASAP7_75t_L g7835 ( 
.A(n_7820),
.B(n_7817),
.Y(n_7835)
);

AND2x4_ASAP7_75t_L g7836 ( 
.A(n_7807),
.B(n_1699),
.Y(n_7836)
);

OAI22xp5_ASAP7_75t_L g7837 ( 
.A1(n_7812),
.A2(n_1699),
.B1(n_1711),
.B2(n_1714),
.Y(n_7837)
);

OAI221xp5_ASAP7_75t_SL g7838 ( 
.A1(n_7815),
.A2(n_1711),
.B1(n_1714),
.B2(n_1737),
.C(n_1742),
.Y(n_7838)
);

NAND2xp5_ASAP7_75t_L g7839 ( 
.A(n_7823),
.B(n_1711),
.Y(n_7839)
);

NAND2xp5_ASAP7_75t_L g7840 ( 
.A(n_7816),
.B(n_1737),
.Y(n_7840)
);

BUFx2_ASAP7_75t_L g7841 ( 
.A(n_7816),
.Y(n_7841)
);

NOR3xp33_ASAP7_75t_L g7842 ( 
.A(n_7841),
.B(n_1737),
.C(n_1742),
.Y(n_7842)
);

INVx2_ASAP7_75t_SL g7843 ( 
.A(n_7824),
.Y(n_7843)
);

NOR3xp33_ASAP7_75t_L g7844 ( 
.A(n_7840),
.B(n_1737),
.C(n_1742),
.Y(n_7844)
);

INVx1_ASAP7_75t_L g7845 ( 
.A(n_7831),
.Y(n_7845)
);

NOR3xp33_ASAP7_75t_L g7846 ( 
.A(n_7830),
.B(n_1737),
.C(n_1742),
.Y(n_7846)
);

INVx1_ASAP7_75t_L g7847 ( 
.A(n_7828),
.Y(n_7847)
);

OR2x2_ASAP7_75t_L g7848 ( 
.A(n_7832),
.B(n_1742),
.Y(n_7848)
);

HB1xp67_ASAP7_75t_L g7849 ( 
.A(n_7826),
.Y(n_7849)
);

AOI221xp5_ASAP7_75t_L g7850 ( 
.A1(n_7826),
.A2(n_1757),
.B1(n_1764),
.B2(n_1794),
.C(n_1809),
.Y(n_7850)
);

BUFx2_ASAP7_75t_L g7851 ( 
.A(n_7836),
.Y(n_7851)
);

OR2x6_ASAP7_75t_L g7852 ( 
.A(n_7835),
.B(n_1903),
.Y(n_7852)
);

INVx1_ASAP7_75t_L g7853 ( 
.A(n_7839),
.Y(n_7853)
);

INVx1_ASAP7_75t_SL g7854 ( 
.A(n_7843),
.Y(n_7854)
);

INVx1_ASAP7_75t_L g7855 ( 
.A(n_7845),
.Y(n_7855)
);

NAND2xp5_ASAP7_75t_SL g7856 ( 
.A(n_7847),
.B(n_7836),
.Y(n_7856)
);

INVx1_ASAP7_75t_SL g7857 ( 
.A(n_7851),
.Y(n_7857)
);

OAI22xp5_ASAP7_75t_L g7858 ( 
.A1(n_7853),
.A2(n_7848),
.B1(n_7849),
.B2(n_7838),
.Y(n_7858)
);

AO22x2_ASAP7_75t_L g7859 ( 
.A1(n_7844),
.A2(n_7837),
.B1(n_7825),
.B2(n_7834),
.Y(n_7859)
);

XNOR2xp5_ASAP7_75t_L g7860 ( 
.A(n_7852),
.B(n_7842),
.Y(n_7860)
);

OAI22xp5_ASAP7_75t_L g7861 ( 
.A1(n_7854),
.A2(n_7852),
.B1(n_7833),
.B2(n_7829),
.Y(n_7861)
);

INVx1_ASAP7_75t_L g7862 ( 
.A(n_7855),
.Y(n_7862)
);

INVx1_ASAP7_75t_L g7863 ( 
.A(n_7857),
.Y(n_7863)
);

OAI221xp5_ASAP7_75t_L g7864 ( 
.A1(n_7860),
.A2(n_7846),
.B1(n_7850),
.B2(n_7827),
.C(n_1809),
.Y(n_7864)
);

CKINVDCx20_ASAP7_75t_R g7865 ( 
.A(n_7863),
.Y(n_7865)
);

CKINVDCx20_ASAP7_75t_R g7866 ( 
.A(n_7862),
.Y(n_7866)
);

NAND2xp33_ASAP7_75t_SL g7867 ( 
.A(n_7861),
.B(n_7856),
.Y(n_7867)
);

NOR2x1p5_ASAP7_75t_L g7868 ( 
.A(n_7865),
.B(n_7858),
.Y(n_7868)
);

XNOR2xp5_ASAP7_75t_L g7869 ( 
.A(n_7866),
.B(n_7859),
.Y(n_7869)
);

AOI22xp5_ASAP7_75t_L g7870 ( 
.A1(n_7868),
.A2(n_7867),
.B1(n_7864),
.B2(n_1794),
.Y(n_7870)
);

OR2x2_ASAP7_75t_L g7871 ( 
.A(n_7869),
.B(n_1757),
.Y(n_7871)
);

INVx1_ASAP7_75t_L g7872 ( 
.A(n_7871),
.Y(n_7872)
);

AOI22xp33_ASAP7_75t_SL g7873 ( 
.A1(n_7872),
.A2(n_7870),
.B1(n_1764),
.B2(n_1794),
.Y(n_7873)
);

OAI21xp5_ASAP7_75t_L g7874 ( 
.A1(n_7872),
.A2(n_1757),
.B(n_1764),
.Y(n_7874)
);

OAI22xp33_ASAP7_75t_L g7875 ( 
.A1(n_7874),
.A2(n_1757),
.B1(n_1764),
.B2(n_1794),
.Y(n_7875)
);

AOI22xp5_ASAP7_75t_SL g7876 ( 
.A1(n_7873),
.A2(n_1757),
.B1(n_1764),
.B2(n_1794),
.Y(n_7876)
);

AOI221xp5_ASAP7_75t_L g7877 ( 
.A1(n_7875),
.A2(n_1809),
.B1(n_1837),
.B2(n_1845),
.C(n_1869),
.Y(n_7877)
);

OR2x6_ASAP7_75t_L g7878 ( 
.A(n_7876),
.B(n_1870),
.Y(n_7878)
);

AOI221xp5_ASAP7_75t_L g7879 ( 
.A1(n_7877),
.A2(n_1809),
.B1(n_1837),
.B2(n_1845),
.C(n_1869),
.Y(n_7879)
);

AOI211xp5_ASAP7_75t_L g7880 ( 
.A1(n_7879),
.A2(n_7878),
.B(n_1837),
.C(n_1845),
.Y(n_7880)
);


endmodule