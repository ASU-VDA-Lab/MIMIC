module fake_netlist_1_6706_n_21 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_21;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_7;
BUFx6f_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
BUFx2_ASAP7_75t_L g8 ( .A(n_0), .Y(n_8) );
AND2x4_ASAP7_75t_L g9 ( .A(n_1), .B(n_4), .Y(n_9) );
NOR2x1p5_ASAP7_75t_L g10 ( .A(n_3), .B(n_0), .Y(n_10) );
BUFx2_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
INVx4_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_2), .Y(n_13) );
AOI21x1_ASAP7_75t_L g14 ( .A1(n_11), .A2(n_2), .B(n_4), .Y(n_14) );
OAI21x1_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_10), .B(n_12), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_9), .A2(n_12), .B(n_8), .Y(n_16) );
AO31x2_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_12), .A3(n_9), .B(n_7), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NOR2x1_ASAP7_75t_L g19 ( .A(n_18), .B(n_7), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AOI21x1_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_14), .B(n_15), .Y(n_21) );
endmodule