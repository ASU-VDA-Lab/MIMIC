module fake_jpeg_31553_n_380 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_380);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_380;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_10),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_53),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_10),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_55),
.Y(n_72)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_57),
.Y(n_79)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_16),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_65),
.A2(n_78),
.B1(n_89),
.B2(n_94),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_20),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_20),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_39),
.B(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_32),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_22),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_22),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_24),
.C(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_57),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_33),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_32),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_25),
.B1(n_35),
.B2(n_29),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_30),
.B(n_29),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_22),
.Y(n_114)
);

OR2x4_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_30),
.Y(n_96)
);

NOR2x1_ASAP7_75t_R g136 ( 
.A(n_96),
.B(n_81),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_97),
.A2(n_100),
.B(n_129),
.Y(n_156)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_30),
.B(n_28),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_60),
.B1(n_58),
.B2(n_34),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g149 ( 
.A1(n_102),
.A2(n_86),
.B1(n_63),
.B2(n_81),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_32),
.B1(n_35),
.B2(n_20),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_103),
.A2(n_110),
.B1(n_127),
.B2(n_131),
.Y(n_154)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_114),
.Y(n_159)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_17),
.B1(n_34),
.B2(n_28),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx2_ASAP7_75t_SL g164 ( 
.A(n_117),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_122),
.Y(n_135)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_125),
.Y(n_147)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_17),
.B1(n_34),
.B2(n_28),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_26),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_78),
.A2(n_17),
.B1(n_26),
.B2(n_37),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_37),
.B1(n_85),
.B2(n_73),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_33),
.B1(n_26),
.B2(n_37),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_75),
.B1(n_80),
.B2(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_133),
.B(n_85),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_155),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_112),
.A3(n_109),
.B1(n_105),
.B2(n_96),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_146),
.Y(n_187)
);

XOR2x1_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_71),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_141),
.A2(n_33),
.B(n_9),
.C(n_11),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_83),
.C(n_84),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_107),
.C(n_116),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_79),
.A3(n_82),
.B1(n_68),
.B2(n_64),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_165),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_82),
.B1(n_81),
.B2(n_79),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_80),
.B1(n_86),
.B2(n_63),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_161),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_77),
.B(n_68),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_102),
.A2(n_80),
.B1(n_86),
.B2(n_77),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_111),
.B1(n_104),
.B2(n_98),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_74),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_170),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_106),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_171),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_106),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_175),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_197),
.B1(n_164),
.B2(n_134),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_126),
.C(n_122),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_120),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_179),
.B(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_182),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_145),
.B(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_180),
.B(n_188),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_161),
.B(n_160),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g226 ( 
.A(n_181),
.B(n_169),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_113),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_108),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_191),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_140),
.B(n_11),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_99),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_124),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_142),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_9),
.Y(n_227)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_150),
.A2(n_117),
.B1(n_9),
.B2(n_11),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_138),
.B(n_6),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_16),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_154),
.B1(n_149),
.B2(n_152),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_222),
.B1(n_230),
.B2(n_179),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_211),
.B(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_149),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_216),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_225),
.B1(n_229),
.B2(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_154),
.Y(n_216)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_220),
.Y(n_258)
);

AO21x1_ASAP7_75t_SL g221 ( 
.A1(n_181),
.A2(n_156),
.B(n_144),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_184),
.B1(n_191),
.B2(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_12),
.C(n_15),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_228),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_144),
.B1(n_157),
.B2(n_134),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_14),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_151),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_157),
.B1(n_158),
.B2(n_6),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_186),
.A2(n_158),
.B1(n_15),
.B2(n_14),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_175),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_178),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_216),
.A2(n_177),
.B(n_186),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_207),
.B(n_221),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_238),
.Y(n_274)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_212),
.A2(n_170),
.B1(n_186),
.B2(n_174),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_239),
.B(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_252),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_202),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_246),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_247),
.A2(n_248),
.B1(n_255),
.B2(n_256),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_173),
.B1(n_168),
.B2(n_171),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_249),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_185),
.Y(n_250)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_199),
.Y(n_251)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_183),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_253),
.Y(n_280)
);

XOR2x2_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_168),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_203),
.C(n_217),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_226),
.A2(n_171),
.B1(n_190),
.B2(n_189),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_195),
.B1(n_193),
.B2(n_12),
.Y(n_256)
);

BUFx12_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_12),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_207),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_215),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_271),
.C(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_237),
.B(n_214),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_265),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_206),
.B(n_217),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_266),
.A2(n_273),
.B(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_267),
.B(n_239),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_261),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_208),
.C(n_217),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_206),
.C(n_204),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_229),
.B(n_209),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_286),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_233),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_251),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_209),
.C(n_218),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_249),
.C(n_242),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_273),
.A2(n_235),
.B(n_232),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_289),
.B(n_302),
.Y(n_315)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_234),
.B1(n_248),
.B2(n_247),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_293),
.A2(n_297),
.B1(n_299),
.B2(n_308),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_241),
.Y(n_294)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_294),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_235),
.B1(n_245),
.B2(n_252),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_296),
.A2(n_282),
.B1(n_277),
.B2(n_264),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_259),
.B1(n_233),
.B2(n_253),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_240),
.C(n_236),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_218),
.C(n_223),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_274),
.B(n_211),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_200),
.C(n_261),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_285),
.C(n_275),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_268),
.B(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_257),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_267),
.A2(n_261),
.B(n_258),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_270),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_281),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_270),
.B1(n_256),
.B2(n_283),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_314),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_272),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_317),
.C(n_319),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_266),
.C(n_279),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_281),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_286),
.C(n_276),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_324),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_312),
.B1(n_296),
.B2(n_325),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_288),
.C(n_289),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_303),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_327),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_290),
.B(n_309),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_331),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_304),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_330),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_332),
.A2(n_333),
.B1(n_1),
.B2(n_3),
.Y(n_352)
);

AOI221xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_307),
.B1(n_280),
.B2(n_262),
.C(n_277),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_293),
.A3(n_280),
.B1(n_297),
.B2(n_287),
.C1(n_282),
.C2(n_264),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_335),
.B(n_340),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_287),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_338),
.Y(n_344)
);

INVx11_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_324),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_0),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_278),
.B(n_257),
.C(n_258),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_342),
.A2(n_331),
.B(n_334),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_314),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_343),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_332),
.A2(n_311),
.B1(n_220),
.B2(n_219),
.Y(n_347)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_347),
.Y(n_356)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_311),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_351),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_350),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_0),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_354),
.Y(n_357)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_338),
.Y(n_354)
);

AOI21x1_ASAP7_75t_L g359 ( 
.A1(n_344),
.A2(n_330),
.B(n_328),
.Y(n_359)
);

O2A1O1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_359),
.A2(n_5),
.B(n_358),
.C(n_355),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_346),
.A2(n_336),
.B1(n_337),
.B2(n_342),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_362),
.A2(n_349),
.B1(n_343),
.B2(n_5),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_353),
.A2(n_336),
.B(n_4),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_363),
.B(n_364),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_3),
.Y(n_364)
);

NOR2x1p5_ASAP7_75t_L g365 ( 
.A(n_363),
.B(n_354),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_366),
.Y(n_372)
);

NOR2x1_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_347),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_351),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_368),
.B(n_370),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_369),
.A2(n_5),
.B1(n_357),
.B2(n_367),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_356),
.A2(n_5),
.B(n_358),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_372),
.B(n_370),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_373),
.C(n_374),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g380 ( 
.A(n_379),
.B(n_377),
.CI(n_372),
.CON(n_380),
.SN(n_380)
);


endmodule