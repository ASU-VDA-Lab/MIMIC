module fake_jpeg_6293_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_17),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_18),
.B1(n_19),
.B2(n_12),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_13),
.B1(n_18),
.B2(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_37),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_23),
.B(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_10),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_10),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_10),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_22),
.C(n_27),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_34),
.C(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_41),
.CI(n_36),
.CON(n_50),
.SN(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_47),
.C(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_50),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_37),
.B(n_33),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_15),
.B(n_38),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_15),
.C(n_38),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_65),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_48),
.B1(n_53),
.B2(n_50),
.Y(n_64)
);

FAx1_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_58),
.CI(n_15),
.CON(n_67),
.SN(n_67)
);

OAI21x1_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_62),
.B(n_61),
.Y(n_69)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_69),
.C(n_66),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_4),
.C(n_6),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_72),
.B(n_70),
.Y(n_73)
);


endmodule