module real_jpeg_22787_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_0),
.B(n_52),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_0),
.B(n_39),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_0),
.B(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_0),
.B(n_17),
.Y(n_220)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_2),
.B(n_44),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_2),
.B(n_47),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_2),
.B(n_28),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_17),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_2),
.B(n_52),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_2),
.B(n_61),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_4),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_4),
.B(n_47),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_4),
.B(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_5),
.B(n_61),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_7),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_7),
.B(n_52),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_7),
.B(n_28),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_7),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_7),
.B(n_61),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_7),
.B(n_47),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_7),
.B(n_39),
.Y(n_232)
);

INVx8_ASAP7_75t_SL g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_9),
.B(n_61),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_9),
.B(n_28),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_9),
.B(n_47),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_9),
.B(n_39),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_9),
.B(n_44),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_11),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_11),
.B(n_61),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_11),
.B(n_47),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_11),
.B(n_52),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_11),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_11),
.B(n_28),
.Y(n_218)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_13),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_13),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_14),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_14),
.B(n_39),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_14),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_14),
.B(n_34),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_14),
.B(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_14),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_14),
.B(n_28),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_14),
.B(n_52),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_17),
.Y(n_136)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_17),
.Y(n_161)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_17),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_149),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.C(n_55),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_22),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_42),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_23),
.B(n_260),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_24),
.B(n_51),
.C(n_54),
.Y(n_113)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.CI(n_33),
.CON(n_24),
.SN(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_27),
.B(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_32),
.B(n_76),
.Y(n_77)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_32),
.Y(n_181)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_36),
.A2(n_37),
.B(n_38),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_36),
.B(n_42),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.C(n_48),
.Y(n_42)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_43),
.B(n_46),
.CI(n_48),
.CON(n_128),
.SN(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_49),
.B(n_55),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.C(n_65),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_56),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.C(n_60),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_57),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_58),
.B(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_59),
.B(n_60),
.Y(n_249)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_90),
.B2(n_123),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_80),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_78),
.B1(n_82),
.B2(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_82),
.C(n_83),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_84),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_86),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.CI(n_89),
.CON(n_86),
.SN(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_112),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.C(n_108),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_97),
.C(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_98),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_108),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_106),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_122),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_118),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_145),
.C(n_147),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_125),
.A2(n_126),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_141),
.C(n_143),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_127),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.C(n_137),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_128),
.B(n_242),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_128),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_129),
.A2(n_130),
.B1(n_137),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_137),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.C(n_140),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_138),
.B(n_139),
.CI(n_140),
.CON(n_228),
.SN(n_228)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_141),
.B(n_143),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_145),
.B(n_147),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_262),
.C(n_263),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_252),
.C(n_253),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_235),
.C(n_236),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_222),
.C(n_223),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_204),
.C(n_205),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_182),
.C(n_183),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_169),
.C(n_174),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_165),
.B2(n_166),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_167),
.C(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_159),
.Y(n_164)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_164),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_178),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_195),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_188),
.C(n_195),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_194),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_203),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_196),
.Y(n_203)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_199),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_202),
.C(n_203),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_213),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_208),
.C(n_213),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_211),
.C(n_212),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_216),
.C(n_217),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_221),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_230),
.C(n_234),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_228),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_230),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.CI(n_233),
.CON(n_230),
.SN(n_230)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_244),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_240),
.C(n_244),
.Y(n_252)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_248),
.C(n_250),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_247),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_248),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_261),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_258),
.C(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);


endmodule