module fake_jpeg_28533_n_540 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_540);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_53),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_57),
.B(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_90),
.Y(n_163)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_24),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_100),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_24),
.B(n_17),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_97),
.Y(n_126)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_18),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_50),
.A2(n_23),
.B1(n_37),
.B2(n_30),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_30),
.B1(n_37),
.B2(n_27),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_102),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_23),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_44),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_108),
.A2(n_65),
.B1(n_70),
.B2(n_69),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_110),
.B(n_45),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_33),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_112),
.B(n_127),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_32),
.B1(n_41),
.B2(n_46),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_120),
.A2(n_129),
.B1(n_150),
.B2(n_0),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_33),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_78),
.A2(n_32),
.B1(n_28),
.B2(n_27),
.Y(n_129)
);

INVx2_ASAP7_75t_R g130 ( 
.A(n_59),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_130),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_56),
.B(n_28),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_133),
.B(n_137),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_73),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_96),
.B(n_49),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_154),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_100),
.A2(n_46),
.B1(n_44),
.B2(n_41),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_100),
.B(n_49),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_103),
.B(n_47),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_161),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_76),
.A2(n_47),
.B1(n_36),
.B2(n_44),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_61),
.B1(n_68),
.B2(n_67),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_60),
.B(n_46),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_74),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_71),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_79),
.B(n_18),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_165),
.B(n_16),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_169),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_120),
.A2(n_93),
.B1(n_84),
.B2(n_64),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_170),
.A2(n_178),
.B1(n_188),
.B2(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_174),
.B(n_175),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_130),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_155),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_176),
.B(n_200),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_177),
.B(n_185),
.Y(n_270)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

BUFx24_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_126),
.B(n_45),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_139),
.A2(n_71),
.B1(n_62),
.B2(n_60),
.Y(n_188)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_128),
.Y(n_189)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_192),
.Y(n_261)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_46),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_201),
.Y(n_236)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_195),
.Y(n_271)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_197),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_126),
.B(n_54),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_199),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_44),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_135),
.B(n_18),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_210),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_150),
.A2(n_52),
.B1(n_114),
.B2(n_134),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_139),
.A2(n_62),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_207),
.A2(n_227),
.B1(n_0),
.B2(n_2),
.Y(n_259)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_147),
.B(n_111),
.Y(n_210)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_213),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_212),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_15),
.Y(n_213)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_109),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_216),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_15),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_157),
.B(n_12),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_219),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_218),
.A2(n_221),
.B1(n_226),
.B2(n_145),
.Y(n_250)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_222),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_122),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_224),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_132),
.B(n_119),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_225),
.Y(n_269)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_177),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_229),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_116),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_162),
.B(n_119),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_231),
.A2(n_195),
.B(n_199),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_175),
.A2(n_151),
.B(n_121),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_234),
.C(n_215),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_196),
.B(n_104),
.Y(n_234)
);

OAI22x1_ASAP7_75t_L g235 ( 
.A1(n_170),
.A2(n_121),
.B1(n_166),
.B2(n_104),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_235),
.A2(n_189),
.B1(n_173),
.B2(n_168),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_171),
.B(n_136),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_248),
.Y(n_300)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_121),
.A3(n_136),
.B1(n_116),
.B2(n_107),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_254),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_167),
.B(n_107),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_181),
.A2(n_145),
.A3(n_131),
.B1(n_124),
.B2(n_122),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_178),
.A2(n_124),
.B1(n_131),
.B2(n_3),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_255),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_259),
.A2(n_253),
.B1(n_268),
.B2(n_235),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_267),
.A2(n_221),
.B1(n_218),
.B2(n_187),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_206),
.B(n_5),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_276),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_5),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_232),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_280),
.B(n_289),
.Y(n_360)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_282),
.Y(n_355)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_284),
.A2(n_292),
.B1(n_262),
.B2(n_268),
.Y(n_330)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_285),
.Y(n_362)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_252),
.B(n_184),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_297),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_302),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_228),
.B(n_188),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_294),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_270),
.B(n_207),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_241),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_298),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_244),
.A2(n_220),
.B1(n_219),
.B2(n_211),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_243),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_304),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_305),
.A2(n_261),
.B(n_264),
.Y(n_358)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_306),
.Y(n_353)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_256),
.Y(n_307)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_222),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_308),
.Y(n_334)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_245),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_233),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_310),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_229),
.B(n_183),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_311),
.B(n_313),
.Y(n_328)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_312),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_230),
.B(n_169),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_315),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_278),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_317),
.Y(n_359)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_225),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_321),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_319),
.A2(n_320),
.B1(n_325),
.B2(n_327),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_275),
.A2(n_267),
.B1(n_244),
.B2(n_276),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_237),
.B(n_263),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_234),
.B(n_193),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_L g349 ( 
.A1(n_322),
.A2(n_323),
.B(n_249),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_234),
.B(n_192),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_236),
.B(n_5),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_248),
.B(n_239),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_273),
.A2(n_226),
.B1(n_180),
.B2(n_8),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_6),
.C(n_7),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_6),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_356),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_330),
.A2(n_332),
.B1(n_345),
.B2(n_348),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_315),
.A2(n_249),
.B1(n_240),
.B2(n_266),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_284),
.A2(n_247),
.B1(n_268),
.B2(n_255),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_242),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_347),
.C(n_368),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_305),
.B(n_291),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_338),
.A2(n_352),
.B(n_358),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_299),
.A2(n_239),
.B1(n_251),
.B2(n_245),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_296),
.B(n_239),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_301),
.A2(n_261),
.B1(n_266),
.B2(n_269),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_320),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_286),
.A2(n_309),
.B1(n_307),
.B2(n_287),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_350),
.A2(n_286),
.B1(n_302),
.B2(n_334),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_293),
.A2(n_264),
.B(n_277),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_300),
.A2(n_308),
.B(n_301),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_364),
.B(n_288),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_SL g366 ( 
.A1(n_294),
.A2(n_240),
.B(n_271),
.C(n_277),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_366),
.A2(n_306),
.B(n_314),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_271),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_289),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_308),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_371),
.B(n_380),
.C(n_396),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_372),
.B(n_395),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_324),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_354),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_344),
.B(n_290),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_378),
.B(n_388),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_359),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_381),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_326),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_359),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_367),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_382),
.B(n_383),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_367),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_335),
.Y(n_384)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_332),
.A2(n_319),
.B1(n_327),
.B2(n_325),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_385),
.A2(n_339),
.B1(n_336),
.B2(n_333),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_360),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_386),
.B(n_387),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_361),
.A2(n_316),
.B1(n_281),
.B2(n_282),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_346),
.B(n_288),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_355),
.Y(n_389)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_358),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_397),
.Y(n_433)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_295),
.Y(n_394)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_394),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_337),
.B(n_288),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_298),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_398),
.A2(n_366),
.B(n_361),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_347),
.B(n_283),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_399),
.B(n_357),
.Y(n_421)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_351),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_400),
.A2(n_351),
.B1(n_333),
.B2(n_336),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_338),
.B(n_285),
.C(n_312),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_402),
.B(n_364),
.C(n_362),
.Y(n_419)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_403),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_404),
.A2(n_400),
.B1(n_411),
.B2(n_429),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_342),
.Y(n_407)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

AOI31xp33_ASAP7_75t_L g408 ( 
.A1(n_372),
.A2(n_329),
.A3(n_342),
.B(n_366),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_408),
.B(n_432),
.Y(n_442)
);

A2O1A1O1Ixp25_ASAP7_75t_L g412 ( 
.A1(n_391),
.A2(n_342),
.B(n_366),
.C(n_334),
.D(n_352),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_398),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_420),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_393),
.A2(n_339),
.B(n_365),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_429),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_418),
.A2(n_387),
.B1(n_375),
.B2(n_369),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_426),
.C(n_427),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_386),
.B(n_343),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_425),
.Y(n_443)
);

XOR2x2_ASAP7_75t_L g425 ( 
.A(n_371),
.B(n_343),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_365),
.C(n_353),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_353),
.C(n_317),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_392),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_393),
.A2(n_9),
.B(n_10),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_401),
.C(n_376),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_437),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_436),
.A2(n_440),
.B1(n_453),
.B2(n_455),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g437 ( 
.A(n_415),
.B(n_396),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_423),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_438),
.B(n_460),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_416),
.A2(n_390),
.B1(n_377),
.B2(n_375),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_424),
.A2(n_385),
.B1(n_374),
.B2(n_397),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_444),
.A2(n_449),
.B1(n_459),
.B2(n_407),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_447),
.A2(n_432),
.B(n_430),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_422),
.A2(n_374),
.B1(n_382),
.B2(n_383),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_451),
.Y(n_464)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_420),
.Y(n_450)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_450),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_414),
.A2(n_391),
.B1(n_379),
.B2(n_381),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_433),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_410),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_418),
.A2(n_402),
.B1(n_403),
.B2(n_389),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_394),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_457),
.C(n_458),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_413),
.A2(n_10),
.B1(n_384),
.B2(n_406),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_408),
.A2(n_10),
.B1(n_406),
.B2(n_407),
.Y(n_456)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_456),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_10),
.C(n_425),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_419),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_424),
.A2(n_433),
.B1(n_423),
.B2(n_431),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_410),
.B(n_414),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_439),
.A2(n_417),
.B(n_431),
.Y(n_462)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_462),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_455),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_471),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_409),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_467),
.Y(n_489)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_443),
.B(n_434),
.CI(n_412),
.CON(n_471),
.SN(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_444),
.A2(n_434),
.B1(n_405),
.B2(n_421),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_477),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_405),
.C(n_411),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_474),
.C(n_481),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_430),
.C(n_428),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_475),
.B(n_447),
.Y(n_482)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_459),
.Y(n_476)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_476),
.Y(n_496)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_440),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_409),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_480),
.Y(n_495)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_456),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_435),
.C(n_457),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_482),
.B(n_498),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_477),
.A2(n_446),
.B1(n_442),
.B2(n_443),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_483),
.A2(n_472),
.B1(n_463),
.B2(n_480),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_464),
.A2(n_453),
.B(n_436),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_484),
.A2(n_497),
.B(n_478),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_487),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_458),
.C(n_437),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_488),
.A2(n_475),
.B1(n_461),
.B2(n_470),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_469),
.B(n_428),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_490),
.Y(n_506)
);

INVx13_ASAP7_75t_L g493 ( 
.A(n_469),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_467),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_464),
.A2(n_465),
.B(n_476),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_481),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_502),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_491),
.A2(n_478),
.B1(n_470),
.B2(n_461),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_507),
.Y(n_514)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_504),
.B(n_505),
.Y(n_521)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_511),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_491),
.A2(n_473),
.B(n_479),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_509),
.B(n_486),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_488),
.Y(n_511)
);

MAJx2_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_466),
.C(n_471),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_498),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_519),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_506),
.A2(n_496),
.B1(n_493),
.B2(n_484),
.Y(n_518)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_518),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_486),
.C(n_466),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_492),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_L g526 ( 
.A1(n_520),
.A2(n_522),
.B(n_512),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_516),
.A2(n_492),
.B(n_496),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_527),
.C(n_514),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_516),
.A2(n_503),
.B1(n_482),
.B2(n_483),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_471),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_510),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_519),
.A2(n_494),
.B(n_510),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_529),
.Y(n_534)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_530),
.Y(n_533)
);

OAI221xp5_ASAP7_75t_L g531 ( 
.A1(n_528),
.A2(n_521),
.B1(n_513),
.B2(n_523),
.C(n_517),
.Y(n_531)
);

INVx6_ASAP7_75t_L g535 ( 
.A(n_533),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_532),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_535),
.B(n_531),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_534),
.B(n_514),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_494),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_468),
.Y(n_540)
);


endmodule