module fake_jpeg_20845_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_41),
.Y(n_43)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx11_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_48),
.B1(n_50),
.B2(n_37),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_25),
.B1(n_31),
.B2(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_37),
.B1(n_26),
.B2(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_28),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_20),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_38),
.B1(n_54),
.B2(n_53),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_23),
.C(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_36),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_23),
.C(n_30),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_42),
.C(n_36),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_37),
.B1(n_38),
.B2(n_36),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_71),
.B1(n_74),
.B2(n_77),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_39),
.B(n_41),
.C(n_26),
.Y(n_62)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_29),
.B(n_42),
.C(n_12),
.D(n_3),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_64),
.B(n_65),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_17),
.B1(n_24),
.B2(n_19),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_89),
.B(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_55),
.B1(n_46),
.B2(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_36),
.Y(n_70)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_17),
.B1(n_24),
.B2(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_32),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_17),
.B1(n_30),
.B2(n_19),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_47),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_49),
.B1(n_45),
.B2(n_48),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_54),
.B1(n_47),
.B2(n_13),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_30),
.B1(n_22),
.B2(n_29),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_42),
.C(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_42),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_47),
.B1(n_50),
.B2(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_90),
.A2(n_72),
.B1(n_76),
.B2(n_79),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_112),
.B1(n_69),
.B2(n_70),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_100),
.C(n_111),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_102),
.B(n_87),
.Y(n_122)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_68),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_28),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_60),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_47),
.B1(n_35),
.B2(n_46),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_61),
.B1(n_86),
.B2(n_66),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_42),
.C(n_35),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_57),
.C(n_55),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_96),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_65),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_134),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_138),
.B1(n_140),
.B2(n_112),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_130),
.B(n_92),
.Y(n_146)
);

OR2x6_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_87),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_131),
.B1(n_110),
.B2(n_105),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_78),
.B(n_68),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_124),
.A2(n_129),
.B(n_105),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_85),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_63),
.CON(n_128),
.SN(n_128)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_128),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_68),
.B(n_81),
.Y(n_129)
);

NOR2xp67_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_62),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_89),
.B1(n_75),
.B2(n_73),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_142),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_64),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_62),
.B1(n_67),
.B2(n_66),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_79),
.B1(n_76),
.B2(n_55),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_72),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_110),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_46),
.B1(n_57),
.B2(n_29),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_134),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_156),
.B1(n_117),
.B2(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_155),
.B1(n_5),
.B2(n_13),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_149),
.Y(n_176)
);

OAI211xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_92),
.B(n_111),
.C(n_101),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_103),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_114),
.B(n_106),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_95),
.B1(n_115),
.B2(n_106),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_123),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_108),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_8),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_6),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_6),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_15),
.C(n_6),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_123),
.C(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_122),
.A3(n_129),
.B1(n_124),
.B2(n_118),
.C1(n_123),
.C2(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_180),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_123),
.B1(n_141),
.B2(n_136),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_174),
.B1(n_189),
.B2(n_149),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_121),
.B1(n_123),
.B2(n_137),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_157),
.B1(n_153),
.B2(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_183),
.B1(n_143),
.B2(n_150),
.Y(n_201)
);

XOR2x1_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_9),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_186),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_9),
.C(n_14),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_167),
.C(n_146),
.Y(n_190)
);

OAI322xp33_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_5),
.A3(n_12),
.B1(n_11),
.B2(n_3),
.C1(n_4),
.C2(n_15),
.Y(n_187)
);

AOI321xp33_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_163),
.A3(n_165),
.B1(n_11),
.B2(n_4),
.C(n_9),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_145),
.A2(n_144),
.B1(n_156),
.B2(n_166),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_199),
.C(n_200),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_157),
.B1(n_150),
.B2(n_162),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_197),
.B1(n_198),
.B2(n_204),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_164),
.C(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_202),
.C(n_180),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_160),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_195),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_154),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_160),
.B1(n_153),
.B2(n_147),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_161),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_153),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_181),
.C(n_175),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_186),
.C(n_185),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_143),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_200),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_175),
.C(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_215),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_179),
.C(n_171),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_184),
.C(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_184),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_194),
.B1(n_188),
.B2(n_177),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_223),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_208),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_211),
.C(n_209),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_195),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_230),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_188),
.B1(n_203),
.B2(n_196),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_187),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_236),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_225),
.C(n_216),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_224),
.B1(n_221),
.B2(n_203),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_12),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_190),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_241),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_232),
.B1(n_235),
.B2(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_244),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_183),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_247),
.B(n_0),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_236),
.B1(n_1),
.B2(n_2),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_2),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_251),
.C(n_245),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_0),
.C(n_1),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_246),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);


endmodule