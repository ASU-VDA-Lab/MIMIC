module fake_jpeg_1636_n_264 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_82;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_62),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_21),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_52),
.Y(n_124)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_28),
.B(n_2),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_5),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_26),
.B(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_79),
.Y(n_94)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_29),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_81),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_6),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_7),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_29),
.B(n_40),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_37),
.B1(n_20),
.B2(n_30),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_55),
.B1(n_24),
.B2(n_36),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_100),
.B1(n_106),
.B2(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_95),
.B(n_89),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_32),
.B1(n_41),
.B2(n_40),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_30),
.B1(n_36),
.B2(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_113),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_38),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_8),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_122),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_52),
.A2(n_81),
.B1(n_76),
.B2(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_10),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_10),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_139),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_127),
.A2(n_147),
.B1(n_140),
.B2(n_129),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_11),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_129),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_91),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_134),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_24),
.B1(n_19),
.B2(n_38),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_151),
.B1(n_117),
.B2(n_142),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_11),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_19),
.B1(n_38),
.B2(n_106),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_154),
.B1(n_147),
.B2(n_160),
.Y(n_185)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_94),
.A2(n_113),
.A3(n_101),
.B1(n_82),
.B2(n_87),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_108),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_99),
.B1(n_101),
.B2(n_98),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_90),
.B(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_159),
.Y(n_181)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_155),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_100),
.A2(n_92),
.B1(n_96),
.B2(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_108),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_160),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_88),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_158),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_109),
.B(n_97),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_129),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_88),
.B1(n_117),
.B2(n_133),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_166),
.B1(n_173),
.B2(n_183),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_88),
.B1(n_117),
.B2(n_128),
.Y(n_166)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_186),
.B(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_126),
.B1(n_156),
.B2(n_149),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_146),
.C(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_153),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_185),
.B(n_188),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_139),
.A2(n_132),
.B(n_136),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_205),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_170),
.B(n_167),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_180),
.A2(n_150),
.B1(n_137),
.B2(n_136),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_167),
.B1(n_168),
.B2(n_179),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_136),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_181),
.A2(n_165),
.B(n_186),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_175),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_197),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_162),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_173),
.Y(n_199)
);

NOR4xp25_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_188),
.C(n_175),
.D(n_183),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_166),
.B1(n_172),
.B2(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_164),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_194),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_197),
.B1(n_195),
.B2(n_193),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_203),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_222),
.A2(n_170),
.B(n_168),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_190),
.B(n_200),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_224),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_225),
.A2(n_229),
.B1(n_234),
.B2(n_214),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_217),
.A2(n_196),
.B(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_221),
.B(n_192),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_227),
.B(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_191),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_235),
.B1(n_215),
.B2(n_210),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_232),
.C(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_201),
.C(n_202),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_204),
.C(n_207),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_179),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_239),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_229),
.B1(n_230),
.B2(n_234),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_214),
.C(n_211),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_215),
.C(n_225),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_249),
.C(n_237),
.Y(n_251)
);

OA21x2_ASAP7_75t_SL g247 ( 
.A1(n_241),
.A2(n_209),
.B(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_223),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_222),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.C(n_249),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_243),
.B(n_242),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_253),
.A2(n_248),
.B(n_240),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_223),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_256),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_225),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_248),
.C(n_225),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_222),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_218),
.C(n_212),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_260),
.C(n_212),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_262),
.Y(n_264)
);


endmodule