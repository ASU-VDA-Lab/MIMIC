module fake_jpeg_12298_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_48),
.Y(n_57)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_44),
.B1(n_42),
.B2(n_4),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_44),
.B1(n_5),
.B2(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_46),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_63),
.B1(n_67),
.B2(n_16),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_39),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_38),
.B1(n_43),
.B2(n_41),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_71),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_68),
.B(n_9),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_10),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_24),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_12),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_31),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_20),
.B(n_23),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_33),
.B(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_90),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_87),
.B(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_98),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_95),
.B1(n_83),
.B2(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_103),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

AOI21x1_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_99),
.B(n_95),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_93),
.Y(n_108)
);


endmodule