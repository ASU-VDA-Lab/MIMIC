module real_jpeg_8989_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_43;
wire n_54;
wire n_57;
wire n_21;
wire n_37;
wire n_73;
wire n_65;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_69;
wire n_58;
wire n_31;
wire n_67;
wire n_49;
wire n_52;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_44;
wire n_28;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_51;
wire n_47;
wire n_71;
wire n_14;
wire n_45;
wire n_25;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_39;
wire n_36;
wire n_70;
wire n_41;
wire n_26;
wire n_56;
wire n_20;
wire n_32;
wire n_48;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_0),
.A2(n_3),
.B(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_0),
.B(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_0),
.A2(n_6),
.B(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_0),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_2),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_3),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_4),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_5),
.C(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_5),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_6),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_8),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_7),
.B(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_8),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

AOI221xp5_ASAP7_75t_L g27 ( 
.A1(n_9),
.A2(n_20),
.B1(n_28),
.B2(n_31),
.C(n_32),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_9),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_10),
.B(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_10),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_10),
.Y(n_73)
);

AOI211xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_48),
.B(n_59),
.C(n_68),
.Y(n_11)
);

A2O1A1Ixp33_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_26),
.B(n_33),
.C(n_37),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_19),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND4xp25_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_25),
.C(n_35),
.D(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_34),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_42),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_40),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);


endmodule