module fake_netlist_6_2741_n_2432 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2432);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2432;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_437;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_1070;
wire n_458;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_346;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_2398;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_2429;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g238 ( 
.A(n_34),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_46),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_19),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_68),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_119),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_76),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_190),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_46),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_184),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_68),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_51),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_139),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_43),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_132),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_138),
.Y(n_258)
);

BUFx2_ASAP7_75t_SL g259 ( 
.A(n_74),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_20),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_170),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_205),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_82),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_36),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_110),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_67),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_35),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_147),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_79),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_232),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_116),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_159),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_195),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_230),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_183),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_36),
.Y(n_281)
);

BUFx8_ASAP7_75t_SL g282 ( 
.A(n_188),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_120),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_149),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_150),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_122),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_0),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_156),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_8),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_52),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_104),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_109),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_85),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_58),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_178),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_60),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_62),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_16),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_185),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_7),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_113),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_112),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_44),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_165),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_45),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_66),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_151),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_56),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_141),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_21),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_225),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_168),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_63),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_179),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_191),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_29),
.Y(n_318)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_61),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_34),
.Y(n_320)
);

BUFx2_ASAP7_75t_SL g321 ( 
.A(n_92),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_137),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_192),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_61),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_228),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_148),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_96),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_26),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_218),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_103),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_174),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_99),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_71),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_29),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_90),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_136),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_25),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_173),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_172),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_181),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_8),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_227),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_93),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_23),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_219),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_164),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_106),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_20),
.Y(n_348)
);

BUFx10_ASAP7_75t_L g349 ( 
.A(n_64),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_54),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_27),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_18),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_101),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_206),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_52),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_204),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_84),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_214),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_57),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_75),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_180),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_21),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_55),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_10),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_126),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_166),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_131),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_67),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_153),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_77),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_223),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_127),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_23),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_107),
.Y(n_374)
);

BUFx5_ASAP7_75t_L g375 ( 
.A(n_108),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_11),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_58),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_26),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_50),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_121),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_146),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_27),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_182),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_213),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_43),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_48),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_86),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_9),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_51),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_41),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_93),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_32),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_145),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_231),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_54),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_14),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_105),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_197),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_71),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_19),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_69),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_114),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_32),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_87),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_63),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_70),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_217),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_102),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_209),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_193),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_125),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_162),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_41),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_163),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_74),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_31),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_37),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_42),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_79),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_99),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_229),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_7),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_78),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_154),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_78),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_6),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_212),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_140),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_111),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_66),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_135),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_83),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_152),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_28),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_207),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_28),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_91),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_100),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_97),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_92),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_24),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_2),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_48),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_44),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_30),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_0),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_11),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_22),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_31),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_22),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_47),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_144),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_59),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_115),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_220),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_187),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_95),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_87),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_25),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_88),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_216),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_42),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_14),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_3),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_57),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_353),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_282),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_335),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_319),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_289),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_454),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_319),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_329),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_319),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_244),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_319),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_319),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_319),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_242),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_291),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_329),
.B(n_1),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_319),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_319),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_249),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_252),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_242),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_255),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_263),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_319),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_335),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_264),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_274),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_265),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_265),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_258),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_275),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_280),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_265),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_265),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_265),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_283),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_265),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_377),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_258),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_377),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_377),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_377),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_377),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_287),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_377),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_385),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_364),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_292),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_293),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_364),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_364),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_330),
.B(n_1),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_364),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_296),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_451),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_240),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_300),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_240),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_359),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_330),
.B(n_2),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_452),
.B(n_3),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_302),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_452),
.B(n_4),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_451),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_359),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_303),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_463),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_314),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_261),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_375),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_306),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_261),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_278),
.B(n_4),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_R g542 ( 
.A(n_314),
.B(n_371),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_439),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_257),
.B(n_5),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_371),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_413),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_439),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_413),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_257),
.B(n_5),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_309),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_416),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_259),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_311),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_375),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_238),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_326),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_331),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_238),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_239),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_372),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_375),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_417),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_259),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_285),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_336),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_338),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_417),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_372),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_239),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_393),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_243),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_299),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_339),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_243),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_248),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_248),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_262),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_340),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_285),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_354),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_262),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_356),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_260),
.B(n_6),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_294),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_241),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_393),
.B(n_9),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_268),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_268),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_358),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_566),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_493),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_493),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_494),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_536),
.B(n_361),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_537),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_537),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_494),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_469),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_498),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_498),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_540),
.B(n_245),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_558),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_565),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_540),
.B(n_245),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_565),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_568),
.B(n_365),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_469),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_472),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_472),
.B(n_278),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_474),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_499),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_553),
.B(n_245),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_474),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_499),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_583),
.B(n_366),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_480),
.B(n_247),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_526),
.B(n_367),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_500),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_500),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_502),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_476),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_518),
.B(n_394),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_503),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_479),
.B(n_295),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_503),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_505),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_477),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_553),
.B(n_394),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_477),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_554),
.B(n_369),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_554),
.B(n_556),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_505),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_478),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_478),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_506),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_518),
.B(n_411),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_482),
.Y(n_644)
);

OA21x2_ASAP7_75t_L g645 ( 
.A1(n_512),
.A2(n_298),
.B(n_281),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_482),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_490),
.A2(n_307),
.B1(n_418),
.B2(n_376),
.Y(n_647)
);

INVx6_ASAP7_75t_L g648 ( 
.A(n_539),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_506),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_556),
.B(n_374),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_517),
.B(n_409),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_483),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_507),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_525),
.B(n_428),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_508),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_483),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_512),
.B(n_411),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_515),
.B(n_278),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_515),
.B(n_278),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_516),
.B(n_260),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_489),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_489),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_589),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_508),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_510),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_510),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_516),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_539),
.B(n_381),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_521),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_539),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_559),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_521),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_528),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_542),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_545),
.B(n_383),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_523),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_523),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_473),
.B(n_270),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_524),
.B(n_530),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_524),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_530),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_590),
.B(n_250),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_562),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_531),
.Y(n_686)
);

NOR2x1_ASAP7_75t_L g687 ( 
.A(n_593),
.B(n_254),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_562),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_481),
.A2(n_420),
.B1(n_446),
.B2(n_442),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_531),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_533),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_651),
.B(n_475),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_602),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_651),
.B(n_480),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_675),
.B(n_484),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_602),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_675),
.B(n_485),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_602),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_613),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_613),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_612),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_612),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_638),
.B(n_470),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_612),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_612),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_654),
.B(n_511),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_612),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_L g708 ( 
.A(n_647),
.B(n_550),
.C(n_548),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_672),
.B(n_270),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

XOR2xp5_ASAP7_75t_L g711 ( 
.A(n_631),
.B(n_466),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_634),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_599),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_602),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_638),
.B(n_471),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_664),
.B(n_511),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_631),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_677),
.B(n_487),
.Y(n_718)
);

CKINVDCx16_ASAP7_75t_R g719 ( 
.A(n_631),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_634),
.Y(n_720)
);

CKINVDCx6p67_ASAP7_75t_R g721 ( 
.A(n_622),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_599),
.Y(n_722)
);

NAND3xp33_ASAP7_75t_L g723 ( 
.A(n_684),
.B(n_567),
.C(n_555),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_615),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_664),
.B(n_488),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_634),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_676),
.B(n_491),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_634),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_606),
.Y(n_729)
);

XOR2xp5_ASAP7_75t_L g730 ( 
.A(n_647),
.B(n_486),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_615),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_675),
.B(n_492),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_634),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_615),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_675),
.B(n_672),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_615),
.Y(n_736)
);

OAI21xp33_ASAP7_75t_SL g737 ( 
.A1(n_623),
.A2(n_680),
.B(n_622),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_599),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_689),
.A2(n_550),
.B1(n_571),
.B2(n_548),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_618),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_618),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_684),
.A2(n_587),
.B1(n_551),
.B2(n_520),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_638),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_636),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_599),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_676),
.B(n_496),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_614),
.B(n_250),
.Y(n_747)
);

AO22x1_ASAP7_75t_L g748 ( 
.A1(n_680),
.A2(n_425),
.B1(n_298),
.B2(n_301),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_636),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_618),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_676),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_672),
.B(n_497),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_618),
.Y(n_753)
);

XOR2x2_ASAP7_75t_L g754 ( 
.A(n_689),
.B(n_588),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_635),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_620),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_636),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_599),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_687),
.A2(n_501),
.B1(n_513),
.B2(n_509),
.Y(n_759)
);

AND2x6_ASAP7_75t_L g760 ( 
.A(n_606),
.B(n_250),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_687),
.B(n_514),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_635),
.B(n_576),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_677),
.B(n_519),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_613),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_R g765 ( 
.A(n_670),
.B(n_522),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_636),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_L g767 ( 
.A(n_637),
.B(n_546),
.C(n_529),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_648),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_648),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_594),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_598),
.B(n_527),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_672),
.B(n_532),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_598),
.B(n_538),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_594),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_599),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_620),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_611),
.B(n_552),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_636),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_611),
.B(n_557),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_620),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_644),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_680),
.A2(n_534),
.B1(n_468),
.B2(n_301),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_621),
.B(n_560),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_637),
.B(n_569),
.C(n_561),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_672),
.B(n_570),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_621),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_670),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_620),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_623),
.B(n_577),
.Y(n_789)
);

AND2x6_ASAP7_75t_L g790 ( 
.A(n_606),
.B(n_250),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_606),
.A2(n_310),
.B1(n_312),
.B2(n_281),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_613),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_650),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_606),
.A2(n_312),
.B1(n_332),
.B2(n_310),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_644),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_650),
.B(n_582),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_635),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_627),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_609),
.B(n_584),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_627),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_617),
.Y(n_801)
);

AND2x6_ASAP7_75t_L g802 ( 
.A(n_609),
.B(n_661),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_627),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_617),
.B(n_571),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_644),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_644),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_658),
.B(n_533),
.Y(n_807)
);

NOR2x1p5_ASAP7_75t_L g808 ( 
.A(n_669),
.B(n_246),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_648),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_599),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_627),
.Y(n_811)
);

OR2x6_ASAP7_75t_L g812 ( 
.A(n_617),
.B(n_321),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_640),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_640),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_640),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_644),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_658),
.B(n_321),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_609),
.B(n_586),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_648),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_609),
.B(n_495),
.Y(n_820)
);

INVxp33_ASAP7_75t_L g821 ( 
.A(n_681),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_609),
.B(n_384),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_658),
.A2(n_333),
.B1(n_334),
.B2(n_332),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_599),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_648),
.B(n_397),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_648),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_614),
.A2(n_334),
.B1(n_352),
.B2(n_333),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_640),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_604),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_629),
.B(n_402),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_646),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_661),
.B(n_250),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_629),
.B(n_407),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_629),
.A2(n_504),
.B1(n_547),
.B2(n_535),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_669),
.B(n_564),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_614),
.A2(n_378),
.B1(n_386),
.B2(n_352),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_613),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_629),
.A2(n_324),
.B1(n_574),
.B2(n_572),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_646),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_646),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_673),
.B(n_467),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_604),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_673),
.B(n_685),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_691),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_604),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_629),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_646),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_691),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_657),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_613),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_643),
.B(n_247),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_657),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_657),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_692),
.B(n_253),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_713),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_846),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_786),
.B(n_251),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_786),
.B(n_408),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_793),
.B(n_412),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_793),
.B(n_414),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_846),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_693),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_718),
.B(n_613),
.Y(n_863)
);

O2A1O1Ixp5_ASAP7_75t_L g864 ( 
.A1(n_735),
.A2(n_659),
.B(n_660),
.C(n_661),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_755),
.B(n_424),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_693),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_696),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_701),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_771),
.B(n_256),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_777),
.B(n_613),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_807),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_743),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_807),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_804),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_696),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_779),
.B(n_266),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_787),
.B(n_641),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_801),
.B(n_427),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_808),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_737),
.A2(n_660),
.B(n_659),
.C(n_267),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_787),
.B(n_641),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_701),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_713),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_789),
.B(n_269),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_703),
.B(n_645),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_844),
.B(n_641),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_703),
.B(n_645),
.Y(n_887)
);

NAND2xp33_ASAP7_75t_L g888 ( 
.A(n_802),
.B(n_614),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_835),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_801),
.B(n_429),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_844),
.B(n_641),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_848),
.B(n_641),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_848),
.B(n_641),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_802),
.B(n_614),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_797),
.B(n_695),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_710),
.B(n_431),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_698),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_702),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_697),
.B(n_641),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_710),
.B(n_433),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_710),
.B(n_435),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_762),
.B(n_456),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_762),
.B(n_461),
.Y(n_903)
);

NOR2xp67_ASAP7_75t_L g904 ( 
.A(n_784),
.B(n_685),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_732),
.B(n_641),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_698),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_826),
.B(n_652),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_714),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_826),
.B(n_843),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_804),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_802),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_763),
.A2(n_643),
.B1(n_614),
.B2(n_659),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_799),
.B(n_652),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_694),
.B(n_273),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_714),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_702),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_706),
.B(n_288),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_704),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_704),
.B(n_652),
.Y(n_919)
);

AOI22x1_ASAP7_75t_L g920 ( 
.A1(n_705),
.A2(n_660),
.B1(n_659),
.B2(n_267),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_705),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_707),
.B(n_652),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_773),
.B(n_290),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_802),
.A2(n_614),
.B1(n_660),
.B2(n_659),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_707),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_712),
.B(n_652),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_765),
.B(n_247),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_821),
.B(n_247),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_759),
.B(n_688),
.Y(n_929)
);

OR2x6_ASAP7_75t_L g930 ( 
.A(n_812),
.B(n_643),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_715),
.B(n_342),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_724),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_724),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_731),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_712),
.B(n_652),
.Y(n_935)
);

AOI221xp5_ASAP7_75t_L g936 ( 
.A1(n_782),
.A2(n_465),
.B1(n_457),
.B2(n_395),
.C(n_396),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_783),
.B(n_297),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_731),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_720),
.B(n_652),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_720),
.B(n_652),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_734),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_726),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_726),
.B(n_728),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_728),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_733),
.B(n_657),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_733),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_802),
.A2(n_614),
.B1(n_660),
.B2(n_645),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_744),
.B(n_662),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_734),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_744),
.B(n_662),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_749),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_749),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_736),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_715),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_742),
.B(n_342),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_736),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_796),
.B(n_305),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_757),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_757),
.B(n_662),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_767),
.B(n_688),
.Y(n_960)
);

AND2x2_ASAP7_75t_SL g961 ( 
.A(n_708),
.B(n_254),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_766),
.Y(n_962)
);

OAI22xp33_ASAP7_75t_L g963 ( 
.A1(n_812),
.A2(n_276),
.B1(n_277),
.B2(n_272),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_770),
.B(n_342),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_802),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_774),
.B(n_308),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_812),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_766),
.B(n_778),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_778),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_740),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_781),
.B(n_662),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_740),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_781),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_795),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_818),
.A2(n_643),
.B1(n_614),
.B2(n_276),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_812),
.B(n_645),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_829),
.A2(n_663),
.B(n_608),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_795),
.B(n_663),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_805),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_770),
.B(n_342),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_805),
.B(n_663),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_751),
.Y(n_982)
);

AND2x2_ASAP7_75t_SL g983 ( 
.A(n_747),
.B(n_380),
.Y(n_983)
);

NAND2x1_ASAP7_75t_L g984 ( 
.A(n_699),
.B(n_614),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_806),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_716),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_721),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_713),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_817),
.B(n_643),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_806),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_816),
.B(n_663),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_729),
.B(n_250),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_816),
.B(n_645),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_709),
.B(n_645),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_839),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_729),
.B(n_271),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_709),
.B(n_604),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_741),
.Y(n_998)
);

NOR3xp33_ASAP7_75t_L g999 ( 
.A(n_838),
.B(n_320),
.C(n_318),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_839),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_729),
.B(n_271),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_817),
.B(n_691),
.Y(n_1002)
);

NAND2x1_ASAP7_75t_L g1003 ( 
.A(n_699),
.B(n_607),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_723),
.B(n_271),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_840),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_741),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_761),
.B(n_271),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_739),
.B(n_271),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_709),
.A2(n_421),
.B1(n_380),
.B2(n_272),
.Y(n_1009)
);

OAI22x1_ASAP7_75t_SL g1010 ( 
.A1(n_717),
.A2(n_328),
.B1(n_337),
.B2(n_327),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_752),
.B(n_604),
.Y(n_1011)
);

BUFx8_ASAP7_75t_L g1012 ( 
.A(n_760),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_750),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_772),
.B(n_604),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_725),
.B(n_341),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_840),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_727),
.B(n_343),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_817),
.A2(n_421),
.B1(n_277),
.B2(n_284),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_785),
.B(n_604),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_847),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_822),
.B(n_604),
.Y(n_1021)
);

NOR2xp67_ASAP7_75t_SL g1022 ( 
.A(n_713),
.B(n_271),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_817),
.B(n_681),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_830),
.B(n_607),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_847),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_849),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_833),
.B(n_607),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_909),
.B(n_748),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_874),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_907),
.A2(n_809),
.B(n_769),
.Y(n_1030)
);

AOI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_854),
.A2(n_746),
.B(n_820),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_869),
.B(n_748),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_870),
.A2(n_809),
.B(n_769),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_876),
.B(n_721),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_910),
.Y(n_1035)
);

INVx3_ASAP7_75t_SL g1036 ( 
.A(n_987),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_863),
.A2(n_819),
.B(n_747),
.Y(n_1037)
);

OAI21xp33_ASAP7_75t_L g1038 ( 
.A1(n_857),
.A2(n_754),
.B(n_841),
.Y(n_1038)
);

OAI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_936),
.A2(n_754),
.B(n_823),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_954),
.A2(n_851),
.B1(n_825),
.B2(n_834),
.Y(n_1040)
);

AO21x1_ASAP7_75t_L g1041 ( 
.A1(n_1008),
.A2(n_284),
.B(n_279),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_913),
.A2(n_819),
.B(n_768),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_864),
.A2(n_849),
.B(n_753),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_954),
.A2(n_751),
.B1(n_790),
.B2(n_760),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_895),
.B(n_791),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_880),
.A2(n_853),
.B(n_753),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_884),
.B(n_794),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_911),
.B(n_713),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_994),
.A2(n_756),
.B(n_750),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_885),
.A2(n_853),
.B(n_776),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_868),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_997),
.A2(n_905),
.B(n_899),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1021),
.A2(n_768),
.B(n_700),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_989),
.Y(n_1054)
);

INVx11_ASAP7_75t_L g1055 ( 
.A(n_1012),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_871),
.B(n_738),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1011),
.A2(n_700),
.B(n_699),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_871),
.B(n_738),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1014),
.A2(n_764),
.B(n_700),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_889),
.B(n_730),
.Y(n_1060)
);

BUFx4f_ASAP7_75t_L g1061 ( 
.A(n_961),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_873),
.B(n_738),
.Y(n_1062)
);

OA22x2_ASAP7_75t_L g1063 ( 
.A1(n_910),
.A2(n_730),
.B1(n_711),
.B2(n_386),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_1003),
.A2(n_891),
.B(n_886),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_L g1065 ( 
.A(n_986),
.B(n_563),
.Y(n_1065)
);

AO22x1_ASAP7_75t_L g1066 ( 
.A1(n_999),
.A2(n_1017),
.B1(n_1015),
.B2(n_937),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_885),
.A2(n_776),
.B(n_756),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1019),
.A2(n_792),
.B(n_764),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_873),
.B(n_745),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1023),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_911),
.B(n_722),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_911),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_911),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_892),
.A2(n_792),
.B(n_764),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_877),
.B(n_745),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_882),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_881),
.B(n_745),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_887),
.B(n_842),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_887),
.B(n_872),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_872),
.B(n_842),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1023),
.A2(n_790),
.B1(n_760),
.B2(n_832),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_989),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_893),
.A2(n_837),
.B(n_792),
.Y(n_1083)
);

O2A1O1Ixp5_ASAP7_75t_L g1084 ( 
.A1(n_1007),
.A2(n_842),
.B(n_788),
.C(n_798),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_882),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_888),
.A2(n_850),
.B(n_837),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_931),
.B(n_837),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_947),
.A2(n_965),
.B1(n_911),
.B2(n_976),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_965),
.A2(n_836),
.B1(n_827),
.B2(n_286),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_888),
.A2(n_850),
.B(n_758),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_894),
.A2(n_850),
.B(n_758),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_898),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_914),
.A2(n_286),
.B(n_304),
.C(n_279),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_856),
.B(n_780),
.Y(n_1094)
);

NAND2x1_ASAP7_75t_L g1095 ( 
.A(n_898),
.B(n_722),
.Y(n_1095)
);

NOR2x1p5_ASAP7_75t_SL g1096 ( 
.A(n_976),
.B(n_780),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_916),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_993),
.A2(n_852),
.B(n_798),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_894),
.A2(n_758),
.B(n_722),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_856),
.B(n_788),
.Y(n_1100)
);

AND2x2_ASAP7_75t_SL g1101 ( 
.A(n_961),
.B(n_304),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_916),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_861),
.B(n_918),
.Y(n_1103)
);

AO21x1_ASAP7_75t_L g1104 ( 
.A1(n_955),
.A2(n_316),
.B(n_313),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1024),
.A2(n_758),
.B(n_722),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_861),
.B(n_918),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_859),
.B(n_800),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_SL g1108 ( 
.A(n_967),
.B(n_313),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_921),
.B(n_852),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1027),
.A2(n_758),
.B(n_722),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_966),
.B(n_719),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_855),
.A2(n_810),
.B(n_775),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_921),
.B(n_800),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_879),
.B(n_563),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_943),
.A2(n_811),
.B(n_803),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_925),
.B(n_803),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_860),
.B(n_811),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_883),
.A2(n_810),
.B(n_775),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_988),
.A2(n_810),
.B(n_775),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_984),
.A2(n_810),
.B(n_775),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_984),
.A2(n_810),
.B(n_775),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1003),
.A2(n_996),
.B(n_992),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_1002),
.Y(n_1123)
);

AOI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_917),
.A2(n_711),
.B(n_317),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_982),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_924),
.A2(n_317),
.B1(n_322),
.B2(n_316),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_925),
.B(n_813),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_942),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_L g1129 ( 
.A(n_858),
.B(n_980),
.C(n_964),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1002),
.B(n_824),
.Y(n_1130)
);

NOR2xp67_ASAP7_75t_L g1131 ( 
.A(n_879),
.B(n_923),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_977),
.A2(n_814),
.B(n_813),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_942),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_944),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_944),
.B(n_814),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_946),
.B(n_815),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1001),
.A2(n_845),
.B(n_824),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_968),
.A2(n_845),
.B(n_824),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_957),
.B(n_815),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_878),
.B(n_681),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_919),
.A2(n_845),
.B(n_824),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1004),
.A2(n_831),
.B(n_828),
.C(n_323),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_987),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_929),
.A2(n_323),
.B(n_325),
.C(n_322),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_922),
.A2(n_845),
.B(n_824),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_926),
.A2(n_845),
.B(n_608),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_946),
.B(n_828),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_935),
.A2(n_608),
.B(n_600),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_951),
.B(n_831),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_951),
.B(n_832),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_890),
.A2(n_350),
.B(n_348),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_952),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_952),
.B(n_832),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_960),
.B(n_896),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_928),
.B(n_351),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_989),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1002),
.B(n_375),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_945),
.A2(n_950),
.B(n_948),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_958),
.B(n_832),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_958),
.B(n_832),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_939),
.A2(n_608),
.B(n_600),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_959),
.A2(n_790),
.B(n_760),
.Y(n_1162)
);

NAND2x2_ASAP7_75t_L g1163 ( 
.A(n_967),
.B(n_691),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_962),
.B(n_832),
.Y(n_1164)
);

BUFx4f_ASAP7_75t_L g1165 ( 
.A(n_930),
.Y(n_1165)
);

AO21x1_ASAP7_75t_L g1166 ( 
.A1(n_963),
.A2(n_345),
.B(n_325),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_865),
.B(n_355),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_930),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_940),
.A2(n_608),
.B(n_600),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_971),
.A2(n_668),
.B(n_683),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_904),
.B(n_345),
.Y(n_1171)
);

O2A1O1Ixp5_ASAP7_75t_L g1172 ( 
.A1(n_902),
.A2(n_347),
.B(n_398),
.C(n_346),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1018),
.A2(n_347),
.B1(n_398),
.B2(n_346),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_962),
.B(n_969),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_912),
.B(n_375),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_975),
.B(n_375),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_969),
.B(n_760),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_973),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_900),
.B(n_357),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_978),
.A2(n_608),
.B(n_600),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_981),
.A2(n_608),
.B(n_600),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_973),
.B(n_375),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_927),
.A2(n_455),
.B(n_410),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_991),
.A2(n_608),
.B(n_600),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1012),
.B(n_299),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_901),
.B(n_903),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_974),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_974),
.B(n_760),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_983),
.B(n_1012),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1010),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_979),
.A2(n_455),
.B(n_410),
.C(n_603),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_979),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_985),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_930),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_930),
.A2(n_608),
.B(n_600),
.Y(n_1195)
);

NOR2x1_ASAP7_75t_R g1196 ( 
.A(n_1010),
.B(n_360),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_985),
.A2(n_600),
.B(n_607),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_990),
.A2(n_600),
.B(n_607),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_990),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1009),
.B(n_790),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_995),
.B(n_362),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_983),
.B(n_375),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_983),
.B(n_299),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_995),
.A2(n_1005),
.B1(n_1016),
.B2(n_1000),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1026),
.A2(n_668),
.B1(n_683),
.B2(n_686),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1026),
.B(n_790),
.Y(n_1206)
);

AND2x2_ASAP7_75t_SL g1207 ( 
.A(n_1000),
.B(n_378),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1005),
.A2(n_610),
.B(n_668),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1016),
.B(n_363),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1025),
.B(n_790),
.Y(n_1210)
);

AND2x2_ASAP7_75t_SL g1211 ( 
.A(n_1020),
.B(n_395),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1025),
.B(n_683),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_920),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1020),
.A2(n_610),
.B(n_668),
.Y(n_1214)
);

INVx6_ASAP7_75t_L g1215 ( 
.A(n_920),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_862),
.A2(n_610),
.B(n_596),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_862),
.B(n_683),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_866),
.A2(n_610),
.B(n_596),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_866),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_867),
.Y(n_1220)
);

INVx11_ASAP7_75t_L g1221 ( 
.A(n_1022),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1124),
.A2(n_404),
.B(n_430),
.C(n_396),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1219),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1028),
.B(n_1032),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1088),
.B(n_867),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1192),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1072),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1034),
.B(n_875),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1207),
.B(n_875),
.Y(n_1229)
);

O2A1O1Ixp5_ASAP7_75t_L g1230 ( 
.A1(n_1066),
.A2(n_1022),
.B(n_906),
.C(n_908),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1029),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1170),
.A2(n_906),
.B(n_897),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1038),
.A2(n_1013),
.B1(n_1006),
.B2(n_998),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1029),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1052),
.A2(n_908),
.B(n_897),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1129),
.A2(n_1013),
.B1(n_1006),
.B2(n_998),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1039),
.B(n_915),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1086),
.A2(n_932),
.B(n_915),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1064),
.A2(n_933),
.B(n_932),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1090),
.A2(n_934),
.B(n_933),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1091),
.A2(n_938),
.B(n_934),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1192),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1076),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1219),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1074),
.A2(n_941),
.B(n_938),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1125),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1051),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1092),
.Y(n_1248)
);

AOI221x1_ASAP7_75t_L g1249 ( 
.A1(n_1031),
.A2(n_972),
.B1(n_970),
.B2(n_956),
.C(n_953),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1036),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1060),
.B(n_941),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1083),
.A2(n_1059),
.B(n_1057),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1097),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1129),
.A2(n_1186),
.B1(n_1047),
.B2(n_1060),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1123),
.B(n_949),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1111),
.B(n_299),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1207),
.B(n_949),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1070),
.B(n_953),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1123),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1035),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1068),
.A2(n_970),
.B(n_956),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1035),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1036),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_R g1264 ( 
.A(n_1185),
.B(n_117),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1070),
.B(n_972),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1078),
.A2(n_610),
.B(n_605),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1093),
.A2(n_458),
.B(n_462),
.C(n_464),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1046),
.A2(n_626),
.B(n_605),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1099),
.A2(n_626),
.B(n_605),
.Y(n_1269)
);

OAI22x1_ASAP7_75t_L g1270 ( 
.A1(n_1190),
.A2(n_368),
.B1(n_370),
.B2(n_373),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1211),
.B(n_683),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_SL g1272 ( 
.A1(n_1202),
.A2(n_1144),
.B(n_1175),
.C(n_1182),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1211),
.B(n_686),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1183),
.A2(n_404),
.B(n_430),
.C(n_445),
.Y(n_1274)
);

NOR3xp33_ASAP7_75t_SL g1275 ( 
.A(n_1151),
.B(n_382),
.C(n_379),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1045),
.B(n_573),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1186),
.A2(n_464),
.B(n_445),
.C(n_447),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1079),
.A2(n_1202),
.B(n_1175),
.Y(n_1278)
);

CKINVDCx16_ASAP7_75t_R g1279 ( 
.A(n_1143),
.Y(n_1279)
);

NOR3xp33_ASAP7_75t_L g1280 ( 
.A(n_1179),
.B(n_388),
.C(n_387),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1201),
.B(n_686),
.Y(n_1281)
);

BUFx12f_ASAP7_75t_L g1282 ( 
.A(n_1123),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1101),
.B(n_389),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1173),
.A2(n_462),
.B(n_458),
.C(n_447),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1123),
.B(n_375),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1072),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1163),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1061),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1101),
.A2(n_448),
.B(n_585),
.C(n_581),
.Y(n_1289)
);

AO22x1_ASAP7_75t_L g1290 ( 
.A1(n_1179),
.A2(n_406),
.B1(n_390),
.B2(n_391),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1201),
.B(n_686),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1171),
.A2(n_448),
.B(n_573),
.C(n_575),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1065),
.B(n_315),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1134),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1209),
.B(n_686),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1072),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1072),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1220),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1209),
.B(n_595),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1085),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1102),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1155),
.A2(n_579),
.B(n_575),
.C(n_580),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1139),
.B(n_595),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1139),
.B(n_1140),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1155),
.B(n_315),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1073),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1204),
.A2(n_392),
.B1(n_399),
.B2(n_400),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_SL g1308 ( 
.A1(n_1182),
.A2(n_591),
.B(n_578),
.C(n_579),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1128),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1133),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1152),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1178),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1050),
.A2(n_630),
.B(n_626),
.Y(n_1313)
);

INVxp67_ASAP7_75t_SL g1314 ( 
.A(n_1073),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1187),
.B(n_597),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1193),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1199),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1040),
.B(n_597),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1103),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1194),
.B(n_578),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1063),
.B(n_1167),
.Y(n_1321)
);

NOR2xp67_ASAP7_75t_L g1322 ( 
.A(n_1131),
.B(n_118),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1055),
.Y(n_1323)
);

NOR3xp33_ASAP7_75t_SL g1324 ( 
.A(n_1167),
.B(n_403),
.C(n_401),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1106),
.Y(n_1325)
);

AND2x6_ASAP7_75t_L g1326 ( 
.A(n_1073),
.B(n_1168),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1094),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1154),
.A2(n_619),
.B1(n_601),
.B2(n_603),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_SL g1329 ( 
.A1(n_1157),
.A2(n_580),
.B(n_581),
.C(n_585),
.Y(n_1329)
);

NAND2x1p5_ASAP7_75t_L g1330 ( 
.A(n_1073),
.B(n_601),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1126),
.A2(n_315),
.B1(n_344),
.B2(n_349),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1054),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1203),
.B(n_315),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1174),
.A2(n_405),
.B1(n_415),
.B2(n_422),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1061),
.A2(n_592),
.B(n_591),
.C(n_432),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_R g1336 ( 
.A(n_1054),
.B(n_123),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1107),
.A2(n_592),
.B(n_423),
.C(n_434),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1067),
.A2(n_630),
.B(n_655),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1082),
.B(n_679),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1100),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1082),
.B(n_679),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1194),
.A2(n_438),
.B1(n_437),
.B2(n_436),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1053),
.A2(n_630),
.B(n_616),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1080),
.B(n_616),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1063),
.B(n_344),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1075),
.A2(n_649),
.B(n_619),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1107),
.A2(n_453),
.B(n_440),
.C(n_441),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1077),
.A2(n_649),
.B(n_624),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1165),
.A2(n_443),
.B1(n_444),
.B2(n_449),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1217),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1109),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1080),
.B(n_624),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1156),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1158),
.A2(n_653),
.B(n_632),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1056),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1168),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_SL g1357 ( 
.A1(n_1157),
.A2(n_653),
.B(n_625),
.C(n_628),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1156),
.B(n_1114),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1168),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1168),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1165),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1058),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1087),
.B(n_679),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1087),
.B(n_625),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1206),
.A2(n_642),
.B(n_628),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1166),
.A2(n_344),
.B1(n_349),
.B2(n_450),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1117),
.A2(n_459),
.B(n_460),
.C(n_549),
.Y(n_1367)
);

NOR2x1_ASAP7_75t_R g1368 ( 
.A(n_1189),
.B(n_541),
.Y(n_1368)
);

AOI22x1_ASAP7_75t_L g1369 ( 
.A1(n_1213),
.A2(n_655),
.B1(n_639),
.B2(n_632),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1113),
.Y(n_1370)
);

OR2x6_ASAP7_75t_L g1371 ( 
.A(n_1130),
.B(n_541),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1117),
.B(n_633),
.Y(n_1372)
);

NAND2xp33_ASAP7_75t_SL g1373 ( 
.A(n_1108),
.B(n_543),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1191),
.A2(n_656),
.B(n_642),
.C(n_639),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_SL g1375 ( 
.A1(n_1176),
.A2(n_666),
.B(n_633),
.C(n_656),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_L g1376 ( 
.A(n_1044),
.B(n_543),
.C(n_544),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1196),
.Y(n_1377)
);

OAI22x1_ASAP7_75t_L g1378 ( 
.A1(n_1048),
.A2(n_549),
.B1(n_544),
.B2(n_349),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1062),
.B(n_665),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1130),
.A2(n_665),
.B(n_666),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1116),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1037),
.A2(n_667),
.B(n_682),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1069),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1095),
.Y(n_1384)
);

AOI221xp5_ASAP7_75t_L g1385 ( 
.A1(n_1089),
.A2(n_667),
.B1(n_344),
.B2(n_349),
.C(n_678),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1172),
.A2(n_690),
.B(n_682),
.C(n_678),
.Y(n_1386)
);

NOR3xp33_ASAP7_75t_SL g1387 ( 
.A(n_1048),
.B(n_10),
.C(n_12),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1127),
.B(n_671),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1250),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1312),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1359),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_SL g1392 ( 
.A1(n_1337),
.A2(n_1071),
.B(n_1176),
.C(n_1150),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1231),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1249),
.A2(n_1104),
.A3(n_1041),
.B(n_1033),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1252),
.A2(n_1030),
.B(n_1042),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1278),
.A2(n_1043),
.B(n_1208),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1254),
.B(n_1081),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1246),
.B(n_1122),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1231),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1263),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1224),
.B(n_1135),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1225),
.A2(n_1110),
.B(n_1105),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1312),
.Y(n_1403)
);

AOI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1222),
.A2(n_1205),
.B1(n_1142),
.B2(n_1149),
.C(n_1147),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1247),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1225),
.A2(n_1138),
.B(n_1071),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1300),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1283),
.A2(n_1163),
.B1(n_1215),
.B2(n_1200),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1304),
.A2(n_1162),
.B(n_1049),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1333),
.B(n_671),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1316),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1223),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1319),
.B(n_1136),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1325),
.B(n_1212),
.Y(n_1414)
);

AOI221xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1277),
.A2(n_1214),
.B1(n_1098),
.B2(n_1115),
.C(n_1164),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1281),
.A2(n_1153),
.B(n_1159),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1291),
.A2(n_1112),
.B(n_1118),
.Y(n_1417)
);

NAND2x1p5_ASAP7_75t_L g1418 ( 
.A(n_1259),
.B(n_1137),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1359),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1295),
.A2(n_1119),
.B(n_1120),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1378),
.A2(n_1145),
.A3(n_1141),
.B(n_1160),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1359),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1301),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1234),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1351),
.B(n_1096),
.Y(n_1425)
);

AOI221x1_ASAP7_75t_L g1426 ( 
.A1(n_1335),
.A2(n_1218),
.B1(n_1216),
.B2(n_1188),
.C(n_1177),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1363),
.A2(n_1121),
.B(n_1210),
.Y(n_1427)
);

AO21x1_ASAP7_75t_L g1428 ( 
.A1(n_1318),
.A2(n_1198),
.B(n_1197),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1239),
.A2(n_1132),
.B(n_1084),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1309),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1230),
.A2(n_1146),
.B(n_1181),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1310),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1283),
.A2(n_1195),
.B(n_1184),
.C(n_1180),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1234),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1370),
.B(n_1215),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1363),
.A2(n_1148),
.B(n_1161),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1244),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1232),
.A2(n_1169),
.B(n_1215),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1311),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1317),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1364),
.A2(n_1221),
.B(n_690),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1280),
.A2(n_690),
.B1(n_682),
.B2(n_678),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1323),
.Y(n_1443)
);

BUFx10_ASAP7_75t_L g1444 ( 
.A(n_1321),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1381),
.B(n_671),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1279),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1321),
.A2(n_1305),
.B(n_1337),
.C(n_1237),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1324),
.B(n_690),
.C(n_682),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1367),
.A2(n_678),
.A3(n_674),
.B(n_671),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_SL g1450 ( 
.A1(n_1347),
.A2(n_674),
.B(n_235),
.C(n_234),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1235),
.A2(n_674),
.B(n_679),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1245),
.A2(n_674),
.B(n_171),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1260),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1298),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1260),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1251),
.B(n_679),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1238),
.A2(n_679),
.B(n_226),
.Y(n_1457)
);

AO21x1_ASAP7_75t_L g1458 ( 
.A1(n_1285),
.A2(n_1228),
.B(n_1372),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1251),
.B(n_679),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1243),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1261),
.A2(n_169),
.B(n_222),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1256),
.B(n_679),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1327),
.B(n_12),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1359),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_SL g1465 ( 
.A1(n_1347),
.A2(n_1367),
.B(n_1289),
.C(n_1335),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1360),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1293),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1237),
.A2(n_13),
.B(n_15),
.C(n_17),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1275),
.A2(n_17),
.B(n_18),
.C(n_24),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1272),
.A2(n_221),
.B(n_208),
.Y(n_1470)
);

AO32x2_ASAP7_75t_L g1471 ( 
.A1(n_1334),
.A2(n_30),
.A3(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_1471)
);

A2O1A1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1275),
.A2(n_33),
.B(n_38),
.C(n_39),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1331),
.A2(n_39),
.B(n_40),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1248),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1253),
.Y(n_1475)
);

BUFx2_ASAP7_75t_R g1476 ( 
.A(n_1361),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1356),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1262),
.B(n_40),
.Y(n_1478)
);

NOR4xp25_ASAP7_75t_L g1479 ( 
.A(n_1277),
.B(n_45),
.C(n_47),
.D(n_49),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1358),
.B(n_49),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1282),
.B(n_202),
.Y(n_1481)
);

O2A1O1Ixp5_ASAP7_75t_SL g1482 ( 
.A1(n_1285),
.A2(n_50),
.B(n_53),
.C(n_55),
.Y(n_1482)
);

AO32x2_ASAP7_75t_L g1483 ( 
.A1(n_1307),
.A2(n_53),
.A3(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_1483)
);

O2A1O1Ixp33_ASAP7_75t_L g1484 ( 
.A1(n_1289),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1340),
.B(n_65),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1382),
.A2(n_201),
.B(n_199),
.Y(n_1486)
);

AOI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1354),
.A2(n_198),
.B(n_196),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1355),
.B(n_69),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1240),
.A2(n_194),
.B(n_186),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1241),
.A2(n_177),
.B(n_176),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1302),
.A2(n_70),
.B(n_72),
.C(n_73),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1362),
.B(n_1383),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1294),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1233),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1276),
.B(n_72),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1343),
.A2(n_1269),
.B(n_1266),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1258),
.B(n_73),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1313),
.A2(n_167),
.B(n_161),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1288),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1338),
.A2(n_1365),
.B(n_1271),
.Y(n_1500)
);

AO31x2_ASAP7_75t_L g1501 ( 
.A1(n_1346),
.A2(n_75),
.A3(n_76),
.B(n_77),
.Y(n_1501)
);

AO31x2_ASAP7_75t_L g1502 ( 
.A1(n_1348),
.A2(n_80),
.A3(n_81),
.B(n_82),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1272),
.A2(n_160),
.B(n_158),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1303),
.A2(n_1299),
.B(n_1388),
.Y(n_1504)
);

NAND2x1_ASAP7_75t_L g1505 ( 
.A(n_1326),
.B(n_157),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1344),
.A2(n_155),
.B(n_143),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1255),
.A2(n_142),
.B(n_134),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1345),
.B(n_80),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1258),
.Y(n_1509)
);

AO32x2_ASAP7_75t_L g1510 ( 
.A1(n_1287),
.A2(n_81),
.A3(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1255),
.A2(n_133),
.B(n_129),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_SL g1512 ( 
.A(n_1368),
.B(n_86),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1352),
.A2(n_128),
.B(n_124),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1349),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1226),
.Y(n_1515)
);

AOI221x1_ASAP7_75t_L g1516 ( 
.A1(n_1270),
.A2(n_89),
.B1(n_91),
.B2(n_94),
.C(n_95),
.Y(n_1516)
);

INVx4_ASAP7_75t_SL g1517 ( 
.A(n_1326),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1265),
.B(n_94),
.Y(n_1518)
);

NAND2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1259),
.B(n_96),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1320),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1324),
.A2(n_1328),
.B(n_1273),
.C(n_1229),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1265),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1339),
.A2(n_98),
.B(n_1341),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1376),
.A2(n_1236),
.B(n_1257),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1290),
.B(n_1320),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1330),
.A2(n_1380),
.B(n_1369),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1360),
.Y(n_1527)
);

NOR2x1_ASAP7_75t_SL g1528 ( 
.A(n_1227),
.B(n_1306),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1350),
.B(n_1242),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1264),
.B(n_1342),
.Y(n_1530)
);

INVx2_ASAP7_75t_SL g1531 ( 
.A(n_1360),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1339),
.A2(n_1341),
.B(n_1379),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1332),
.B(n_1353),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1331),
.B(n_1366),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1332),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1386),
.A2(n_1268),
.B(n_1375),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1314),
.A2(n_1268),
.B(n_1315),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1284),
.A2(n_1322),
.B(n_1267),
.C(n_1366),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1353),
.B(n_1286),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1371),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1286),
.B(n_1296),
.Y(n_1541)
);

BUFx2_ASAP7_75t_R g1542 ( 
.A(n_1296),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1326),
.B(n_1371),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1377),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1264),
.B(n_1227),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1371),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1384),
.A2(n_1268),
.B(n_1227),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1330),
.Y(n_1548)
);

AOI221x1_ASAP7_75t_L g1549 ( 
.A1(n_1373),
.A2(n_1387),
.B1(n_1384),
.B2(n_1227),
.C(n_1297),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1308),
.Y(n_1550)
);

AO31x2_ASAP7_75t_L g1551 ( 
.A1(n_1375),
.A2(n_1357),
.A3(n_1329),
.B(n_1387),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1308),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1297),
.B(n_1306),
.Y(n_1553)
);

BUFx4_ASAP7_75t_SL g1554 ( 
.A(n_1336),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1297),
.A2(n_1306),
.B(n_1357),
.Y(n_1555)
);

AO31x2_ASAP7_75t_L g1556 ( 
.A1(n_1329),
.A2(n_1374),
.A3(n_1326),
.B(n_1385),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1326),
.A2(n_1297),
.B1(n_1306),
.B2(n_1336),
.Y(n_1557)
);

AO31x2_ASAP7_75t_L g1558 ( 
.A1(n_1274),
.A2(n_1249),
.A3(n_1252),
.B(n_1378),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1292),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1239),
.A2(n_1232),
.B(n_1170),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1252),
.A2(n_863),
.B(n_870),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1312),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1333),
.B(n_1251),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1312),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1252),
.A2(n_863),
.B(n_870),
.Y(n_1565)
);

OAI22x1_ASAP7_75t_L g1566 ( 
.A1(n_1254),
.A2(n_1321),
.B1(n_1283),
.B2(n_730),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1246),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1252),
.A2(n_863),
.B(n_870),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1224),
.B(n_1319),
.Y(n_1569)
);

AO31x2_ASAP7_75t_L g1570 ( 
.A1(n_1249),
.A2(n_1252),
.A3(n_1378),
.B(n_880),
.Y(n_1570)
);

AO31x2_ASAP7_75t_L g1571 ( 
.A1(n_1249),
.A2(n_1252),
.A3(n_1378),
.B(n_880),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1249),
.A2(n_1230),
.B(n_1232),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1400),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1391),
.Y(n_1574)
);

INVx6_ASAP7_75t_L g1575 ( 
.A(n_1517),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_1514),
.B2(n_1563),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1397),
.A2(n_1530),
.B1(n_1467),
.B2(n_1512),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1544),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1391),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1405),
.Y(n_1580)
);

BUFx4f_ASAP7_75t_SL g1581 ( 
.A(n_1443),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1473),
.A2(n_1516),
.B(n_1520),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1411),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1512),
.A2(n_1525),
.B1(n_1508),
.B2(n_1495),
.Y(n_1584)
);

INVx4_ASAP7_75t_L g1585 ( 
.A(n_1517),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1495),
.A2(n_1518),
.B1(n_1497),
.B2(n_1480),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1533),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1439),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1407),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1519),
.A2(n_1444),
.B1(n_1497),
.B2(n_1518),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1403),
.Y(n_1591)
);

BUFx10_ASAP7_75t_L g1592 ( 
.A(n_1389),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1499),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1519),
.A2(n_1444),
.B1(n_1477),
.B2(n_1569),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1569),
.A2(n_1473),
.B1(n_1481),
.B2(n_1509),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1446),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1447),
.A2(n_1522),
.B1(n_1492),
.B2(n_1413),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1533),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1564),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1488),
.A2(n_1485),
.B1(n_1463),
.B2(n_1494),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1423),
.Y(n_1601)
);

NAND2x1p5_ASAP7_75t_L g1602 ( 
.A(n_1455),
.B(n_1393),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1488),
.A2(n_1485),
.B1(n_1463),
.B2(n_1500),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1424),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1492),
.A2(n_1413),
.B1(n_1408),
.B2(n_1521),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1562),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1430),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1454),
.Y(n_1608)
);

INVx6_ASAP7_75t_L g1609 ( 
.A(n_1517),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1479),
.A2(n_1481),
.B1(n_1478),
.B2(n_1393),
.Y(n_1610)
);

INVx3_ASAP7_75t_SL g1611 ( 
.A(n_1567),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1434),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1500),
.A2(n_1401),
.B1(n_1481),
.B2(n_1410),
.Y(n_1613)
);

INVx6_ASAP7_75t_L g1614 ( 
.A(n_1391),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1401),
.A2(n_1524),
.B1(n_1559),
.B2(n_1432),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_SL g1616 ( 
.A1(n_1540),
.A2(n_1503),
.B1(n_1470),
.B2(n_1399),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1412),
.B(n_1437),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1474),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1476),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1479),
.A2(n_1453),
.B1(n_1546),
.B2(n_1543),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1440),
.Y(n_1621)
);

INVx6_ASAP7_75t_L g1622 ( 
.A(n_1422),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1475),
.Y(n_1623)
);

NAND2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1545),
.B(n_1557),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1493),
.Y(n_1625)
);

BUFx12f_ASAP7_75t_L g1626 ( 
.A(n_1422),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1553),
.Y(n_1627)
);

BUFx8_ASAP7_75t_SL g1628 ( 
.A(n_1422),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1529),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1529),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1561),
.A2(n_1568),
.B(n_1565),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1535),
.B(n_1460),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1515),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1476),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1539),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1524),
.A2(n_1414),
.B1(n_1458),
.B2(n_1503),
.Y(n_1636)
);

INVx6_ASAP7_75t_L g1637 ( 
.A(n_1464),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1462),
.A2(n_1538),
.B1(n_1465),
.B2(n_1472),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1539),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1414),
.A2(n_1435),
.B1(n_1543),
.B2(n_1542),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1445),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1435),
.B(n_1541),
.Y(n_1642)
);

CKINVDCx6p67_ASAP7_75t_R g1643 ( 
.A(n_1464),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1542),
.A2(n_1425),
.B1(n_1548),
.B2(n_1469),
.Y(n_1644)
);

INVx8_ASAP7_75t_L g1645 ( 
.A(n_1464),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1425),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1504),
.A2(n_1523),
.B1(n_1456),
.B2(n_1459),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1398),
.A2(n_1468),
.B1(n_1505),
.B2(n_1448),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1466),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_1466),
.Y(n_1650)
);

OAI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1549),
.A2(n_1445),
.B1(n_1510),
.B2(n_1483),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1506),
.A2(n_1513),
.B1(n_1396),
.B2(n_1404),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1466),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1532),
.A2(n_1409),
.B1(n_1404),
.B2(n_1541),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1429),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1554),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1419),
.Y(n_1657)
);

CKINVDCx11_ASAP7_75t_R g1658 ( 
.A(n_1550),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1419),
.Y(n_1659)
);

INVx6_ASAP7_75t_L g1660 ( 
.A(n_1528),
.Y(n_1660)
);

INVx6_ASAP7_75t_L g1661 ( 
.A(n_1531),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1396),
.A2(n_1552),
.B1(n_1428),
.B2(n_1483),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1433),
.A2(n_1441),
.B1(n_1537),
.B2(n_1547),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1527),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1560),
.Y(n_1665)
);

CKINVDCx16_ASAP7_75t_R g1666 ( 
.A(n_1442),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1484),
.B(n_1491),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1483),
.A2(n_1537),
.B1(n_1471),
.B2(n_1406),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1449),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1498),
.A2(n_1486),
.B1(n_1461),
.B2(n_1490),
.Y(n_1670)
);

BUFx8_ASAP7_75t_L g1671 ( 
.A(n_1510),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1501),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1555),
.Y(n_1673)
);

CKINVDCx14_ASAP7_75t_R g1674 ( 
.A(n_1471),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1501),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1431),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1501),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1502),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1510),
.A2(n_1471),
.B1(n_1426),
.B2(n_1536),
.Y(n_1679)
);

BUFx10_ASAP7_75t_L g1680 ( 
.A(n_1482),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1457),
.A2(n_1536),
.B1(n_1402),
.B2(n_1427),
.Y(n_1681)
);

OAI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1418),
.A2(n_1487),
.B1(n_1431),
.B2(n_1420),
.Y(n_1682)
);

INVxp33_ASAP7_75t_SL g1683 ( 
.A(n_1507),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1502),
.Y(n_1684)
);

BUFx12f_ASAP7_75t_L g1685 ( 
.A(n_1418),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1489),
.A2(n_1572),
.B1(n_1511),
.B2(n_1526),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1570),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1572),
.A2(n_1496),
.B1(n_1417),
.B2(n_1452),
.Y(n_1688)
);

CKINVDCx6p67_ASAP7_75t_R g1689 ( 
.A(n_1450),
.Y(n_1689)
);

CKINVDCx6p67_ASAP7_75t_R g1690 ( 
.A(n_1392),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1449),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1570),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1449),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1421),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1395),
.A2(n_1556),
.B1(n_1438),
.B2(n_1551),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1558),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1451),
.A2(n_1415),
.B1(n_1556),
.B2(n_1558),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1421),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_SL g1699 ( 
.A1(n_1556),
.A2(n_1551),
.B1(n_1416),
.B2(n_1558),
.Y(n_1699)
);

OAI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1436),
.A2(n_1415),
.B1(n_1551),
.B2(n_1570),
.Y(n_1700)
);

OAI21xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1571),
.A2(n_1421),
.B(n_1394),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1571),
.A2(n_1534),
.B1(n_1566),
.B2(n_854),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1571),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1394),
.Y(n_1704)
);

INVx4_ASAP7_75t_L g1705 ( 
.A(n_1394),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_854),
.B2(n_1038),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1424),
.Y(n_1707)
);

INVx6_ASAP7_75t_L g1708 ( 
.A(n_1517),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1390),
.Y(n_1709)
);

OAI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1512),
.A2(n_1473),
.B1(n_1467),
.B2(n_1254),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1534),
.A2(n_1283),
.B1(n_854),
.B2(n_1305),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1405),
.Y(n_1712)
);

BUFx3_ASAP7_75t_L g1713 ( 
.A(n_1477),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_SL g1714 ( 
.A1(n_1534),
.A2(n_1283),
.B1(n_854),
.B2(n_1305),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1405),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1407),
.Y(n_1716)
);

OAI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1512),
.A2(n_1473),
.B1(n_1467),
.B2(n_1254),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1405),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1400),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_854),
.B2(n_1038),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_854),
.B2(n_1038),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1405),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1443),
.Y(n_1723)
);

OAI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1512),
.A2(n_1473),
.B1(n_1467),
.B2(n_1254),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1405),
.Y(n_1725)
);

BUFx4_ASAP7_75t_SL g1726 ( 
.A(n_1544),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1407),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1424),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_854),
.B2(n_1038),
.Y(n_1729)
);

INVx6_ASAP7_75t_L g1730 ( 
.A(n_1517),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1424),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_854),
.B2(n_1038),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_854),
.B2(n_1038),
.Y(n_1733)
);

INVx6_ASAP7_75t_L g1734 ( 
.A(n_1517),
.Y(n_1734)
);

NAND2x1p5_ASAP7_75t_L g1735 ( 
.A(n_1455),
.B(n_1393),
.Y(n_1735)
);

CKINVDCx11_ASAP7_75t_R g1736 ( 
.A(n_1400),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1499),
.Y(n_1737)
);

BUFx12f_ASAP7_75t_L g1738 ( 
.A(n_1400),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1477),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1390),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1400),
.Y(n_1741)
);

INVx8_ASAP7_75t_L g1742 ( 
.A(n_1391),
.Y(n_1742)
);

BUFx12f_ASAP7_75t_L g1743 ( 
.A(n_1400),
.Y(n_1743)
);

BUFx8_ASAP7_75t_SL g1744 ( 
.A(n_1544),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1534),
.A2(n_1283),
.B1(n_854),
.B2(n_1305),
.Y(n_1745)
);

INVx8_ASAP7_75t_L g1746 ( 
.A(n_1391),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1499),
.Y(n_1747)
);

INVx8_ASAP7_75t_L g1748 ( 
.A(n_1391),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1405),
.Y(n_1749)
);

BUFx12f_ASAP7_75t_L g1750 ( 
.A(n_1400),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1443),
.Y(n_1751)
);

OAI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1447),
.A2(n_854),
.B(n_1038),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1499),
.Y(n_1753)
);

CKINVDCx11_ASAP7_75t_R g1754 ( 
.A(n_1400),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_854),
.B2(n_1038),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1477),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_SL g1757 ( 
.A1(n_1534),
.A2(n_1283),
.B1(n_854),
.B2(n_1305),
.Y(n_1757)
);

CKINVDCx20_ASAP7_75t_R g1758 ( 
.A(n_1400),
.Y(n_1758)
);

CKINVDCx11_ASAP7_75t_R g1759 ( 
.A(n_1400),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_SL g1760 ( 
.A1(n_1534),
.A2(n_1283),
.B1(n_854),
.B2(n_1305),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1424),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_SL g1762 ( 
.A1(n_1534),
.A2(n_1283),
.B1(n_854),
.B2(n_1305),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1477),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1534),
.A2(n_1566),
.B1(n_854),
.B2(n_1038),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1424),
.Y(n_1765)
);

CKINVDCx11_ASAP7_75t_R g1766 ( 
.A(n_1400),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1391),
.Y(n_1767)
);

BUFx2_ASAP7_75t_SL g1768 ( 
.A(n_1443),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1569),
.A2(n_854),
.B1(n_889),
.B2(n_1038),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1393),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1534),
.A2(n_1283),
.B1(n_854),
.B2(n_1305),
.Y(n_1771)
);

BUFx10_ASAP7_75t_L g1772 ( 
.A(n_1389),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1405),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1672),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1675),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1593),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1677),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1678),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1684),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1655),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1770),
.Y(n_1781)
);

BUFx2_ASAP7_75t_L g1782 ( 
.A(n_1587),
.Y(n_1782)
);

AND2x2_ASAP7_75t_SL g1783 ( 
.A(n_1668),
.B(n_1671),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1674),
.B(n_1646),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1655),
.Y(n_1785)
);

AO31x2_ASAP7_75t_L g1786 ( 
.A1(n_1663),
.A2(n_1691),
.A3(n_1693),
.B(n_1705),
.Y(n_1786)
);

AO21x2_ASAP7_75t_L g1787 ( 
.A1(n_1682),
.A2(n_1631),
.B(n_1700),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1685),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1704),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1703),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1669),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1669),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1598),
.Y(n_1793)
);

AOI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1654),
.A2(n_1667),
.B(n_1696),
.Y(n_1794)
);

OAI21x1_ASAP7_75t_L g1795 ( 
.A1(n_1688),
.A2(n_1686),
.B(n_1681),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1710),
.A2(n_1717),
.B1(n_1724),
.B2(n_1752),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1591),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1668),
.A2(n_1701),
.B(n_1662),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1710),
.A2(n_1717),
.B1(n_1724),
.B2(n_1711),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1585),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1687),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1599),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1585),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1737),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1714),
.A2(n_1757),
.B(n_1745),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1688),
.A2(n_1686),
.B(n_1681),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1707),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1692),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1696),
.Y(n_1809)
);

OAI21x1_ASAP7_75t_L g1810 ( 
.A1(n_1665),
.A2(n_1697),
.B(n_1694),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1698),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1705),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1575),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1690),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1674),
.B(n_1702),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1604),
.B(n_1612),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1580),
.Y(n_1817)
);

OR2x6_ASAP7_75t_L g1818 ( 
.A(n_1624),
.B(n_1610),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1583),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1712),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1728),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1715),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1676),
.Y(n_1823)
);

OAI21x1_ASAP7_75t_L g1824 ( 
.A1(n_1697),
.A2(n_1636),
.B(n_1652),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1718),
.Y(n_1825)
);

CKINVDCx14_ASAP7_75t_R g1826 ( 
.A(n_1736),
.Y(n_1826)
);

OAI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1582),
.A2(n_1666),
.B1(n_1769),
.B2(n_1644),
.Y(n_1827)
);

NOR2xp67_ASAP7_75t_SL g1828 ( 
.A(n_1768),
.B(n_1738),
.Y(n_1828)
);

NAND2x1p5_ASAP7_75t_L g1829 ( 
.A(n_1673),
.B(n_1648),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1642),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1602),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1575),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1575),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1709),
.B(n_1740),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1760),
.B(n_1762),
.Y(n_1835)
);

OAI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1636),
.A2(n_1652),
.B(n_1662),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1602),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1722),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1731),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1725),
.Y(n_1840)
);

OAI21x1_ASAP7_75t_L g1841 ( 
.A1(n_1647),
.A2(n_1641),
.B(n_1605),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1702),
.B(n_1639),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1771),
.B(n_1584),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1749),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1773),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1609),
.Y(n_1846)
);

OAI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1647),
.A2(n_1641),
.B(n_1597),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1635),
.B(n_1603),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1679),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1679),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1594),
.B(n_1595),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1700),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1588),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1603),
.B(n_1627),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1608),
.Y(n_1855)
);

AO31x2_ASAP7_75t_L g1856 ( 
.A1(n_1699),
.A2(n_1640),
.A3(n_1695),
.B(n_1625),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1770),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1609),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1618),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1577),
.A2(n_1733),
.B1(n_1732),
.B2(n_1729),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1623),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1606),
.Y(n_1862)
);

OR2x6_ASAP7_75t_L g1863 ( 
.A(n_1624),
.B(n_1620),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1629),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1630),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1607),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1609),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1708),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1607),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1651),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1735),
.Y(n_1871)
);

AOI21x1_ASAP7_75t_L g1872 ( 
.A1(n_1617),
.A2(n_1632),
.B(n_1657),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1651),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1671),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1600),
.B(n_1586),
.Y(n_1875)
);

OAI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1638),
.A2(n_1615),
.B(n_1600),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1589),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1601),
.Y(n_1878)
);

INVx4_ASAP7_75t_L g1879 ( 
.A(n_1708),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1621),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1577),
.A2(n_1755),
.B1(n_1706),
.B2(n_1729),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1716),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1727),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1706),
.A2(n_1755),
.B1(n_1732),
.B2(n_1764),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1586),
.B(n_1576),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1576),
.B(n_1615),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1708),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1720),
.B(n_1721),
.Y(n_1888)
);

INVx3_ASAP7_75t_SL g1889 ( 
.A(n_1730),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1747),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1633),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1720),
.B(n_1721),
.Y(n_1892)
);

BUFx3_ASAP7_75t_L g1893 ( 
.A(n_1650),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1659),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1682),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1613),
.B(n_1764),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1613),
.B(n_1733),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1590),
.A2(n_1739),
.B1(n_1756),
.B2(n_1763),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1730),
.Y(n_1899)
);

OAI21x1_ASAP7_75t_L g1900 ( 
.A1(n_1670),
.A2(n_1767),
.B(n_1683),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1680),
.Y(n_1901)
);

CKINVDCx6p67_ASAP7_75t_R g1902 ( 
.A(n_1754),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1680),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1616),
.A2(n_1689),
.B(n_1748),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1659),
.Y(n_1905)
);

AOI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1761),
.A2(n_1765),
.B1(n_1753),
.B2(n_1763),
.C(n_1756),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1659),
.B(n_1767),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1664),
.Y(n_1908)
);

OA21x2_ASAP7_75t_L g1909 ( 
.A1(n_1634),
.A2(n_1660),
.B(n_1723),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1660),
.Y(n_1910)
);

OAI21x1_ASAP7_75t_L g1911 ( 
.A1(n_1730),
.A2(n_1734),
.B(n_1660),
.Y(n_1911)
);

INVx3_ASAP7_75t_L g1912 ( 
.A(n_1734),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_R g1913 ( 
.A(n_1759),
.B(n_1766),
.Y(n_1913)
);

AOI21x1_ASAP7_75t_L g1914 ( 
.A1(n_1751),
.A2(n_1643),
.B(n_1661),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1734),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1574),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1574),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1579),
.Y(n_1918)
);

OAI21xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1649),
.A2(n_1658),
.B(n_1748),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1579),
.Y(n_1920)
);

OAI21x1_ASAP7_75t_L g1921 ( 
.A1(n_1645),
.A2(n_1748),
.B(n_1742),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1661),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1713),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1661),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1614),
.Y(n_1925)
);

INVx2_ASAP7_75t_SL g1926 ( 
.A(n_1713),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1614),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1645),
.A2(n_1746),
.B(n_1742),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1614),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1622),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1739),
.B(n_1637),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1622),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1611),
.Y(n_1933)
);

AO21x1_ASAP7_75t_L g1934 ( 
.A1(n_1637),
.A2(n_1645),
.B(n_1742),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1653),
.B(n_1611),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1596),
.B(n_1573),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1626),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1628),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1726),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1656),
.B(n_1741),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1581),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1581),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1758),
.B(n_1719),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1578),
.B(n_1619),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1743),
.A2(n_1750),
.B1(n_1592),
.B2(n_1772),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1592),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1772),
.B(n_1726),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1744),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1830),
.B(n_1784),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1902),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1796),
.A2(n_1799),
.B1(n_1881),
.B2(n_1860),
.C(n_1805),
.Y(n_1951)
);

NOR2x1_ASAP7_75t_SL g1952 ( 
.A(n_1863),
.B(n_1872),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1902),
.Y(n_1953)
);

AO32x2_ASAP7_75t_L g1954 ( 
.A1(n_1857),
.A2(n_1926),
.A3(n_1923),
.B1(n_1873),
.B2(n_1870),
.Y(n_1954)
);

O2A1O1Ixp33_ASAP7_75t_L g1955 ( 
.A1(n_1843),
.A2(n_1827),
.B(n_1892),
.C(n_1888),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1871),
.B(n_1831),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1893),
.Y(n_1957)
);

OAI22xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1799),
.A2(n_1884),
.B1(n_1835),
.B2(n_1818),
.Y(n_1958)
);

NAND3xp33_ASAP7_75t_L g1959 ( 
.A(n_1884),
.B(n_1885),
.C(n_1875),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1817),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1857),
.B(n_1781),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1854),
.B(n_1831),
.Y(n_1962)
);

A2O1A1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1876),
.A2(n_1851),
.B(n_1885),
.C(n_1836),
.Y(n_1963)
);

INVxp33_ASAP7_75t_SL g1964 ( 
.A(n_1913),
.Y(n_1964)
);

OR2x6_ASAP7_75t_L g1965 ( 
.A(n_1863),
.B(n_1900),
.Y(n_1965)
);

AOI22x1_ASAP7_75t_SL g1966 ( 
.A1(n_1948),
.A2(n_1814),
.B1(n_1874),
.B2(n_1938),
.Y(n_1966)
);

A2O1A1Ixp33_ASAP7_75t_L g1967 ( 
.A1(n_1876),
.A2(n_1836),
.B(n_1875),
.C(n_1896),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1871),
.B(n_1837),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1829),
.A2(n_1824),
.B(n_1841),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1886),
.A2(n_1897),
.B1(n_1896),
.B2(n_1873),
.C(n_1870),
.Y(n_1970)
);

AO21x2_ASAP7_75t_L g1971 ( 
.A1(n_1901),
.A2(n_1903),
.B(n_1806),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1818),
.A2(n_1863),
.B1(n_1826),
.B2(n_1898),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1909),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1943),
.Y(n_1974)
);

OA21x2_ASAP7_75t_L g1975 ( 
.A1(n_1795),
.A2(n_1806),
.B(n_1824),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1823),
.B(n_1874),
.Y(n_1976)
);

OAI211xp5_ASAP7_75t_L g1977 ( 
.A1(n_1897),
.A2(n_1886),
.B(n_1906),
.C(n_1919),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1848),
.B(n_1782),
.Y(n_1978)
);

A2O1A1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1904),
.A2(n_1841),
.B(n_1847),
.C(n_1919),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1914),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1845),
.B(n_1911),
.Y(n_1981)
);

O2A1O1Ixp33_ASAP7_75t_SL g1982 ( 
.A1(n_1814),
.A2(n_1948),
.B(n_1939),
.C(n_1933),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_SL g1983 ( 
.A1(n_1818),
.A2(n_1863),
.B1(n_1945),
.B2(n_1941),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1842),
.B(n_1815),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_SL g1985 ( 
.A1(n_1818),
.A2(n_1863),
.B1(n_1783),
.B2(n_1815),
.Y(n_1985)
);

O2A1O1Ixp33_ASAP7_75t_SL g1986 ( 
.A1(n_1814),
.A2(n_1910),
.B(n_1938),
.C(n_1937),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1807),
.B(n_1821),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1793),
.B(n_1819),
.Y(n_1988)
);

AND2x4_ASAP7_75t_L g1989 ( 
.A(n_1911),
.B(n_1797),
.Y(n_1989)
);

INVx6_ASAP7_75t_SL g1990 ( 
.A(n_1943),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1842),
.B(n_1848),
.Y(n_1991)
);

O2A1O1Ixp33_ASAP7_75t_SL g1992 ( 
.A1(n_1910),
.A2(n_1937),
.B(n_1942),
.C(n_1941),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1931),
.B(n_1909),
.Y(n_1993)
);

CKINVDCx20_ASAP7_75t_R g1994 ( 
.A(n_1944),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1931),
.B(n_1909),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1909),
.B(n_1818),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1819),
.B(n_1820),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1797),
.B(n_1802),
.Y(n_1998)
);

O2A1O1Ixp33_ASAP7_75t_SL g1999 ( 
.A1(n_1942),
.A2(n_1946),
.B(n_1936),
.C(n_1924),
.Y(n_1999)
);

OA21x2_ASAP7_75t_L g2000 ( 
.A1(n_1852),
.A2(n_1895),
.B(n_1810),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1864),
.B(n_1865),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1907),
.B(n_1893),
.Y(n_2002)
);

A2O1A1Ixp33_ASAP7_75t_L g2003 ( 
.A1(n_1783),
.A2(n_1850),
.B(n_1849),
.C(n_1828),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1787),
.A2(n_1829),
.B(n_1783),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1820),
.B(n_1822),
.Y(n_2005)
);

A2O1A1Ixp33_ASAP7_75t_L g2006 ( 
.A1(n_1850),
.A2(n_1828),
.B(n_1895),
.C(n_1946),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1935),
.B(n_1822),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1788),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1825),
.B(n_1838),
.Y(n_2009)
);

OAI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1829),
.A2(n_1794),
.B(n_1852),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1853),
.B(n_1855),
.Y(n_2011)
);

AO32x2_ASAP7_75t_L g2012 ( 
.A1(n_1798),
.A2(n_1879),
.A3(n_1794),
.B1(n_1809),
.B2(n_1856),
.Y(n_2012)
);

INVx4_ASAP7_75t_L g2013 ( 
.A(n_1889),
.Y(n_2013)
);

A2O1A1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_1788),
.A2(n_1832),
.B(n_1833),
.C(n_1846),
.Y(n_2014)
);

OAI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1776),
.A2(n_1804),
.B(n_1890),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1940),
.A2(n_1947),
.B1(n_1839),
.B2(n_1816),
.Y(n_2016)
);

BUFx2_ASAP7_75t_L g2017 ( 
.A(n_1788),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1840),
.B(n_1844),
.Y(n_2018)
);

INVx3_ASAP7_75t_SL g2019 ( 
.A(n_1940),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1889),
.A2(n_1798),
.B1(n_1879),
.B2(n_1844),
.Y(n_2020)
);

AOI221xp5_ASAP7_75t_L g2021 ( 
.A1(n_1859),
.A2(n_1861),
.B1(n_1891),
.B2(n_1862),
.C(n_1787),
.Y(n_2021)
);

OAI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1914),
.A2(n_1891),
.B(n_1834),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1940),
.A2(n_1947),
.B1(n_1868),
.B2(n_1867),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_1889),
.A2(n_1798),
.B1(n_1879),
.B2(n_1859),
.Y(n_2024)
);

A2O1A1Ixp33_ASAP7_75t_L g2025 ( 
.A1(n_1832),
.A2(n_1833),
.B(n_1912),
.C(n_1846),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1834),
.B(n_1905),
.Y(n_2026)
);

A2O1A1Ixp33_ASAP7_75t_L g2027 ( 
.A1(n_1832),
.A2(n_1868),
.B(n_1846),
.C(n_1867),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1790),
.Y(n_2028)
);

AO21x1_ASAP7_75t_L g2029 ( 
.A1(n_1862),
.A2(n_1812),
.B(n_1916),
.Y(n_2029)
);

O2A1O1Ixp33_ASAP7_75t_SL g2030 ( 
.A1(n_1924),
.A2(n_1925),
.B(n_1927),
.C(n_1833),
.Y(n_2030)
);

NAND2x1p5_ASAP7_75t_L g2031 ( 
.A(n_1800),
.B(n_1879),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1834),
.B(n_1894),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1789),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1798),
.A2(n_1912),
.B1(n_1867),
.B2(n_1868),
.Y(n_2034)
);

AO21x2_ASAP7_75t_L g2035 ( 
.A1(n_1787),
.A2(n_1774),
.B(n_1775),
.Y(n_2035)
);

OR2x2_ASAP7_75t_L g2036 ( 
.A(n_1791),
.B(n_1792),
.Y(n_2036)
);

A2O1A1Ixp33_ASAP7_75t_L g2037 ( 
.A1(n_1899),
.A2(n_1912),
.B(n_1803),
.C(n_1915),
.Y(n_2037)
);

AO32x2_ASAP7_75t_L g2038 ( 
.A1(n_1856),
.A2(n_1800),
.A3(n_1791),
.B1(n_1792),
.B2(n_1778),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1774),
.Y(n_2039)
);

OAI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_1834),
.A2(n_1880),
.B(n_1877),
.Y(n_2040)
);

OAI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1899),
.A2(n_1858),
.B1(n_1813),
.B2(n_1887),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1917),
.B(n_1918),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1940),
.A2(n_1943),
.B1(n_1915),
.B2(n_1922),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1866),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1775),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_1777),
.B(n_1779),
.Y(n_2046)
);

AND2x4_ASAP7_75t_SL g2047 ( 
.A(n_1943),
.B(n_1858),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1866),
.B(n_1869),
.Y(n_2048)
);

AND2x2_ASAP7_75t_SL g2049 ( 
.A(n_2021),
.B(n_1800),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1993),
.B(n_1995),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_1951),
.A2(n_1800),
.B1(n_1908),
.B2(n_1858),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_2028),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2033),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_SL g2054 ( 
.A(n_1965),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1978),
.B(n_1786),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_1951),
.A2(n_1858),
.B1(n_1887),
.B2(n_1813),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1991),
.B(n_1856),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2039),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_1981),
.B(n_1786),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1950),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1981),
.B(n_1786),
.Y(n_2061)
);

BUFx2_ASAP7_75t_SL g2062 ( 
.A(n_2029),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1989),
.B(n_1786),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2045),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1984),
.B(n_1856),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2048),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2048),
.Y(n_2067)
);

BUFx2_ASAP7_75t_L g2068 ( 
.A(n_1954),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1958),
.A2(n_1887),
.B1(n_1813),
.B2(n_1858),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1960),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1962),
.B(n_1856),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1949),
.B(n_1786),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1978),
.B(n_1780),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_2019),
.B(n_1913),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2007),
.B(n_1883),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_1959),
.A2(n_1887),
.B1(n_1813),
.B2(n_1922),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_1961),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2046),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2011),
.Y(n_2079)
);

OR2x6_ASAP7_75t_L g2080 ( 
.A(n_1965),
.B(n_1785),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1998),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_1987),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1996),
.B(n_2026),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1959),
.B(n_1877),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2032),
.B(n_2018),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2036),
.Y(n_2086)
);

AND2x4_ASAP7_75t_SL g2087 ( 
.A(n_2013),
.B(n_1887),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1957),
.B(n_1932),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1970),
.B(n_1878),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1977),
.A2(n_1908),
.B1(n_1932),
.B2(n_1930),
.Y(n_2090)
);

INVxp67_ASAP7_75t_SL g2091 ( 
.A(n_2044),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2035),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1970),
.B(n_1882),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1997),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2012),
.B(n_1811),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1972),
.A2(n_1930),
.B1(n_1929),
.B2(n_1882),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1954),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2012),
.B(n_1801),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2005),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_1988),
.Y(n_2100)
);

AND2x4_ASAP7_75t_SL g2101 ( 
.A(n_1956),
.B(n_1808),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_1973),
.B(n_1869),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1969),
.B(n_1920),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2009),
.Y(n_2104)
);

AOI33xp33_ASAP7_75t_L g2105 ( 
.A1(n_2057),
.A2(n_1955),
.A3(n_1985),
.B1(n_2021),
.B2(n_2043),
.B3(n_1982),
.Y(n_2105)
);

BUFx2_ASAP7_75t_L g2106 ( 
.A(n_2059),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2052),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_2084),
.B(n_1974),
.Y(n_2108)
);

BUFx3_ASAP7_75t_L g2109 ( 
.A(n_2087),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2050),
.B(n_1973),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2050),
.B(n_1954),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_2074),
.B(n_2023),
.Y(n_2112)
);

AOI211xp5_ASAP7_75t_L g2113 ( 
.A1(n_2051),
.A2(n_1977),
.B(n_1983),
.C(n_1963),
.Y(n_2113)
);

INVxp67_ASAP7_75t_L g2114 ( 
.A(n_2100),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_2082),
.B(n_1964),
.Y(n_2115)
);

NAND3xp33_ASAP7_75t_L g2116 ( 
.A(n_2090),
.B(n_2006),
.C(n_1967),
.Y(n_2116)
);

OAI221xp5_ASAP7_75t_L g2117 ( 
.A1(n_2069),
.A2(n_1979),
.B1(n_2016),
.B2(n_2015),
.C(n_2004),
.Y(n_2117)
);

INVx5_ASAP7_75t_L g2118 ( 
.A(n_2080),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2083),
.B(n_1971),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2098),
.Y(n_2120)
);

NOR2x1_ASAP7_75t_L g2121 ( 
.A(n_2062),
.B(n_1980),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2098),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2064),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2083),
.B(n_2072),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2055),
.B(n_2000),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2072),
.B(n_1971),
.Y(n_2126)
);

NAND3xp33_ASAP7_75t_L g2127 ( 
.A(n_2090),
.B(n_2010),
.C(n_2003),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_2051),
.B(n_1953),
.Y(n_2128)
);

AO21x2_ASAP7_75t_L g2129 ( 
.A1(n_2092),
.A2(n_2010),
.B(n_2004),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_2077),
.Y(n_2130)
);

AOI211xp5_ASAP7_75t_L g2131 ( 
.A1(n_2065),
.A2(n_2020),
.B(n_2024),
.C(n_2015),
.Y(n_2131)
);

INVx4_ASAP7_75t_L g2132 ( 
.A(n_2087),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2085),
.B(n_1976),
.Y(n_2133)
);

NAND3xp33_ASAP7_75t_L g2134 ( 
.A(n_2056),
.B(n_1999),
.C(n_2014),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2102),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_2059),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2085),
.B(n_2038),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2102),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2057),
.B(n_2038),
.Y(n_2139)
);

INVx5_ASAP7_75t_L g2140 ( 
.A(n_2080),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2053),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2053),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2095),
.Y(n_2143)
);

INVx1_ASAP7_75t_SL g2144 ( 
.A(n_2101),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2058),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_2059),
.B(n_1952),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_2073),
.Y(n_2147)
);

AOI33xp33_ASAP7_75t_L g2148 ( 
.A1(n_2065),
.A2(n_1992),
.A3(n_1986),
.B1(n_2002),
.B2(n_2047),
.B3(n_2042),
.Y(n_2148)
);

OAI33xp33_ASAP7_75t_L g2149 ( 
.A1(n_2055),
.A2(n_2024),
.A3(n_2020),
.B1(n_2034),
.B2(n_2001),
.B3(n_2041),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2066),
.B(n_2038),
.Y(n_2150)
);

INVx4_ASAP7_75t_L g2151 ( 
.A(n_2087),
.Y(n_2151)
);

OR2x2_ASAP7_75t_L g2152 ( 
.A(n_2073),
.B(n_2000),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2095),
.Y(n_2153)
);

AOI211xp5_ASAP7_75t_L g2154 ( 
.A1(n_2089),
.A2(n_2034),
.B(n_2041),
.C(n_2025),
.Y(n_2154)
);

NAND4xp25_ASAP7_75t_L g2155 ( 
.A(n_2093),
.B(n_2027),
.C(n_2022),
.D(n_2037),
.Y(n_2155)
);

OAI211xp5_ASAP7_75t_L g2156 ( 
.A1(n_2068),
.A2(n_2022),
.B(n_1975),
.C(n_2040),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2066),
.B(n_1968),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2058),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2066),
.B(n_1968),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2070),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2126),
.B(n_2078),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2106),
.B(n_2068),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2126),
.B(n_2078),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2106),
.B(n_2097),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2141),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2123),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2136),
.B(n_2097),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2111),
.B(n_2094),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2111),
.B(n_2094),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2123),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2141),
.B(n_2099),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2125),
.B(n_2067),
.Y(n_2172)
);

NOR2x2_ASAP7_75t_L g2173 ( 
.A(n_2120),
.B(n_1966),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2136),
.B(n_2080),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2142),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2142),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2137),
.B(n_2080),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2145),
.B(n_2104),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2158),
.B(n_2104),
.Y(n_2179)
);

INVx4_ASAP7_75t_L g2180 ( 
.A(n_2132),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_2146),
.B(n_2061),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2137),
.B(n_2080),
.Y(n_2182)
);

INVxp33_ASAP7_75t_SL g2183 ( 
.A(n_2115),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2158),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2160),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2160),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2124),
.B(n_2081),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2125),
.B(n_2081),
.Y(n_2188)
);

INVxp67_ASAP7_75t_L g2189 ( 
.A(n_2130),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2147),
.B(n_2086),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2124),
.B(n_2081),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2123),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2139),
.B(n_2135),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2139),
.B(n_2086),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2135),
.B(n_2079),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_2112),
.B(n_2008),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2119),
.B(n_2061),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_2152),
.B(n_2091),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2138),
.B(n_2079),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2107),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2119),
.B(n_2061),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2110),
.B(n_2146),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2110),
.B(n_2061),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2146),
.B(n_2063),
.Y(n_2204)
);

INVx1_ASAP7_75t_SL g2205 ( 
.A(n_2144),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2152),
.B(n_2075),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_2146),
.B(n_2063),
.Y(n_2207)
);

OR2x2_ASAP7_75t_L g2208 ( 
.A(n_2138),
.B(n_2062),
.Y(n_2208)
);

OAI21xp5_ASAP7_75t_L g2209 ( 
.A1(n_2116),
.A2(n_2049),
.B(n_2096),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2165),
.Y(n_2210)
);

OR2x2_ASAP7_75t_L g2211 ( 
.A(n_2193),
.B(n_2156),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2202),
.B(n_2120),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_2181),
.B(n_2118),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2166),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2166),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2166),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2183),
.B(n_2060),
.Y(n_2217)
);

NOR2x1_ASAP7_75t_L g2218 ( 
.A(n_2180),
.B(n_2121),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2202),
.B(n_2181),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2181),
.B(n_2120),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2181),
.B(n_2122),
.Y(n_2221)
);

AOI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2209),
.A2(n_2116),
.B1(n_2113),
.B2(n_2127),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2170),
.Y(n_2223)
);

OAI21xp33_ASAP7_75t_L g2224 ( 
.A1(n_2209),
.A2(n_2105),
.B(n_2127),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2170),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2196),
.B(n_2114),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2165),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2175),
.Y(n_2228)
);

OAI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_2196),
.A2(n_2113),
.B1(n_2117),
.B2(n_2134),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_2180),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2193),
.B(n_2143),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2207),
.B(n_2122),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2175),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2207),
.B(n_2122),
.Y(n_2234)
);

NAND2xp67_ASAP7_75t_SL g2235 ( 
.A(n_2162),
.B(n_2103),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2161),
.B(n_2143),
.Y(n_2236)
);

OR2x2_ASAP7_75t_L g2237 ( 
.A(n_2161),
.B(n_2143),
.Y(n_2237)
);

INVxp67_ASAP7_75t_L g2238 ( 
.A(n_2189),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2176),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_2189),
.B(n_2148),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2163),
.B(n_2153),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2190),
.B(n_2154),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2176),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2170),
.Y(n_2244)
);

NAND2x1_ASAP7_75t_L g2245 ( 
.A(n_2180),
.B(n_2121),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2184),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2207),
.B(n_2157),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2184),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_2163),
.B(n_2153),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2207),
.B(n_2157),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2177),
.B(n_2182),
.Y(n_2251)
);

OAI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_2208),
.A2(n_2134),
.B(n_2128),
.Y(n_2252)
);

AND2x2_ASAP7_75t_SL g2253 ( 
.A(n_2180),
.B(n_2049),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2208),
.B(n_2153),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2192),
.Y(n_2255)
);

INVx2_ASAP7_75t_SL g2256 ( 
.A(n_2174),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2185),
.Y(n_2257)
);

INVx1_ASAP7_75t_SL g2258 ( 
.A(n_2173),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2177),
.B(n_2159),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2192),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2185),
.Y(n_2261)
);

AOI32xp33_ASAP7_75t_L g2262 ( 
.A1(n_2162),
.A2(n_2131),
.A3(n_2154),
.B1(n_2071),
.B2(n_2076),
.Y(n_2262)
);

NOR2xp33_ASAP7_75t_L g2263 ( 
.A(n_2205),
.B(n_2155),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2182),
.B(n_2159),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2192),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_2205),
.B(n_2131),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2251),
.B(n_2204),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2210),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2210),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2238),
.B(n_2194),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2251),
.B(n_2204),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2222),
.B(n_2187),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2219),
.B(n_2259),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2222),
.B(n_2187),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2224),
.A2(n_2229),
.B1(n_2258),
.B2(n_2266),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_2218),
.B(n_2219),
.Y(n_2276)
);

OR2x2_ASAP7_75t_L g2277 ( 
.A(n_2211),
.B(n_2194),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2224),
.B(n_2191),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2211),
.B(n_2198),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2227),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2259),
.B(n_2162),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2227),
.Y(n_2282)
);

BUFx2_ASAP7_75t_L g2283 ( 
.A(n_2218),
.Y(n_2283)
);

A2O1A1Ixp33_ASAP7_75t_L g2284 ( 
.A1(n_2262),
.A2(n_2155),
.B(n_2049),
.C(n_2108),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2263),
.B(n_2191),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_2242),
.B(n_2198),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2230),
.B(n_2164),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2228),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2220),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2228),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2264),
.B(n_2197),
.Y(n_2291)
);

NOR3xp33_ASAP7_75t_L g2292 ( 
.A(n_2252),
.B(n_2149),
.C(n_2017),
.Y(n_2292)
);

NAND2x1_ASAP7_75t_L g2293 ( 
.A(n_2213),
.B(n_2164),
.Y(n_2293)
);

NOR2x1_ASAP7_75t_L g2294 ( 
.A(n_2230),
.B(n_2186),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_L g2295 ( 
.A(n_2217),
.B(n_1994),
.Y(n_2295)
);

INVx2_ASAP7_75t_SL g2296 ( 
.A(n_2245),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2240),
.B(n_2190),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2262),
.B(n_2133),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2226),
.B(n_2133),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_2230),
.B(n_2167),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2264),
.B(n_2197),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2247),
.B(n_2250),
.Y(n_2302)
);

OR2x2_ASAP7_75t_L g2303 ( 
.A(n_2256),
.B(n_2168),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2256),
.B(n_2168),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2247),
.B(n_2169),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2250),
.B(n_2201),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2213),
.B(n_2201),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2212),
.B(n_2169),
.Y(n_2308)
);

INVx2_ASAP7_75t_SL g2309 ( 
.A(n_2245),
.Y(n_2309)
);

OAI211xp5_ASAP7_75t_SL g2310 ( 
.A1(n_2275),
.A2(n_2230),
.B(n_2225),
.C(n_2260),
.Y(n_2310)
);

NOR2xp33_ASAP7_75t_L g2311 ( 
.A(n_2295),
.B(n_2213),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2268),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2278),
.B(n_2233),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2297),
.B(n_2212),
.Y(n_2314)
);

AOI211xp5_ASAP7_75t_L g2315 ( 
.A1(n_2284),
.A2(n_2213),
.B(n_2261),
.C(n_2233),
.Y(n_2315)
);

NAND3xp33_ASAP7_75t_L g2316 ( 
.A(n_2284),
.B(n_2253),
.C(n_2243),
.Y(n_2316)
);

NAND2xp33_ASAP7_75t_L g2317 ( 
.A(n_2292),
.B(n_2118),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2272),
.B(n_2274),
.Y(n_2318)
);

AND2x4_ASAP7_75t_L g2319 ( 
.A(n_2276),
.B(n_2220),
.Y(n_2319)
);

AOI211xp5_ASAP7_75t_L g2320 ( 
.A1(n_2298),
.A2(n_2239),
.B(n_2261),
.C(n_2243),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2286),
.B(n_2239),
.Y(n_2321)
);

OAI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2283),
.A2(n_2253),
.B(n_2167),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2299),
.B(n_2206),
.Y(n_2323)
);

OAI21xp5_ASAP7_75t_SL g2324 ( 
.A1(n_2283),
.A2(n_2253),
.B(n_2232),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2273),
.Y(n_2325)
);

AOI21xp33_ASAP7_75t_L g2326 ( 
.A1(n_2286),
.A2(n_2129),
.B(n_2246),
.Y(n_2326)
);

OAI21xp33_ASAP7_75t_L g2327 ( 
.A1(n_2285),
.A2(n_2232),
.B(n_2221),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2273),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2302),
.Y(n_2329)
);

OAI21xp33_ASAP7_75t_L g2330 ( 
.A1(n_2270),
.A2(n_2221),
.B(n_2234),
.Y(n_2330)
);

AOI32xp33_ASAP7_75t_L g2331 ( 
.A1(n_2276),
.A2(n_2234),
.A3(n_2174),
.B1(n_2235),
.B2(n_2254),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_L g2332 ( 
.A1(n_2307),
.A2(n_2054),
.B1(n_2129),
.B2(n_2140),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2269),
.Y(n_2333)
);

OR2x2_ASAP7_75t_L g2334 ( 
.A(n_2279),
.B(n_2254),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2280),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2282),
.Y(n_2336)
);

OAI221xp5_ASAP7_75t_L g2337 ( 
.A1(n_2293),
.A2(n_2231),
.B1(n_2246),
.B2(n_2257),
.C(n_2248),
.Y(n_2337)
);

OR2x2_ASAP7_75t_L g2338 ( 
.A(n_2279),
.B(n_2231),
.Y(n_2338)
);

AOI32xp33_ASAP7_75t_L g2339 ( 
.A1(n_2276),
.A2(n_2235),
.A3(n_2144),
.B1(n_2071),
.B2(n_2248),
.Y(n_2339)
);

INVx1_ASAP7_75t_SL g2340 ( 
.A(n_2334),
.Y(n_2340)
);

NAND3xp33_ASAP7_75t_L g2341 ( 
.A(n_2315),
.B(n_2294),
.C(n_2270),
.Y(n_2341)
);

NOR2x1_ASAP7_75t_L g2342 ( 
.A(n_2316),
.B(n_2288),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2325),
.B(n_2302),
.Y(n_2343)
);

OAI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2318),
.A2(n_2309),
.B1(n_2296),
.B2(n_2277),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2328),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2329),
.B(n_2281),
.Y(n_2346)
);

HB1xp67_ASAP7_75t_L g2347 ( 
.A(n_2338),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2312),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2319),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2333),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2320),
.B(n_2281),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_2322),
.B(n_2296),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2314),
.B(n_2267),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2322),
.A2(n_2324),
.B1(n_2311),
.B2(n_2309),
.Y(n_2354)
);

OAI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_2339),
.A2(n_2277),
.B1(n_2271),
.B2(n_2267),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2319),
.B(n_2271),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2313),
.B(n_2291),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2337),
.A2(n_2305),
.B1(n_2291),
.B2(n_2301),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2335),
.Y(n_2359)
);

INVxp67_ASAP7_75t_L g2360 ( 
.A(n_2313),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2336),
.Y(n_2361)
);

A2O1A1Ixp33_ASAP7_75t_L g2362 ( 
.A1(n_2342),
.A2(n_2331),
.B(n_2317),
.C(n_2310),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2347),
.Y(n_2363)
);

AOI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2354),
.A2(n_2330),
.B1(n_2327),
.B2(n_2300),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2347),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2346),
.Y(n_2366)
);

AOI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2352),
.A2(n_2321),
.B(n_2326),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2340),
.B(n_2321),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2345),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2343),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2349),
.Y(n_2371)
);

AOI21xp33_ASAP7_75t_L g2372 ( 
.A1(n_2352),
.A2(n_2323),
.B(n_2300),
.Y(n_2372)
);

INVx1_ASAP7_75t_SL g2373 ( 
.A(n_2349),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2356),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2356),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2373),
.B(n_2374),
.Y(n_2376)
);

OA22x2_ASAP7_75t_L g2377 ( 
.A1(n_2373),
.A2(n_2360),
.B1(n_2344),
.B2(n_2351),
.Y(n_2377)
);

INVx1_ASAP7_75t_SL g2378 ( 
.A(n_2363),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2365),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2375),
.Y(n_2380)
);

NOR3xp33_ASAP7_75t_L g2381 ( 
.A(n_2370),
.B(n_2341),
.C(n_2348),
.Y(n_2381)
);

OAI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2362),
.A2(n_2367),
.B(n_2372),
.Y(n_2382)
);

NOR3xp33_ASAP7_75t_SL g2383 ( 
.A(n_2366),
.B(n_2358),
.C(n_2355),
.Y(n_2383)
);

INVxp67_ASAP7_75t_SL g2384 ( 
.A(n_2368),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2371),
.B(n_2353),
.Y(n_2385)
);

NAND3xp33_ASAP7_75t_SL g2386 ( 
.A(n_2364),
.B(n_2357),
.C(n_2350),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2369),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2363),
.Y(n_2388)
);

AND4x1_ASAP7_75t_L g2389 ( 
.A(n_2382),
.B(n_2383),
.C(n_2376),
.D(n_2381),
.Y(n_2389)
);

OAI32xp33_ASAP7_75t_L g2390 ( 
.A1(n_2378),
.A2(n_2361),
.A3(n_2359),
.B1(n_2326),
.B2(n_2303),
.Y(n_2390)
);

AOI221xp5_ASAP7_75t_L g2391 ( 
.A1(n_2386),
.A2(n_2332),
.B1(n_2290),
.B2(n_2287),
.C(n_2300),
.Y(n_2391)
);

INVxp67_ASAP7_75t_L g2392 ( 
.A(n_2384),
.Y(n_2392)
);

OAI211xp5_ASAP7_75t_L g2393 ( 
.A1(n_2378),
.A2(n_2289),
.B(n_2307),
.C(n_2304),
.Y(n_2393)
);

AOI221xp5_ASAP7_75t_L g2394 ( 
.A1(n_2388),
.A2(n_2287),
.B1(n_2289),
.B2(n_2303),
.C(n_2308),
.Y(n_2394)
);

OAI21xp33_ASAP7_75t_L g2395 ( 
.A1(n_2377),
.A2(n_2287),
.B(n_2306),
.Y(n_2395)
);

AOI321xp33_ASAP7_75t_L g2396 ( 
.A1(n_2385),
.A2(n_2306),
.A3(n_2301),
.B1(n_2225),
.B2(n_2260),
.C(n_2255),
.Y(n_2396)
);

AOI211xp5_ASAP7_75t_L g2397 ( 
.A1(n_2380),
.A2(n_2379),
.B(n_2387),
.C(n_2377),
.Y(n_2397)
);

OAI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2382),
.A2(n_2257),
.B1(n_2237),
.B2(n_2236),
.Y(n_2398)
);

OAI211xp5_ASAP7_75t_SL g2399 ( 
.A1(n_2392),
.A2(n_2225),
.B(n_2260),
.C(n_2255),
.Y(n_2399)
);

AOI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2390),
.A2(n_2255),
.B1(n_2265),
.B2(n_2244),
.C(n_2223),
.Y(n_2400)
);

AOI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2397),
.A2(n_2395),
.B(n_2391),
.Y(n_2401)
);

NOR3xp33_ASAP7_75t_L g2402 ( 
.A(n_2393),
.B(n_2265),
.C(n_2215),
.Y(n_2402)
);

NAND3x1_ASAP7_75t_SL g2403 ( 
.A(n_2394),
.B(n_1990),
.C(n_2150),
.Y(n_2403)
);

NAND4xp25_ASAP7_75t_L g2404 ( 
.A(n_2396),
.B(n_2088),
.C(n_2132),
.D(n_2151),
.Y(n_2404)
);

OAI221xp5_ASAP7_75t_L g2405 ( 
.A1(n_2389),
.A2(n_2214),
.B1(n_2244),
.B2(n_2215),
.C(n_2216),
.Y(n_2405)
);

HB1xp67_ASAP7_75t_L g2406 ( 
.A(n_2398),
.Y(n_2406)
);

OAI322xp33_ASAP7_75t_L g2407 ( 
.A1(n_2392),
.A2(n_2214),
.A3(n_2223),
.B1(n_2216),
.B2(n_2249),
.C1(n_2236),
.C2(n_2241),
.Y(n_2407)
);

NOR2xp67_ASAP7_75t_L g2408 ( 
.A(n_2404),
.B(n_2237),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2406),
.Y(n_2409)
);

NOR2x1_ASAP7_75t_L g2410 ( 
.A(n_2401),
.B(n_2241),
.Y(n_2410)
);

INVx2_ASAP7_75t_SL g2411 ( 
.A(n_2403),
.Y(n_2411)
);

NAND4xp75_ASAP7_75t_L g2412 ( 
.A(n_2400),
.B(n_1934),
.C(n_2195),
.D(n_2199),
.Y(n_2412)
);

NAND4xp75_ASAP7_75t_L g2413 ( 
.A(n_2405),
.B(n_1934),
.C(n_2195),
.D(n_2199),
.Y(n_2413)
);

AND3x4_ASAP7_75t_L g2414 ( 
.A(n_2402),
.B(n_2109),
.C(n_1990),
.Y(n_2414)
);

AOI21xp33_ASAP7_75t_SL g2415 ( 
.A1(n_2409),
.A2(n_2399),
.B(n_2407),
.Y(n_2415)
);

XNOR2xp5_ASAP7_75t_L g2416 ( 
.A(n_2410),
.B(n_2031),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2414),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2408),
.B(n_2249),
.Y(n_2418)
);

NOR3xp33_ASAP7_75t_L g2419 ( 
.A(n_2417),
.B(n_2411),
.C(n_2413),
.Y(n_2419)
);

OAI22xp5_ASAP7_75t_L g2420 ( 
.A1(n_2418),
.A2(n_2412),
.B1(n_2172),
.B2(n_2188),
.Y(n_2420)
);

OAI22x1_ASAP7_75t_L g2421 ( 
.A1(n_2419),
.A2(n_2416),
.B1(n_2415),
.B2(n_2132),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2421),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2421),
.Y(n_2423)
);

OAI22x1_ASAP7_75t_L g2424 ( 
.A1(n_2422),
.A2(n_2420),
.B1(n_2132),
.B2(n_2151),
.Y(n_2424)
);

AOI22xp33_ASAP7_75t_SL g2425 ( 
.A1(n_2423),
.A2(n_2118),
.B1(n_2140),
.B2(n_2151),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2424),
.B(n_2203),
.Y(n_2426)
);

OAI21x1_ASAP7_75t_L g2427 ( 
.A1(n_2425),
.A2(n_2200),
.B(n_2186),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2426),
.B(n_2200),
.Y(n_2428)
);

AOI22xp33_ASAP7_75t_L g2429 ( 
.A1(n_2428),
.A2(n_2427),
.B1(n_2151),
.B2(n_2109),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_2429),
.Y(n_2430)
);

OAI221xp5_ASAP7_75t_R g2431 ( 
.A1(n_2430),
.A2(n_2427),
.B1(n_2179),
.B2(n_2178),
.C(n_2171),
.Y(n_2431)
);

AOI211xp5_ASAP7_75t_L g2432 ( 
.A1(n_2431),
.A2(n_1928),
.B(n_1921),
.C(n_2030),
.Y(n_2432)
);


endmodule