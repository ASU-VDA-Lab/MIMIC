module fake_jpeg_1037_n_229 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_229);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_15),
.B(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_21),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_27),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_5),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_6),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_84),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_79),
.Y(n_89)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_45),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_55),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_52),
.B1(n_72),
.B2(n_73),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_76),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_73),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_102),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_108),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_77),
.B1(n_56),
.B2(n_54),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_106),
.B1(n_86),
.B2(n_89),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_77),
.B1(n_56),
.B2(n_54),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_65),
.B(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_115),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_82),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_82),
.B1(n_65),
.B2(n_67),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_119),
.B1(n_73),
.B2(n_49),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_52),
.B1(n_72),
.B2(n_61),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_96),
.A3(n_85),
.B1(n_62),
.B2(n_71),
.Y(n_131)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_74),
.B1(n_70),
.B2(n_61),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_69),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_126),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_115),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_86),
.B1(n_85),
.B2(n_95),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_135),
.B1(n_139),
.B2(n_68),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_66),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_115),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_50),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_138),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_83),
.B1(n_58),
.B2(n_53),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_59),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_83),
.B1(n_58),
.B2(n_53),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_116),
.B1(n_118),
.B2(n_117),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_142),
.Y(n_186)
);

OAI21x1_ASAP7_75t_SL g168 ( 
.A1(n_145),
.A2(n_154),
.B(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_151),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_71),
.B1(n_62),
.B2(n_41),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_150),
.B1(n_155),
.B2(n_159),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_2),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_33),
.C(n_32),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_26),
.Y(n_174)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_3),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_164),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_5),
.B(n_7),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_14),
.B(n_16),
.Y(n_175)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_163),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_175),
.Y(n_195)
);

BUFx12f_ASAP7_75t_SL g197 ( 
.A(n_168),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_139),
.B(n_135),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_170),
.B(n_173),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_12),
.B(n_13),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_12),
.B(n_13),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_178),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_145),
.B(n_148),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_25),
.B(n_24),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_20),
.B(n_21),
.Y(n_196)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_141),
.B1(n_155),
.B2(n_156),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_200),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_181),
.A2(n_159),
.B1(n_16),
.B2(n_17),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_179),
.B1(n_184),
.B2(n_183),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_191),
.A2(n_198),
.B1(n_183),
.B2(n_184),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_18),
.C(n_19),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_199),
.C(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_172),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_22),
.B1(n_169),
.B2(n_185),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_180),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_171),
.C(n_170),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_173),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_209),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_205),
.B1(n_198),
.B2(n_197),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_207),
.Y(n_214)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_174),
.B(n_195),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_192),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_210),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_201),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_216),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_210),
.C(n_204),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_221),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_214),
.C(n_217),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_220),
.C(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_227),
.B(n_211),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_196),
.Y(n_229)
);


endmodule