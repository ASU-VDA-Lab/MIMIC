module fake_jpeg_30867_n_234 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.C(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_57),
.Y(n_73)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_47),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx6p67_ASAP7_75t_R g90 ( 
.A(n_44),
.Y(n_90)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_8),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_22),
.B(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_58),
.Y(n_80)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_2),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_36),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_11),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_27),
.Y(n_81)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_62),
.Y(n_94)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_36),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_88),
.C(n_6),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_75),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_67),
.B(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_91),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_31),
.B1(n_21),
.B2(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_32),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_21),
.B1(n_30),
.B2(n_24),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_21),
.B1(n_30),
.B2(n_24),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_95),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_34),
.B1(n_33),
.B2(n_38),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_50),
.B1(n_40),
.B2(n_7),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_30),
.B1(n_34),
.B2(n_38),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_37),
.B1(n_25),
.B2(n_20),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_37),
.B(n_25),
.C(n_20),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_50),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_11),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_100),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_122),
.B1(n_90),
.B2(n_65),
.Y(n_129)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_12),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_12),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_113),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_121),
.Y(n_133)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_120),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_6),
.B1(n_7),
.B2(n_14),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_63),
.B1(n_94),
.B2(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_15),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_15),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_64),
.B1(n_89),
.B2(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_78),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_116),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_144),
.B1(n_103),
.B2(n_109),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_125),
.A2(n_108),
.B1(n_112),
.B2(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_146),
.B1(n_117),
.B2(n_119),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_94),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_94),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_96),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_84),
.B1(n_65),
.B2(n_70),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_70),
.B1(n_83),
.B2(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_83),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_147),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_149),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_97),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_113),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_157),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_110),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_107),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_170),
.B1(n_141),
.B2(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_168),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_169),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_136),
.C(n_143),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_129),
.C(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_102),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_157),
.B(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_159),
.A2(n_146),
.B1(n_128),
.B2(n_130),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_186),
.B1(n_126),
.B2(n_164),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_169),
.A2(n_145),
.B(n_130),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_168),
.B(n_153),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_136),
.B(n_144),
.C(n_134),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_161),
.B(n_166),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_167),
.C(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_191),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_199),
.C(n_181),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_197),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_194),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_170),
.B1(n_151),
.B2(n_158),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_196),
.B(n_185),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_162),
.B1(n_155),
.B2(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_163),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_198),
.A2(n_183),
.B1(n_185),
.B2(n_182),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_139),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_205),
.B1(n_207),
.B2(n_199),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_193),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_175),
.B1(n_172),
.B2(n_184),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_171),
.A3(n_187),
.B1(n_179),
.B2(n_180),
.C1(n_176),
.C2(n_100),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_210),
.Y(n_215)
);

AOI31xp33_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_179),
.A3(n_180),
.B(n_115),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_196),
.B(n_191),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_189),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_197),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_203),
.C(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_220),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_207),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_202),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_204),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_226),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_208),
.B1(n_192),
.B2(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_227),
.B(n_222),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_230),
.C(n_208),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_225),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_224),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_232),
.C(n_223),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_233),
.Y(n_234)
);


endmodule