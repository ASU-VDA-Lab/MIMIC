module real_aes_8214_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g439 ( .A(n_0), .Y(n_439) );
INVx1_ASAP7_75t_L g504 ( .A(n_1), .Y(n_504) );
INVx1_ASAP7_75t_L g185 ( .A(n_2), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_3), .A2(n_37), .B1(n_157), .B2(n_513), .Y(n_512) );
AOI21xp33_ASAP7_75t_L g196 ( .A1(n_4), .A2(n_114), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_5), .B(n_144), .Y(n_496) );
AND2x6_ASAP7_75t_L g119 ( .A(n_6), .B(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_7), .A2(n_165), .B(n_166), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_8), .B(n_38), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_9), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g202 ( .A(n_10), .Y(n_202) );
INVx1_ASAP7_75t_L g140 ( .A(n_11), .Y(n_140) );
INVx1_ASAP7_75t_L g500 ( .A(n_12), .Y(n_500) );
INVx1_ASAP7_75t_L g173 ( .A(n_13), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_14), .B(n_188), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_15), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_16), .B(n_136), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_17), .A2(n_41), .B1(n_745), .B2(n_746), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_17), .Y(n_746) );
AO32x2_ASAP7_75t_L g510 ( .A1(n_18), .A2(n_135), .A3(n_144), .B1(n_482), .B2(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_19), .B(n_157), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_20), .B(n_130), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_21), .B(n_136), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_22), .A2(n_49), .B1(n_157), .B2(n_513), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_23), .B(n_114), .Y(n_113) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_24), .A2(n_75), .B1(n_157), .B2(n_188), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_25), .B(n_157), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_26), .B(n_195), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_27), .A2(n_170), .B(n_172), .C(n_174), .Y(n_169) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_28), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_29), .B(n_148), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_30), .B(n_155), .Y(n_186) );
INVx1_ASAP7_75t_L g212 ( .A(n_31), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_32), .B(n_148), .Y(n_526) );
INVx2_ASAP7_75t_L g117 ( .A(n_33), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_34), .B(n_157), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_35), .B(n_148), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g121 ( .A1(n_36), .A2(n_119), .B(n_122), .C(n_125), .Y(n_121) );
INVx1_ASAP7_75t_L g210 ( .A(n_39), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_40), .B(n_155), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_41), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_42), .B(n_157), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_43), .A2(n_86), .B1(n_133), .B2(n_513), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_44), .B(n_157), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_45), .B(n_157), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_46), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_47), .B(n_480), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_48), .B(n_114), .Y(n_158) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_50), .A2(n_59), .B1(n_157), .B2(n_188), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_51), .A2(n_122), .B1(n_188), .B2(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_52), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_53), .B(n_157), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_54), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_55), .B(n_157), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_56), .A2(n_200), .B(n_201), .C(n_203), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_57), .Y(n_250) );
INVx1_ASAP7_75t_L g198 ( .A(n_58), .Y(n_198) );
INVx1_ASAP7_75t_L g120 ( .A(n_60), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_61), .B(n_157), .Y(n_505) );
INVx1_ASAP7_75t_L g139 ( .A(n_62), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_63), .Y(n_452) );
AO32x2_ASAP7_75t_L g546 ( .A1(n_64), .A2(n_144), .A3(n_147), .B1(n_482), .B2(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g478 ( .A(n_65), .Y(n_478) );
INVx1_ASAP7_75t_L g521 ( .A(n_66), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_SL g220 ( .A1(n_67), .A2(n_130), .B(n_203), .C(n_221), .Y(n_220) );
INVxp67_ASAP7_75t_L g222 ( .A(n_68), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_69), .B(n_188), .Y(n_522) );
INVx1_ASAP7_75t_L g455 ( .A(n_70), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_71), .Y(n_215) );
INVx1_ASAP7_75t_L g243 ( .A(n_72), .Y(n_243) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_73), .A2(n_103), .B1(n_447), .B2(n_456), .C1(n_753), .C2(n_758), .Y(n_102) );
OAI321xp33_ASAP7_75t_L g103 ( .A1(n_73), .A2(n_104), .A3(n_434), .B1(n_441), .B2(n_442), .C(n_444), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_73), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_74), .A2(n_88), .B1(n_432), .B2(n_433), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_74), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_76), .A2(n_119), .B(n_122), .C(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_77), .B(n_513), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_78), .A2(n_743), .B1(n_744), .B2(n_747), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_78), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_79), .B(n_188), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_80), .B(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_82), .B(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_83), .B(n_188), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_84), .A2(n_119), .B(n_122), .C(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g436 ( .A(n_85), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g461 ( .A(n_85), .B(n_438), .Y(n_461) );
INVx2_ASAP7_75t_L g465 ( .A(n_85), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_87), .A2(n_101), .B1(n_188), .B2(n_189), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_88), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_89), .B(n_148), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_90), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_91), .A2(n_119), .B(n_122), .C(n_151), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_92), .Y(n_160) );
INVx1_ASAP7_75t_L g219 ( .A(n_93), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g167 ( .A(n_94), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_95), .B(n_127), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_96), .B(n_188), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_97), .B(n_144), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_98), .A2(n_114), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_99), .B(n_455), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_100), .A2(n_458), .B1(n_741), .B2(n_742), .C1(n_748), .C2(n_751), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_104), .B(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_106), .B1(n_430), .B2(n_431), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_105), .A2(n_461), .B1(n_462), .B2(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_106), .A2(n_459), .B1(n_462), .B2(n_466), .Y(n_458) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_399), .Y(n_106) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_292), .C(n_365), .Y(n_107) );
OAI211xp5_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_177), .B(n_224), .C(n_276), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_145), .Y(n_110) );
AND2x2_ASAP7_75t_L g240 ( .A(n_111), .B(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g259 ( .A(n_111), .Y(n_259) );
INVx2_ASAP7_75t_L g274 ( .A(n_111), .Y(n_274) );
INVx1_ASAP7_75t_L g304 ( .A(n_111), .Y(n_304) );
AND2x2_ASAP7_75t_L g354 ( .A(n_111), .B(n_275), .Y(n_354) );
AOI32xp33_ASAP7_75t_L g381 ( .A1(n_111), .A2(n_309), .A3(n_382), .B1(n_384), .B2(n_385), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_111), .B(n_230), .Y(n_387) );
AND2x2_ASAP7_75t_L g414 ( .A(n_111), .B(n_257), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_111), .B(n_423), .Y(n_422) );
OR2x6_ASAP7_75t_L g111 ( .A(n_112), .B(n_141), .Y(n_111) );
AOI21xp5_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_121), .B(n_134), .Y(n_112) );
BUFx2_ASAP7_75t_L g165 ( .A(n_114), .Y(n_165) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_119), .Y(n_114) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_115), .B(n_119), .Y(n_182) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_118), .Y(n_115) );
INVx1_ASAP7_75t_L g480 ( .A(n_116), .Y(n_480) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g123 ( .A(n_117), .Y(n_123) );
INVx1_ASAP7_75t_L g189 ( .A(n_117), .Y(n_189) );
INVx1_ASAP7_75t_L g124 ( .A(n_118), .Y(n_124) );
INVx3_ASAP7_75t_L g128 ( .A(n_118), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_118), .Y(n_130) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_118), .Y(n_171) );
INVx4_ASAP7_75t_SL g175 ( .A(n_119), .Y(n_175) );
BUFx3_ASAP7_75t_L g482 ( .A(n_119), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_119), .A2(n_489), .B(n_492), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_119), .A2(n_499), .B(n_503), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_119), .A2(n_520), .B(n_523), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_119), .A2(n_529), .B(n_533), .Y(n_528) );
INVx5_ASAP7_75t_L g168 ( .A(n_122), .Y(n_168) );
AND2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
BUFx3_ASAP7_75t_L g133 ( .A(n_123), .Y(n_133) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
INVx1_ASAP7_75t_L g513 ( .A(n_123), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B(n_131), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_127), .A2(n_185), .B(n_186), .C(n_187), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_127), .A2(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_127), .A2(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g495 ( .A(n_127), .Y(n_495) );
O2A1O1Ixp5_ASAP7_75t_SL g520 ( .A1(n_127), .A2(n_203), .B(n_521), .C(n_522), .Y(n_520) );
INVx5_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_128), .B(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_128), .B(n_222), .Y(n_221) );
OAI22xp5_ASAP7_75t_SL g547 ( .A1(n_128), .A2(n_155), .B1(n_548), .B2(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g532 ( .A(n_130), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_131), .A2(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
INVx1_ASAP7_75t_L g248 ( .A(n_134), .Y(n_248) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_134), .A2(n_473), .B(n_483), .Y(n_472) );
OA21x2_ASAP7_75t_L g497 ( .A1(n_134), .A2(n_498), .B(n_506), .Y(n_497) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_135), .A2(n_180), .B(n_190), .Y(n_179) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_135), .A2(n_207), .B(n_214), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_135), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_137), .B(n_138), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
NOR2xp33_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
INVx3_ASAP7_75t_L g195 ( .A(n_143), .Y(n_195) );
AO21x1_ASAP7_75t_L g558 ( .A1(n_143), .A2(n_559), .B(n_562), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_143), .B(n_482), .C(n_559), .Y(n_583) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_144), .A2(n_217), .B(n_223), .Y(n_216) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_144), .A2(n_488), .B(n_496), .Y(n_487) );
AND2x2_ASAP7_75t_L g303 ( .A(n_145), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g325 ( .A(n_145), .Y(n_325) );
AND2x2_ASAP7_75t_L g410 ( .A(n_145), .B(n_240), .Y(n_410) );
AND2x2_ASAP7_75t_L g413 ( .A(n_145), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_162), .Y(n_145) );
INVx2_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_146), .B(n_257), .Y(n_263) );
AND2x2_ASAP7_75t_L g273 ( .A(n_146), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g309 ( .A(n_146), .Y(n_309) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_159), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_148), .A2(n_164), .B(n_176), .Y(n_163) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_148), .A2(n_519), .B(n_526), .Y(n_518) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_148), .A2(n_528), .B(n_536), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_158), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_156), .Y(n_151) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_155), .A2(n_495), .B1(n_512), .B2(n_514), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_155), .A2(n_495), .B1(n_560), .B2(n_561), .Y(n_559) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_161), .B(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_161), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g251 ( .A(n_162), .B(n_232), .Y(n_251) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g233 ( .A(n_163), .Y(n_233) );
AND2x2_ASAP7_75t_L g275 ( .A(n_163), .B(n_257), .Y(n_275) );
AND2x2_ASAP7_75t_L g344 ( .A(n_163), .B(n_241), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_169), .C(n_175), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_168), .A2(n_175), .B(n_198), .C(n_199), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_168), .A2(n_175), .B(n_219), .C(n_220), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_170), .B(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g502 ( .A(n_170), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_170), .A2(n_524), .B(n_525), .Y(n_523) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g209 ( .A1(n_171), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_209) );
INVx2_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g207 ( .A1(n_175), .A2(n_182), .B1(n_208), .B2(n_213), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_192), .Y(n_177) );
OR2x2_ASAP7_75t_L g238 ( .A(n_178), .B(n_206), .Y(n_238) );
INVx1_ASAP7_75t_L g317 ( .A(n_178), .Y(n_317) );
AND2x2_ASAP7_75t_L g331 ( .A(n_178), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_178), .B(n_205), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_178), .B(n_329), .Y(n_383) );
AND2x2_ASAP7_75t_L g391 ( .A(n_178), .B(n_392), .Y(n_391) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g228 ( .A(n_179), .Y(n_228) );
AND2x2_ASAP7_75t_L g298 ( .A(n_179), .B(n_206), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_182), .A2(n_243), .B(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_187), .A2(n_500), .B(n_501), .C(n_502), .Y(n_499) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_192), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g425 ( .A(n_192), .Y(n_425) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_205), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_193), .B(n_269), .Y(n_291) );
OR2x2_ASAP7_75t_L g320 ( .A(n_193), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g352 ( .A(n_193), .B(n_332), .Y(n_352) );
INVx1_ASAP7_75t_SL g372 ( .A(n_193), .Y(n_372) );
AND2x2_ASAP7_75t_L g376 ( .A(n_193), .B(n_237), .Y(n_376) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_SL g229 ( .A(n_194), .B(n_205), .Y(n_229) );
AND2x2_ASAP7_75t_L g236 ( .A(n_194), .B(n_216), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_194), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g279 ( .A(n_194), .B(n_261), .Y(n_279) );
INVx1_ASAP7_75t_SL g286 ( .A(n_194), .Y(n_286) );
BUFx2_ASAP7_75t_L g297 ( .A(n_194), .Y(n_297) );
AND2x2_ASAP7_75t_L g313 ( .A(n_194), .B(n_228), .Y(n_313) );
AND2x2_ASAP7_75t_L g328 ( .A(n_194), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g392 ( .A(n_194), .B(n_206), .Y(n_392) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_204), .Y(n_194) );
O2A1O1Ixp5_ASAP7_75t_L g477 ( .A1(n_200), .A2(n_478), .B(n_479), .C(n_481), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_200), .A2(n_534), .B(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_205), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g316 ( .A(n_205), .B(n_317), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_205), .A2(n_334), .B1(n_337), .B2(n_340), .C(n_345), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_205), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_216), .Y(n_205) );
INVx3_ASAP7_75t_L g261 ( .A(n_206), .Y(n_261) );
BUFx2_ASAP7_75t_L g271 ( .A(n_216), .Y(n_271) );
AND2x2_ASAP7_75t_L g285 ( .A(n_216), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g302 ( .A(n_216), .Y(n_302) );
OR2x2_ASAP7_75t_L g321 ( .A(n_216), .B(n_261), .Y(n_321) );
INVx3_ASAP7_75t_L g329 ( .A(n_216), .Y(n_329) );
AND2x2_ASAP7_75t_L g332 ( .A(n_216), .B(n_261), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_230), .B1(n_234), .B2(n_239), .C(n_252), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_227), .B(n_301), .Y(n_426) );
OR2x2_ASAP7_75t_L g429 ( .A(n_227), .B(n_260), .Y(n_429) );
INVx1_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
OAI221xp5_ASAP7_75t_SL g252 ( .A1(n_228), .A2(n_253), .B1(n_260), .B2(n_262), .C(n_265), .Y(n_252) );
AND2x2_ASAP7_75t_L g269 ( .A(n_228), .B(n_261), .Y(n_269) );
AND2x2_ASAP7_75t_L g277 ( .A(n_228), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_228), .B(n_285), .Y(n_284) );
NAND2x1_ASAP7_75t_L g327 ( .A(n_228), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g379 ( .A(n_228), .B(n_321), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_230), .A2(n_339), .B1(n_368), .B2(n_370), .Y(n_367) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AOI322xp5_ASAP7_75t_L g276 ( .A1(n_231), .A2(n_240), .A3(n_277), .B1(n_280), .B2(n_283), .C1(n_287), .C2(n_290), .Y(n_276) );
OR2x2_ASAP7_75t_L g288 ( .A(n_231), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_232), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g267 ( .A(n_232), .B(n_241), .Y(n_267) );
INVx1_ASAP7_75t_L g282 ( .A(n_232), .Y(n_282) );
AND2x2_ASAP7_75t_L g348 ( .A(n_232), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g258 ( .A(n_233), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g349 ( .A(n_233), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_233), .B(n_257), .Y(n_423) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_237), .B(n_372), .Y(n_371) );
INVx3_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g323 ( .A(n_238), .B(n_270), .Y(n_323) );
OR2x2_ASAP7_75t_L g420 ( .A(n_238), .B(n_271), .Y(n_420) );
INVx1_ASAP7_75t_L g401 ( .A(n_239), .Y(n_401) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_251), .Y(n_239) );
INVx4_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_240), .B(n_308), .Y(n_314) );
INVx2_ASAP7_75t_L g257 ( .A(n_241), .Y(n_257) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_248), .B(n_249), .Y(n_241) );
INVx1_ASAP7_75t_L g339 ( .A(n_251), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_251), .B(n_311), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g326 ( .A1(n_253), .A2(n_327), .B(n_330), .Y(n_326) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g311 ( .A(n_257), .Y(n_311) );
INVx1_ASAP7_75t_L g338 ( .A(n_257), .Y(n_338) );
INVx1_ASAP7_75t_L g264 ( .A(n_258), .Y(n_264) );
AND2x2_ASAP7_75t_L g266 ( .A(n_258), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g362 ( .A(n_259), .B(n_348), .Y(n_362) );
AND2x2_ASAP7_75t_L g384 ( .A(n_259), .B(n_344), .Y(n_384) );
BUFx2_ASAP7_75t_L g336 ( .A(n_261), .Y(n_336) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AOI32xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_268), .A3(n_269), .B1(n_270), .B2(n_272), .Y(n_265) );
INVx1_ASAP7_75t_L g346 ( .A(n_266), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_266), .A2(n_394), .B1(n_395), .B2(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_269), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_269), .B(n_328), .Y(n_369) );
AND2x2_ASAP7_75t_L g416 ( .A(n_269), .B(n_301), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_270), .B(n_317), .Y(n_364) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g417 ( .A(n_272), .Y(n_417) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_L g342 ( .A(n_273), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_275), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g389 ( .A(n_275), .B(n_309), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_275), .B(n_304), .Y(n_396) );
INVx1_ASAP7_75t_SL g378 ( .A(n_277), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_278), .B(n_329), .Y(n_356) );
NOR4xp25_ASAP7_75t_L g402 ( .A(n_278), .B(n_301), .C(n_403), .D(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_279), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVxp67_ASAP7_75t_L g359 ( .A(n_282), .Y(n_359) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_285), .A2(n_376), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g301 ( .A(n_286), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g350 ( .A(n_289), .Y(n_350) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND4xp25_ASAP7_75t_SL g292 ( .A(n_293), .B(n_318), .C(n_333), .D(n_353), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_299), .B(n_303), .C(n_305), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g385 ( .A(n_298), .B(n_328), .Y(n_385) );
AND2x2_ASAP7_75t_L g394 ( .A(n_298), .B(n_372), .Y(n_394) );
INVx3_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_301), .B(n_336), .Y(n_398) );
AND2x2_ASAP7_75t_L g310 ( .A(n_304), .B(n_311), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_312), .B1(n_314), .B2(n_315), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
AND2x2_ASAP7_75t_L g408 ( .A(n_308), .B(n_354), .Y(n_408) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_310), .B(n_359), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_311), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B(n_324), .C(n_326), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_319), .A2(n_354), .B1(n_355), .B2(n_357), .C(n_360), .Y(n_353) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_327), .A2(n_412), .B1(n_415), .B2(n_417), .C(n_418), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_328), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_336), .B(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g366 ( .A(n_338), .Y(n_366) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_341), .A2(n_361), .B1(n_363), .B2(n_364), .Y(n_360) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI21xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B(n_351), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_350), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_361), .A2(n_387), .B1(n_425), .B2(n_426), .C(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g406 ( .A(n_363), .Y(n_406) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_373), .C(n_393), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI211xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B(n_377), .C(n_386), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_380), .C(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g405 ( .A(n_383), .Y(n_405) );
OAI21xp5_ASAP7_75t_SL g427 ( .A1(n_384), .A2(n_410), .B(n_428), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI21xp5_ASAP7_75t_SL g419 ( .A1(n_396), .A2(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_411), .C(n_424), .Y(n_399) );
OAI211xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_407), .C(n_409), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
CKINVDCx14_ASAP7_75t_R g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g443 ( .A(n_436), .Y(n_443) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_436), .Y(n_446) );
INVx1_ASAP7_75t_SL g757 ( .A(n_436), .Y(n_757) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_437), .B(n_465), .Y(n_750) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g464 ( .A(n_438), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
OA21x2_ASAP7_75t_L g759 ( .A1(n_443), .A2(n_452), .B(n_453), .Y(n_759) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_448), .Y(n_447) );
CKINVDCx6p67_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NOR2xp33_ASAP7_75t_SL g755 ( .A(n_452), .B(n_454), .Y(n_755) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g752 ( .A(n_466), .Y(n_752) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR3x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_669), .C(n_718), .Y(n_467) );
NAND5xp2_ASAP7_75t_L g468 ( .A(n_469), .B(n_584), .C(n_612), .D(n_642), .E(n_656), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_507), .B1(n_537), .B2(n_542), .C(n_551), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_484), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_471), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g564 ( .A(n_472), .Y(n_564) );
AND2x2_ASAP7_75t_L g572 ( .A(n_472), .B(n_487), .Y(n_572) );
AND2x2_ASAP7_75t_L g595 ( .A(n_472), .B(n_486), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_472), .B(n_497), .Y(n_610) );
OR2x2_ASAP7_75t_L g619 ( .A(n_472), .B(n_558), .Y(n_619) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_472), .Y(n_622) );
AND2x2_ASAP7_75t_L g730 ( .A(n_472), .B(n_558), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_477), .B(n_482), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_479), .A2(n_495), .B(n_504), .C(n_505), .Y(n_503) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_484), .B(n_622), .Y(n_678) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
OAI311xp33_ASAP7_75t_L g620 ( .A1(n_485), .A2(n_621), .A3(n_622), .B1(n_623), .C1(n_638), .Y(n_620) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_497), .Y(n_485) );
AND2x2_ASAP7_75t_L g581 ( .A(n_486), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g588 ( .A(n_486), .Y(n_588) );
AND2x2_ASAP7_75t_L g709 ( .A(n_486), .B(n_541), .Y(n_709) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_487), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g565 ( .A(n_487), .B(n_497), .Y(n_565) );
AND2x2_ASAP7_75t_L g617 ( .A(n_487), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g631 ( .A(n_487), .B(n_564), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B(n_495), .Y(n_492) );
INVx2_ASAP7_75t_L g541 ( .A(n_497), .Y(n_541) );
AND2x2_ASAP7_75t_L g580 ( .A(n_497), .B(n_564), .Y(n_580) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_515), .Y(n_507) );
OR2x2_ASAP7_75t_L g675 ( .A(n_508), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_508), .B(n_681), .Y(n_692) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_509), .B(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g550 ( .A(n_510), .Y(n_550) );
AND2x2_ASAP7_75t_L g616 ( .A(n_510), .B(n_546), .Y(n_616) );
AND2x2_ASAP7_75t_L g627 ( .A(n_510), .B(n_527), .Y(n_627) );
AND2x2_ASAP7_75t_L g636 ( .A(n_510), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_515), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_515), .B(n_577), .Y(n_621) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g608 ( .A(n_516), .B(n_567), .Y(n_608) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_527), .Y(n_516) );
INVx2_ASAP7_75t_L g544 ( .A(n_517), .Y(n_544) );
AND2x2_ASAP7_75t_L g635 ( .A(n_517), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g554 ( .A(n_518), .Y(n_554) );
OR2x2_ASAP7_75t_L g652 ( .A(n_518), .B(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_518), .Y(n_715) );
AND2x2_ASAP7_75t_L g555 ( .A(n_527), .B(n_550), .Y(n_555) );
INVx1_ASAP7_75t_L g575 ( .A(n_527), .Y(n_575) );
AND2x2_ASAP7_75t_L g596 ( .A(n_527), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g637 ( .A(n_527), .Y(n_637) );
INVx1_ASAP7_75t_L g653 ( .A(n_527), .Y(n_653) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_527), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
INVxp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_539), .B(n_641), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_539), .A2(n_626), .B1(n_675), .B2(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
OAI211xp5_ASAP7_75t_SL g718 ( .A1(n_540), .A2(n_719), .B(n_721), .C(n_739), .Y(n_718) );
INVx2_ASAP7_75t_L g571 ( .A(n_541), .Y(n_571) );
AND2x2_ASAP7_75t_L g629 ( .A(n_541), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g640 ( .A(n_541), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_542), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
AND2x2_ASAP7_75t_L g613 ( .A(n_543), .B(n_577), .Y(n_613) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g645 ( .A(n_544), .B(n_636), .Y(n_645) );
AND2x2_ASAP7_75t_L g664 ( .A(n_544), .B(n_578), .Y(n_664) );
AND2x4_ASAP7_75t_L g600 ( .A(n_545), .B(n_574), .Y(n_600) );
AND2x2_ASAP7_75t_L g738 ( .A(n_545), .B(n_714), .Y(n_738) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_550), .Y(n_545) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_546), .Y(n_567) );
INVx1_ASAP7_75t_L g578 ( .A(n_546), .Y(n_578) );
INVx1_ASAP7_75t_L g677 ( .A(n_546), .Y(n_677) );
OR2x2_ASAP7_75t_L g568 ( .A(n_550), .B(n_554), .Y(n_568) );
AND2x2_ASAP7_75t_L g577 ( .A(n_550), .B(n_578), .Y(n_577) );
NOR2xp67_ASAP7_75t_L g597 ( .A(n_550), .B(n_598), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_556), .B1(n_566), .B2(n_569), .C(n_573), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_553), .A2(n_574), .B(n_576), .C(n_579), .Y(n_573) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g598 ( .A(n_554), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_554), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_SL g681 ( .A(n_554), .B(n_575), .Y(n_681) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_554), .Y(n_688) );
AND2x2_ASAP7_75t_L g606 ( .A(n_555), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g643 ( .A(n_555), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_565), .Y(n_556) );
INVx2_ASAP7_75t_L g634 ( .A(n_557), .Y(n_634) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_557), .A2(n_567), .B1(n_684), .B2(n_686), .C1(n_687), .C2(n_689), .Y(n_683) );
AND2x2_ASAP7_75t_L g740 ( .A(n_557), .B(n_709), .Y(n_740) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_564), .Y(n_557) );
INVx1_ASAP7_75t_L g630 ( .A(n_558), .Y(n_630) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g582 ( .A(n_563), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g668 ( .A(n_565), .B(n_602), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g679 ( .A1(n_566), .A2(n_680), .B(n_682), .Y(n_679) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx2_ASAP7_75t_L g607 ( .A(n_567), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_567), .B(n_574), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_567), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx3_ASAP7_75t_L g633 ( .A(n_571), .Y(n_633) );
OR2x2_ASAP7_75t_L g685 ( .A(n_571), .B(n_607), .Y(n_685) );
AND2x2_ASAP7_75t_L g601 ( .A(n_572), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g639 ( .A(n_572), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_572), .B(n_633), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_572), .B(n_629), .Y(n_655) );
AND2x2_ASAP7_75t_L g659 ( .A(n_572), .B(n_641), .Y(n_659) );
INVxp67_ASAP7_75t_L g591 ( .A(n_574), .Y(n_591) );
BUFx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_576), .A2(n_649), .B1(n_654), .B2(n_655), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_576), .B(n_681), .Y(n_711) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g697 ( .A(n_577), .B(n_688), .Y(n_697) );
AND2x2_ASAP7_75t_L g726 ( .A(n_577), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g731 ( .A(n_577), .B(n_681), .Y(n_731) );
INVx1_ASAP7_75t_L g644 ( .A(n_578), .Y(n_644) );
BUFx2_ASAP7_75t_L g650 ( .A(n_578), .Y(n_650) );
INVx1_ASAP7_75t_L g735 ( .A(n_579), .Y(n_735) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_580), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g611 ( .A(n_581), .Y(n_611) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_582), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g594 ( .A(n_582), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g603 ( .A(n_582), .Y(n_603) );
INVx3_ASAP7_75t_L g641 ( .A(n_582), .Y(n_641) );
OR2x2_ASAP7_75t_L g707 ( .A(n_582), .B(n_708), .Y(n_707) );
AOI211xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_589), .B(n_592), .C(n_604), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_585), .A2(n_722), .B1(n_729), .B2(n_731), .C(n_732), .Y(n_721) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_593), .B(n_599), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_595), .B(n_633), .Y(n_647) );
AND2x2_ASAP7_75t_L g689 ( .A(n_595), .B(n_629), .Y(n_689) );
INVx1_ASAP7_75t_SL g702 ( .A(n_596), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_596), .B(n_650), .Y(n_705) );
INVx1_ASAP7_75t_L g723 ( .A(n_597), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_601), .A2(n_691), .B1(n_693), .B2(n_697), .C(n_698), .Y(n_690) );
AND2x2_ASAP7_75t_L g717 ( .A(n_602), .B(n_709), .Y(n_717) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g701 ( .A(n_603), .Y(n_701) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_608), .B(n_609), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g672 ( .A(n_607), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g658 ( .A(n_608), .Y(n_658) );
INVx1_ASAP7_75t_L g686 ( .A(n_609), .Y(n_686) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B(n_617), .C(n_620), .Y(n_612) );
OAI31xp33_ASAP7_75t_L g739 ( .A1(n_613), .A2(n_651), .A3(n_738), .B(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g713 ( .A(n_616), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g734 ( .A(n_616), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_618), .B(n_633), .Y(n_661) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g736 ( .A(n_619), .B(n_633), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_628), .B1(n_632), .B2(n_635), .Y(n_623) );
NAND2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_627), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g663 ( .A(n_627), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g666 ( .A(n_627), .B(n_650), .Y(n_666) );
AND2x2_ASAP7_75t_L g720 ( .A(n_627), .B(n_715), .Y(n_720) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g695 ( .A(n_631), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
OAI32xp33_ASAP7_75t_L g698 ( .A1(n_633), .A2(n_667), .A3(n_699), .B1(n_701), .B2(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g673 ( .A(n_636), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_636), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g696 ( .A(n_640), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B(n_646), .C(n_648), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_644), .B(n_681), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_645), .A2(n_657), .B1(n_658), .B2(n_659), .C(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g657 ( .A(n_655), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_665), .B2(n_667), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND4xp25_ASAP7_75t_SL g722 ( .A(n_665), .B(n_723), .C(n_724), .D(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
NAND4xp25_ASAP7_75t_SL g669 ( .A(n_670), .B(n_683), .C(n_690), .D(n_703), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B(n_678), .C(n_679), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g700 ( .A(n_676), .Y(n_700) );
INVx2_ASAP7_75t_L g724 ( .A(n_681), .Y(n_724) );
OR2x2_ASAP7_75t_L g733 ( .A(n_688), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_706), .B(n_710), .Y(n_703) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g729 ( .A(n_709), .B(n_730), .Y(n_729) );
AOI21xp33_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_712), .B(n_716), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
CKINVDCx16_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
NAND2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
endmodule