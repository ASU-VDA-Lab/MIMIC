module fake_jpeg_7978_n_170 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx10_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_20),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_11),
.B1(n_19),
.B2(n_18),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_28),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_26),
.B1(n_24),
.B2(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_42),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_29),
.B(n_21),
.C(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_46),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_26),
.B1(n_24),
.B2(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_27),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_19),
.B(n_16),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.C(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_25),
.Y(n_51)
);

OR2x2_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_20),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_12),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_56),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_62),
.B1(n_65),
.B2(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_64),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_26),
.B1(n_24),
.B2(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_65),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_30),
.C(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_23),
.B1(n_36),
.B2(n_22),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_23),
.B1(n_36),
.B2(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_16),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_46),
.B1(n_52),
.B2(n_48),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_78),
.B(n_61),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_32),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_94),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_56),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_89),
.C(n_58),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_60),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_53),
.B(n_55),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_94),
.B(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_79),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_75),
.B1(n_73),
.B2(n_76),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_107),
.B1(n_111),
.B2(n_21),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_103),
.Y(n_117)
);

XNOR2x1_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_106),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_87),
.C(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_57),
.B(n_58),
.Y(n_107)
);

NAND2x1p5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_25),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_13),
.B1(n_33),
.B2(n_17),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_18),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_7),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_114),
.C(n_118),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_13),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_103),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_33),
.C(n_27),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_13),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_126),
.C(n_109),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_100),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_123),
.A2(n_125),
.B(n_108),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_129),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_135),
.B(n_5),
.Y(n_146)
);

AOI31xp67_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_109),
.A3(n_104),
.B(n_115),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_132),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_134),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_96),
.C(n_13),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_7),
.B(n_10),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_6),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_33),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_117),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_132),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_144),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_124),
.Y(n_144)
);

NAND4xp25_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_121),
.C(n_118),
.D(n_7),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_4),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_141),
.B(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_139),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_0),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_6),
.C(n_9),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_8),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_146),
.B1(n_141),
.B2(n_9),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_150),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_156),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_158),
.B(n_159),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_143),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_153),
.B(n_151),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_162),
.B(n_164),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_15),
.B(n_17),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_3),
.B(n_9),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_17),
.C(n_15),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_166),
.A2(n_167),
.B(n_3),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_3),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_169),
.Y(n_170)
);

OAI321xp33_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_15),
.C(n_154),
.Y(n_169)
);


endmodule