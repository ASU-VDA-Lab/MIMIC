module fake_jpeg_1537_n_227 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_227);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_0),
.B(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_0),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_78),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_54),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_58),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_55),
.B1(n_57),
.B2(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_99),
.B1(n_79),
.B2(n_61),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_97),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_61),
.B1(n_57),
.B2(n_70),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_58),
.B1(n_83),
.B2(n_75),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_74),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_70),
.B1(n_60),
.B2(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_113),
.B1(n_73),
.B2(n_71),
.Y(n_129)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_58),
.B1(n_52),
.B2(n_74),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_118),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_52),
.B1(n_65),
.B2(n_68),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_115),
.A2(n_95),
.B1(n_98),
.B2(n_91),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_120),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_65),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_1),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_95),
.B1(n_91),
.B2(n_75),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_69),
.B(n_77),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_130),
.B(n_133),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_67),
.B(n_64),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_53),
.B1(n_66),
.B2(n_56),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_138),
.B1(n_107),
.B2(n_106),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_116),
.B(n_104),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_38),
.C(n_50),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_110),
.C(n_111),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_63),
.B1(n_2),
.B2(n_3),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_141),
.B(n_26),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_147),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_111),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_35),
.C(n_46),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_157),
.C(n_31),
.Y(n_172)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_63),
.B1(n_4),
.B2(n_5),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_45),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_162),
.B1(n_13),
.B2(n_14),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_1),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_159),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_44),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_43),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_4),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_5),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_40),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_39),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_131),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_164),
.B(n_165),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_6),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_6),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_7),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_34),
.B(n_32),
.Y(n_171)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_167),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_176),
.B(n_187),
.Y(n_193)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_23),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_177),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_14),
.B(n_16),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_158),
.B1(n_149),
.B2(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_183),
.Y(n_202)
);

AO22x1_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_17),
.C(n_18),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_157),
.C(n_150),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_177),
.B1(n_169),
.B2(n_188),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_20),
.B(n_22),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_162),
.B(n_161),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_191),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_180),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_195),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_23),
.B(n_182),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_198),
.C(n_200),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_189),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_176),
.C(n_185),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_196),
.B(n_179),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_209),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_173),
.B1(n_179),
.B2(n_186),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_190),
.B1(n_198),
.B2(n_194),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_202),
.B(n_178),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_172),
.C(n_183),
.Y(n_210)
);

AOI31xp33_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_199),
.A3(n_194),
.B(n_193),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_216),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_207),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_214),
.B(n_193),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_203),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_206),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_217),
.B(n_216),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_218),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_222),
.B(n_218),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_213),
.Y(n_227)
);


endmodule