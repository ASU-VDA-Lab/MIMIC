module fake_jpeg_1653_n_476 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_48),
.Y(n_122)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_49),
.Y(n_127)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_14),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_63),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_14),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_13),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_71),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_35),
.B(n_13),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_17),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_12),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_80),
.Y(n_126)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_12),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_12),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_36),
.B(n_11),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_11),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_36),
.B(n_11),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_98),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_31),
.B(n_9),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_34),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_106),
.A2(n_108),
.B1(n_121),
.B2(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_56),
.B1(n_42),
.B2(n_48),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_157),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_42),
.B1(n_38),
.B2(n_23),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_39),
.B1(n_33),
.B2(n_26),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_150),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_62),
.A2(n_39),
.B1(n_33),
.B2(n_26),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_134),
.A2(n_135),
.B1(n_100),
.B2(n_81),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_25),
.B1(n_23),
.B2(n_29),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_49),
.A2(n_25),
.B1(n_29),
.B2(n_44),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_144),
.A2(n_148),
.B1(n_100),
.B2(n_72),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_52),
.A2(n_44),
.B1(n_15),
.B2(n_40),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_60),
.A2(n_34),
.B1(n_15),
.B2(n_22),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_91),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_95),
.A2(n_22),
.B1(n_40),
.B2(n_9),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_151),
.A2(n_90),
.B1(n_93),
.B2(n_99),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_68),
.A2(n_40),
.B1(n_1),
.B2(n_2),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_71),
.B(n_64),
.C(n_86),
.Y(n_176)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_70),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_163),
.B(n_166),
.Y(n_222)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_152),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_103),
.B(n_57),
.C(n_87),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_167),
.B(n_189),
.C(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_82),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_168),
.B(n_170),
.Y(n_244)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_119),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_9),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_174),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_209),
.B1(n_153),
.B2(n_145),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_180),
.Y(n_216)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_190),
.Y(n_230)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_59),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_116),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_115),
.B1(n_114),
.B2(n_148),
.Y(n_217)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_112),
.B(n_55),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_92),
.B(n_85),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_192),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_194),
.Y(n_239)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_224)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_96),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_208),
.Y(n_238)
);

BUFx2_ASAP7_75t_SL g204 ( 
.A(n_137),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_109),
.B(n_78),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_153),
.Y(n_236)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_134),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_217),
.A2(n_220),
.B1(n_252),
.B2(n_118),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_172),
.A2(n_135),
.B1(n_144),
.B2(n_158),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_172),
.A2(n_186),
.B1(n_167),
.B2(n_206),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_248),
.B1(n_250),
.B2(n_200),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_165),
.B(n_104),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_251),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_181),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_158),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_246),
.C(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_117),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_235),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_117),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_183),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_189),
.B(n_127),
.C(n_162),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_179),
.B(n_127),
.C(n_140),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_176),
.B1(n_212),
.B2(n_189),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_184),
.A2(n_147),
.B1(n_159),
.B2(n_143),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_184),
.B(n_118),
.C(n_157),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_192),
.A2(n_159),
.B1(n_147),
.B2(n_143),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_230),
.A2(n_200),
.B(n_185),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_253),
.A2(n_257),
.B(n_268),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_273),
.B1(n_274),
.B2(n_279),
.Y(n_288)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_256),
.B(n_258),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_203),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_263),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_198),
.B(n_188),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_260),
.A2(n_247),
.B(n_239),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_199),
.B1(n_197),
.B2(n_195),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_261),
.A2(n_218),
.B1(n_215),
.B2(n_227),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_262),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_216),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_270),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_220),
.A2(n_202),
.B1(n_193),
.B2(n_194),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_175),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_164),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_271),
.B(n_281),
.Y(n_309)
);

INVxp67_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_280),
.B(n_224),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_221),
.A2(n_110),
.B1(n_125),
.B2(n_173),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_276),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_216),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_229),
.A2(n_125),
.B1(n_162),
.B2(n_154),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_243),
.A2(n_169),
.B1(n_113),
.B2(n_154),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_1),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_226),
.B(n_1),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_282),
.B(n_251),
.Y(n_303)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_291),
.A2(n_307),
.B1(n_274),
.B2(n_279),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_254),
.A2(n_232),
.B1(n_226),
.B2(n_222),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_292),
.A2(n_298),
.B1(n_300),
.B2(n_266),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_225),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_308),
.C(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_274),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_297),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_260),
.A2(n_222),
.B1(n_236),
.B2(n_233),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_214),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_270),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_260),
.A2(n_252),
.B1(n_250),
.B2(n_214),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_264),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_304),
.Y(n_327)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_237),
.C(n_239),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_315),
.Y(n_343)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_294),
.B(n_272),
.CI(n_264),
.CON(n_311),
.SN(n_311)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_318),
.C(n_293),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_263),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_314),
.B(n_329),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_269),
.Y(n_316)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_283),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_321),
.Y(n_336)
);

OA21x2_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_272),
.B(n_267),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_332),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_283),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_287),
.B(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_286),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_282),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_334),
.C(n_303),
.Y(n_335)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_288),
.A2(n_274),
.B1(n_273),
.B2(n_261),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_330),
.A2(n_331),
.B1(n_304),
.B2(n_297),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_288),
.A2(n_257),
.B1(n_276),
.B2(n_281),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_296),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_277),
.Y(n_333)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_333),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_282),
.C(n_281),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_350),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_338),
.A2(n_342),
.B1(n_351),
.B2(n_359),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_316),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_345),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_341),
.B(n_311),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_331),
.A2(n_321),
.B1(n_317),
.B2(n_329),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_325),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_347),
.A2(n_291),
.B1(n_280),
.B2(n_312),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_325),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_349),
.B(n_328),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_292),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_327),
.A2(n_306),
.B1(n_285),
.B2(n_301),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_303),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_358),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_301),
.Y(n_353)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_353),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_289),
.C(n_285),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_357),
.C(n_284),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_289),
.C(n_284),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_309),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_327),
.A2(n_297),
.B1(n_300),
.B2(n_298),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_296),
.Y(n_360)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_360),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_320),
.B(n_326),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_379),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_342),
.A2(n_330),
.B1(n_268),
.B2(n_319),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_363),
.B1(n_372),
.B2(n_380),
.Y(n_385)
);

AOI21xp33_ASAP7_75t_L g364 ( 
.A1(n_346),
.A2(n_253),
.B(n_286),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_364),
.B(n_368),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_355),
.Y(n_367)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_367),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_360),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_335),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_325),
.Y(n_371)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_336),
.Y(n_372)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_338),
.A2(n_319),
.B1(n_326),
.B2(n_309),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_373),
.A2(n_380),
.B1(n_381),
.B2(n_359),
.Y(n_386)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_384),
.Y(n_390)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_348),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

NOR3xp33_ASAP7_75t_SL g393 ( 
.A(n_382),
.B(n_344),
.C(n_337),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_311),
.C(n_253),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_383),
.B(n_350),
.C(n_352),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_256),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_385),
.A2(n_395),
.B1(n_381),
.B2(n_361),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_386),
.A2(n_401),
.B1(n_402),
.B2(n_365),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_365),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_392),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_375),
.Y(n_392)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_363),
.A2(n_347),
.B1(n_357),
.B2(n_356),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_341),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_371),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_358),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_379),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_373),
.A2(n_272),
.B1(n_354),
.B2(n_259),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_367),
.A2(n_271),
.B1(n_354),
.B2(n_312),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_369),
.Y(n_404)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_375),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_408),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_383),
.C(n_377),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_362),
.C(n_366),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_412),
.C(n_415),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_370),
.Y(n_411)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_411),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_366),
.C(n_378),
.Y(n_412)
);

BUFx24_ASAP7_75t_SL g413 ( 
.A(n_394),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_417),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_414),
.A2(n_397),
.B1(n_401),
.B2(n_391),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_376),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_416),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_242),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_305),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_420),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_385),
.A2(n_382),
.B1(n_305),
.B2(n_218),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_422),
.A2(n_228),
.B1(n_223),
.B2(n_234),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_409),
.A2(n_397),
.B(n_399),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_424),
.A2(n_426),
.B(n_407),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_406),
.A2(n_396),
.B(n_390),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_412),
.A2(n_398),
.B(n_390),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_431),
.B(n_223),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_435),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_408),
.A2(n_396),
.B(n_242),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_433),
.B(n_238),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_241),
.C(n_234),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_436),
.A2(n_440),
.B(n_445),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_410),
.C(n_241),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_438),
.Y(n_452)
);

AOI211xp5_ASAP7_75t_L g440 ( 
.A1(n_434),
.A2(n_245),
.B(n_219),
.C(n_215),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_425),
.B(n_245),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_441),
.B(n_442),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_421),
.B(n_227),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_444),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_228),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_228),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_446),
.B(n_433),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_426),
.A2(n_223),
.B(n_249),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_447),
.A2(n_422),
.B1(n_431),
.B2(n_435),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_423),
.Y(n_448)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_448),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_454),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_436),
.A2(n_432),
.B(n_428),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_451),
.A2(n_457),
.B(n_8),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_428),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_455),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_444),
.B(n_432),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_448),
.A2(n_438),
.B1(n_443),
.B2(n_249),
.Y(n_458)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

NOR3xp33_ASAP7_75t_SL g460 ( 
.A(n_451),
.B(n_8),
.C(n_4),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_460),
.A2(n_463),
.B(n_464),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_456),
.A2(n_452),
.B(n_450),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_453),
.C(n_4),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_3),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_461),
.A2(n_3),
.B(n_4),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_467),
.A2(n_3),
.B(n_5),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_462),
.C(n_4),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_469),
.A2(n_5),
.B(n_6),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g473 ( 
.A1(n_470),
.A2(n_471),
.B(n_466),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_472),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_473),
.C(n_6),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_475),
.A2(n_5),
.B(n_7),
.Y(n_476)
);


endmodule