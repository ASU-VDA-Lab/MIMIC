module fake_jpeg_29567_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_47),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_16),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_74),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_79),
.Y(n_93)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_64),
.B1(n_62),
.B2(n_68),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_64),
.B1(n_62),
.B2(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_89),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_68),
.B1(n_53),
.B2(n_60),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_90),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_69),
.B1(n_53),
.B2(n_58),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_108),
.B1(n_109),
.B2(n_96),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_55),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_9),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_110),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_58),
.B(n_54),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_109),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_67),
.B1(n_25),
.B2(n_27),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_2),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_9),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_115),
.B1(n_122),
.B2(n_99),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

OAI211xp5_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_28),
.B(n_48),
.C(n_46),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_130),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_20),
.C(n_42),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_119),
.C(n_131),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_19),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_8),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_129),
.Y(n_133)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_30),
.C(n_40),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_29),
.A3(n_39),
.B1(n_35),
.B2(n_14),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_32),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_10),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_23),
.B(n_31),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_139),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_34),
.B(n_50),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_123),
.B(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_126),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_128),
.B1(n_147),
.B2(n_138),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_142),
.B(n_134),
.C(n_147),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_141),
.B(n_133),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_155),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_149),
.C(n_156),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_153),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_148),
.B1(n_151),
.B2(n_146),
.C(n_143),
.Y(n_162)
);


endmodule