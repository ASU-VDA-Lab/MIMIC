module fake_netlist_1_2966_n_26 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
NAND2xp5_ASAP7_75t_L g12 ( .A(n_9), .B(n_11), .Y(n_12) );
BUFx3_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
NAND2xp33_ASAP7_75t_SL g14 ( .A(n_1), .B(n_2), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_7), .B(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_13), .B(n_0), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_15), .B(n_4), .Y(n_18) );
AO31x2_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_12), .A3(n_14), .B(n_16), .Y(n_19) );
AOI211xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_18), .B(n_15), .C(n_10), .Y(n_20) );
NAND2x1_ASAP7_75t_L g21 ( .A(n_20), .B(n_5), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_6), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_23), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVxp67_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
endmodule