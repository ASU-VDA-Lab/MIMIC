module fake_aes_8118_n_803 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_191, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_803);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_803;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_384;
wire n_227;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_560;
wire n_517;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_771;
wire n_696;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_198;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g195 ( .A(n_36), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_14), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_101), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_98), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_22), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_49), .Y(n_202) );
INVx1_ASAP7_75t_SL g203 ( .A(n_106), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_4), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_71), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_126), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_103), .Y(n_207) );
CKINVDCx14_ASAP7_75t_R g208 ( .A(n_176), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_69), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_72), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_14), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_191), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_76), .Y(n_214) );
INVx1_ASAP7_75t_SL g215 ( .A(n_65), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_83), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_122), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_172), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_47), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_50), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_76), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_173), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_141), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_121), .Y(n_224) );
BUFx8_ASAP7_75t_SL g225 ( .A(n_145), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_108), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_150), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_42), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_87), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_30), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_84), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_11), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_139), .Y(n_234) );
NOR2xp67_ASAP7_75t_L g235 ( .A(n_93), .B(n_48), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_183), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_180), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_104), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_127), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_136), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_188), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_115), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_102), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_8), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_129), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_181), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_128), .Y(n_247) );
NOR2xp67_ASAP7_75t_L g248 ( .A(n_80), .B(n_157), .Y(n_248) );
BUFx2_ASAP7_75t_SL g249 ( .A(n_21), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_165), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_94), .Y(n_251) );
BUFx5_ASAP7_75t_L g252 ( .A(n_193), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_175), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_186), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_112), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_162), .Y(n_256) );
BUFx2_ASAP7_75t_SL g257 ( .A(n_134), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_4), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_159), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_138), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_137), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_177), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_133), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_163), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_51), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_187), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_192), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g268 ( .A(n_64), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_37), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_58), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_20), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_68), .Y(n_272) );
INVxp67_ASAP7_75t_L g273 ( .A(n_100), .Y(n_273) );
BUFx5_ASAP7_75t_L g274 ( .A(n_143), .Y(n_274) );
INVxp67_ASAP7_75t_L g275 ( .A(n_117), .Y(n_275) );
NOR2xp67_ASAP7_75t_L g276 ( .A(n_13), .B(n_144), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_54), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_55), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_99), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_65), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_97), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_130), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_182), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_110), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_53), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_124), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_82), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_161), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_184), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_190), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_116), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_18), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_17), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_174), .B(n_153), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_140), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_88), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_146), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_148), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_89), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_149), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_61), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_132), .Y(n_302) );
INVxp67_ASAP7_75t_L g303 ( .A(n_135), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_34), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_154), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_1), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_62), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_210), .B(n_0), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_252), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_207), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_233), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_263), .B(n_0), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_282), .B(n_1), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_277), .Y(n_314) );
OAI22x1_ASAP7_75t_L g315 ( .A1(n_285), .A2(n_5), .B1(n_2), .B2(n_3), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_210), .Y(n_316) );
AND2x6_ASAP7_75t_L g317 ( .A(n_253), .B(n_90), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_252), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_301), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_252), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_207), .Y(n_321) );
NAND2xp33_ASAP7_75t_L g322 ( .A(n_252), .B(n_194), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_252), .Y(n_323) );
NOR2x1_ASAP7_75t_L g324 ( .A(n_301), .B(n_3), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_196), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_243), .B(n_5), .Y(n_326) );
OAI22xp5_ASAP7_75t_SL g327 ( .A1(n_214), .A2(n_9), .B1(n_6), .B2(n_7), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_252), .Y(n_328) );
OA21x2_ASAP7_75t_L g329 ( .A1(n_217), .A2(n_92), .B(n_91), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_209), .B(n_6), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_306), .B(n_7), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_253), .B(n_10), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_268), .A2(n_15), .B1(n_12), .B2(n_13), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_198), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_217), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_199), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_252), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_274), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_260), .B(n_12), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_256), .B(n_15), .Y(n_340) );
INVx5_ASAP7_75t_L g341 ( .A(n_207), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_225), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_206), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_307), .B(n_16), .Y(n_344) );
OR2x6_ASAP7_75t_L g345 ( .A(n_342), .B(n_249), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_309), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_325), .B(n_228), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_317), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_332), .Y(n_349) );
INVx5_ASAP7_75t_L g350 ( .A(n_317), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
NAND3xp33_ASAP7_75t_L g353 ( .A(n_313), .B(n_231), .C(n_211), .Y(n_353) );
NOR2x1p5_ASAP7_75t_L g354 ( .A(n_342), .B(n_223), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_310), .Y(n_355) );
AND2x6_ASAP7_75t_L g356 ( .A(n_332), .B(n_260), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
AND2x6_ASAP7_75t_L g358 ( .A(n_332), .B(n_261), .Y(n_358) );
NAND2xp33_ASAP7_75t_SL g359 ( .A(n_330), .B(n_312), .Y(n_359) );
NAND3xp33_ASAP7_75t_L g360 ( .A(n_313), .B(n_265), .C(n_258), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_332), .Y(n_361) );
NOR2x1p5_ASAP7_75t_L g362 ( .A(n_326), .B(n_223), .Y(n_362) );
NOR2x1p5_ASAP7_75t_L g363 ( .A(n_326), .B(n_255), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_310), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_308), .A2(n_197), .B1(n_201), .B2(n_195), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_339), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_340), .B(n_331), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_310), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_333), .A2(n_230), .B1(n_238), .B2(n_222), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_339), .Y(n_370) );
BUFx4f_ASAP7_75t_L g371 ( .A(n_317), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_339), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_318), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_318), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_317), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_334), .B(n_336), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_339), .B(n_319), .Y(n_377) );
OR2x6_ASAP7_75t_L g378 ( .A(n_327), .B(n_257), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_371), .B(n_320), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_367), .Y(n_380) );
INVx4_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_347), .B(n_343), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_367), .B(n_340), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_377), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_359), .A2(n_333), .B1(n_230), .B2(n_238), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_376), .B(n_319), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_362), .B(n_316), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_363), .B(n_284), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_378), .A2(n_219), .B1(n_232), .B2(n_214), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_371), .B(n_320), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_377), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_353), .B(n_344), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_377), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_365), .B(n_322), .C(n_269), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_356), .B(n_286), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_356), .B(n_288), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_345), .B(n_324), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_352), .Y(n_400) );
AND2x6_ASAP7_75t_L g401 ( .A(n_366), .B(n_324), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_352), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_358), .B(n_289), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_358), .B(n_208), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_371), .B(n_320), .Y(n_405) );
AND2x6_ASAP7_75t_SL g406 ( .A(n_378), .B(n_202), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_345), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_350), .B(n_323), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_360), .A2(n_270), .B1(n_215), .B2(n_205), .C(n_216), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_349), .A2(n_329), .B(n_328), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_357), .B(n_311), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_357), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_366), .A2(n_335), .B1(n_317), .B2(n_328), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_350), .B(n_323), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_366), .B(n_335), .Y(n_415) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_378), .A2(n_219), .B1(n_244), .B2(n_232), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_372), .B(n_314), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_372), .B(n_314), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_349), .B(n_224), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_350), .B(n_328), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_361), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_361), .B(n_227), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_370), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_370), .A2(n_317), .B1(n_338), .B2(n_337), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_346), .B(n_234), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_351), .B(n_237), .Y(n_426) );
NOR2xp33_ASAP7_75t_SL g427 ( .A(n_345), .B(n_244), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_354), .A2(n_315), .B1(n_204), .B2(n_221), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_348), .B(n_220), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_351), .B(n_200), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_375), .B(n_229), .Y(n_431) );
NOR2xp67_ASAP7_75t_L g432 ( .A(n_369), .B(n_337), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_410), .A2(n_391), .B(n_379), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_380), .B(n_383), .Y(n_434) );
OAI21xp33_ASAP7_75t_SL g435 ( .A1(n_382), .A2(n_378), .B(n_374), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_382), .B(n_373), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_393), .A2(n_373), .B(n_338), .C(n_337), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_394), .Y(n_438) );
O2A1O1Ixp5_ASAP7_75t_SL g439 ( .A1(n_388), .A2(n_213), .B(n_218), .C(n_212), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_427), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_385), .Y(n_441) );
OAI21x1_ASAP7_75t_L g442 ( .A1(n_424), .A2(n_329), .B(n_355), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_405), .A2(n_329), .B(n_226), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_385), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_392), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_432), .A2(n_271), .B1(n_278), .B2(n_272), .Y(n_446) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_384), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_407), .B(n_280), .Y(n_448) );
BUFx12f_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
CKINVDCx11_ASAP7_75t_R g450 ( .A(n_399), .Y(n_450) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_428), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_393), .B(n_287), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_409), .A2(n_293), .B(n_304), .C(n_292), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_402), .A2(n_317), .B(n_240), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_430), .B(n_264), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_386), .A2(n_235), .B1(n_276), .B2(n_248), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_430), .B(n_273), .Y(n_457) );
AOI33xp33_ASAP7_75t_L g458 ( .A1(n_390), .A2(n_281), .A3(n_247), .B1(n_239), .B2(n_241), .B3(n_305), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_387), .A2(n_246), .B1(n_251), .B2(n_242), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_400), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_401), .B(n_275), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_401), .B(n_303), .Y(n_462) );
INVx4_ASAP7_75t_L g463 ( .A(n_395), .Y(n_463) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_397), .A2(n_236), .B(n_203), .Y(n_464) );
INVx8_ASAP7_75t_L g465 ( .A(n_401), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_395), .Y(n_466) );
AOI21x1_ASAP7_75t_L g467 ( .A1(n_404), .A2(n_364), .B(n_355), .Y(n_467) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_396), .B(n_283), .C(n_267), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_411), .A2(n_299), .B(n_254), .C(n_262), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_398), .B(n_266), .Y(n_470) );
NOR2xp67_ASAP7_75t_L g471 ( .A(n_389), .B(n_17), .Y(n_471) );
BUFx4f_ASAP7_75t_L g472 ( .A(n_429), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_390), .Y(n_474) );
BUFx12f_ASAP7_75t_L g475 ( .A(n_429), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_403), .B(n_296), .Y(n_476) );
CKINVDCx6p67_ASAP7_75t_R g477 ( .A(n_431), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_418), .A2(n_262), .B(n_279), .C(n_250), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_415), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_412), .A2(n_290), .B(n_291), .C(n_279), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_416), .B(n_302), .C(n_294), .Y(n_481) );
AO32x1_ASAP7_75t_L g482 ( .A1(n_421), .A2(n_298), .A3(n_290), .B1(n_291), .B2(n_295), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_423), .A2(n_297), .B1(n_298), .B2(n_295), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_419), .Y(n_484) );
NOR3xp33_ASAP7_75t_L g485 ( .A(n_416), .B(n_368), .C(n_364), .Y(n_485) );
INVx8_ASAP7_75t_L g486 ( .A(n_413), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_422), .B(n_18), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_426), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_425), .B(n_19), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_408), .A2(n_245), .B(n_259), .C(n_207), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_414), .A2(n_259), .B1(n_300), .B2(n_245), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_420), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_410), .A2(n_341), .B(n_300), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_380), .B(n_274), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_381), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_380), .B(n_274), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g497 ( .A(n_390), .B(n_23), .C(n_24), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_385), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_385), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_410), .A2(n_341), .B(n_321), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_380), .B(n_274), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_380), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_380), .B(n_25), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_380), .Y(n_504) );
BUFx12f_ASAP7_75t_L g505 ( .A(n_406), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_380), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_385), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_410), .A2(n_96), .B(n_95), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_380), .B(n_26), .Y(n_509) );
AO31x2_ASAP7_75t_L g510 ( .A1(n_443), .A2(n_29), .A3(n_27), .B(n_28), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_495), .Y(n_511) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_433), .A2(n_31), .A3(n_29), .B(n_30), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_484), .B(n_32), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_504), .B(n_32), .Y(n_514) );
OAI22x1_ASAP7_75t_L g515 ( .A1(n_474), .A2(n_35), .B1(n_33), .B2(n_34), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_506), .B(n_33), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_444), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_445), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_473), .B(n_35), .Y(n_519) );
OAI22x1_ASAP7_75t_L g520 ( .A1(n_440), .A2(n_38), .B1(n_36), .B2(n_37), .Y(n_520) );
BUFx3_ASAP7_75t_L g521 ( .A(n_475), .Y(n_521) );
AND2x2_ASAP7_75t_SL g522 ( .A(n_472), .B(n_39), .Y(n_522) );
AO31x2_ASAP7_75t_L g523 ( .A1(n_480), .A2(n_40), .A3(n_41), .B(n_43), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_446), .B(n_43), .Y(n_525) );
AO31x2_ASAP7_75t_L g526 ( .A1(n_508), .A2(n_44), .A3(n_45), .B(n_46), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_488), .B(n_46), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_477), .Y(n_528) );
OAI21x1_ASAP7_75t_L g529 ( .A1(n_467), .A2(n_107), .B(n_105), .Y(n_529) );
OR2x6_ASAP7_75t_L g530 ( .A(n_505), .B(n_48), .Y(n_530) );
OAI21x1_ASAP7_75t_L g531 ( .A1(n_500), .A2(n_111), .B(n_109), .Y(n_531) );
BUFx12f_ASAP7_75t_L g532 ( .A(n_450), .Y(n_532) );
INVx4_ASAP7_75t_L g533 ( .A(n_472), .Y(n_533) );
INVx3_ASAP7_75t_SL g534 ( .A(n_509), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_495), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_503), .Y(n_536) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_436), .A2(n_114), .B(n_113), .Y(n_537) );
BUFx8_ASAP7_75t_L g538 ( .A(n_448), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_479), .A2(n_119), .B(n_118), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_458), .B(n_52), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_454), .A2(n_123), .B(n_120), .Y(n_541) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_499), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_454), .A2(n_142), .B(n_189), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_452), .B(n_56), .Y(n_545) );
INVx3_ASAP7_75t_SL g546 ( .A(n_448), .Y(n_546) );
CKINVDCx11_ASAP7_75t_R g547 ( .A(n_465), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_451), .B(n_57), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_494), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_496), .Y(n_550) );
AO31x2_ASAP7_75t_L g551 ( .A1(n_491), .A2(n_58), .A3(n_59), .B(n_60), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_497), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_507), .Y(n_553) );
AOI221x1_ASAP7_75t_L g554 ( .A1(n_491), .A2(n_63), .B1(n_66), .B2(n_67), .C(n_69), .Y(n_554) );
AOI221x1_ASAP7_75t_L g555 ( .A1(n_459), .A2(n_70), .B1(n_71), .B2(n_72), .C(n_73), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_447), .Y(n_556) );
OR2x6_ASAP7_75t_L g557 ( .A(n_465), .B(n_74), .Y(n_557) );
NOR2x1_ASAP7_75t_SL g558 ( .A(n_495), .B(n_75), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_455), .B(n_457), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_501), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_470), .A2(n_152), .B(n_179), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_438), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_466), .Y(n_563) );
AO31x2_ASAP7_75t_L g564 ( .A1(n_490), .A2(n_77), .A3(n_78), .B(n_79), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_489), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_464), .A2(n_478), .B(n_462), .C(n_461), .Y(n_566) );
AND2x4_ASAP7_75t_L g567 ( .A(n_498), .B(n_81), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_441), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_476), .A2(n_155), .B(n_178), .Y(n_569) );
AO32x2_ASAP7_75t_L g570 ( .A1(n_482), .A2(n_463), .A3(n_468), .B1(n_486), .B2(n_483), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_471), .A2(n_85), .B(n_86), .C(n_125), .Y(n_571) );
AO31x2_ASAP7_75t_L g572 ( .A1(n_482), .A2(n_131), .A3(n_147), .B(n_156), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_492), .A2(n_164), .B1(n_166), .B2(n_167), .Y(n_573) );
AOI221xp5_ASAP7_75t_SL g574 ( .A1(n_460), .A2(n_168), .B1(n_169), .B2(n_170), .C(n_171), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_493), .A2(n_410), .B(n_433), .Y(n_575) );
O2A1O1Ixp33_ASAP7_75t_L g576 ( .A1(n_456), .A2(n_453), .B(n_435), .C(n_469), .Y(n_576) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_466), .Y(n_577) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_493), .A2(n_442), .B(n_467), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_502), .B(n_380), .Y(n_579) );
BUFx3_ASAP7_75t_L g580 ( .A(n_475), .Y(n_580) );
AO31x2_ASAP7_75t_L g581 ( .A1(n_443), .A2(n_493), .A3(n_433), .B(n_469), .Y(n_581) );
BUFx4f_ASAP7_75t_SL g582 ( .A(n_449), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_439), .A2(n_433), .B(n_437), .Y(n_583) );
OA21x2_ASAP7_75t_L g584 ( .A1(n_443), .A2(n_410), .B(n_442), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_493), .A2(n_410), .B(n_433), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_485), .A2(n_380), .B1(n_481), .B2(n_474), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_434), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g588 ( .A1(n_435), .A2(n_382), .B(n_393), .C(n_487), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_444), .Y(n_589) );
BUFx3_ASAP7_75t_L g590 ( .A(n_521), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_522), .B(n_534), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_559), .B(n_588), .Y(n_592) );
INVx4_ASAP7_75t_L g593 ( .A(n_547), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_587), .B(n_565), .Y(n_594) );
AOI21xp5_ASAP7_75t_SL g595 ( .A1(n_527), .A2(n_557), .B(n_513), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_546), .B(n_513), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_584), .A2(n_566), .B(n_576), .Y(n_597) );
OA21x2_ASAP7_75t_L g598 ( .A1(n_574), .A2(n_529), .B(n_531), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_514), .Y(n_599) );
AO31x2_ASAP7_75t_L g600 ( .A1(n_554), .A2(n_555), .A3(n_544), .B(n_541), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_545), .A2(n_540), .B(n_519), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_586), .B(n_536), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_556), .B(n_548), .Y(n_603) );
OR2x6_ASAP7_75t_L g604 ( .A(n_557), .B(n_533), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_568), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_580), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_550), .B(n_560), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_516), .B(n_528), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_518), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_567), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_543), .Y(n_612) );
OA21x2_ASAP7_75t_L g613 ( .A1(n_571), .A2(n_569), .B(n_561), .Y(n_613) );
BUFx12f_ASAP7_75t_L g614 ( .A(n_530), .Y(n_614) );
CKINVDCx11_ASAP7_75t_R g615 ( .A(n_530), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_553), .B(n_589), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_549), .B(n_525), .Y(n_617) );
OA21x2_ASAP7_75t_L g618 ( .A1(n_570), .A2(n_573), .B(n_552), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_581), .B(n_535), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_510), .Y(n_620) );
OR2x6_ASAP7_75t_L g621 ( .A(n_515), .B(n_520), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_581), .B(n_563), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_523), .Y(n_623) );
OAI21x1_ASAP7_75t_L g624 ( .A1(n_581), .A2(n_577), .B(n_524), .Y(n_624) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_524), .A2(n_542), .B(n_563), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_542), .B(n_523), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_572), .A2(n_526), .B(n_512), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_551), .B(n_564), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_551), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_579), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_579), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_533), .B(n_380), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_579), .Y(n_633) );
AOI21xp5_ASAP7_75t_SL g634 ( .A1(n_527), .A2(n_557), .B(n_513), .Y(n_634) );
INVx6_ASAP7_75t_L g635 ( .A(n_538), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_562), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_533), .B(n_472), .Y(n_637) );
NAND2x1_ASAP7_75t_L g638 ( .A(n_511), .B(n_535), .Y(n_638) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_533), .B(n_472), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_562), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_579), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_562), .Y(n_642) );
AO31x2_ASAP7_75t_L g643 ( .A1(n_575), .A2(n_585), .A3(n_588), .B(n_443), .Y(n_643) );
AO31x2_ASAP7_75t_L g644 ( .A1(n_575), .A2(n_585), .A3(n_588), .B(n_443), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_579), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_533), .B(n_380), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_522), .B(n_380), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_559), .B(n_473), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_522), .B(n_380), .Y(n_649) );
OA21x2_ASAP7_75t_L g650 ( .A1(n_578), .A2(n_574), .B(n_583), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g651 ( .A(n_582), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_559), .B(n_473), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_562), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_579), .Y(n_654) );
OAI21x1_ASAP7_75t_SL g655 ( .A1(n_558), .A2(n_539), .B(n_537), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_579), .Y(n_656) );
OAI21x1_ASAP7_75t_SL g657 ( .A1(n_558), .A2(n_539), .B(n_537), .Y(n_657) );
BUFx8_ASAP7_75t_L g658 ( .A(n_532), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_559), .B(n_473), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_562), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_559), .B(n_473), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_559), .B(n_473), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_629), .Y(n_663) );
OR2x6_ASAP7_75t_L g664 ( .A(n_595), .B(n_634), .Y(n_664) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_611), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_592), .B(n_607), .Y(n_666) );
AO21x2_ASAP7_75t_L g667 ( .A1(n_627), .A2(n_628), .B(n_597), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_643), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_619), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_637), .Y(n_670) );
BUFx3_ASAP7_75t_L g671 ( .A(n_590), .Y(n_671) );
BUFx3_ASAP7_75t_L g672 ( .A(n_606), .Y(n_672) );
BUFx3_ASAP7_75t_L g673 ( .A(n_632), .Y(n_673) );
OR2x6_ASAP7_75t_L g674 ( .A(n_604), .B(n_621), .Y(n_674) );
INVx8_ASAP7_75t_L g675 ( .A(n_604), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_623), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_635), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_636), .B(n_640), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_630), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_631), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_642), .B(n_653), .Y(n_681) );
BUFx12f_ASAP7_75t_L g682 ( .A(n_658), .Y(n_682) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_616), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_648), .B(n_652), .Y(n_684) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_593), .B(n_614), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_644), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_620), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_644), .Y(n_688) );
OR2x6_ASAP7_75t_L g689 ( .A(n_604), .B(n_621), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_633), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_659), .B(n_661), .Y(n_691) );
BUFx12f_ASAP7_75t_L g692 ( .A(n_658), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_660), .B(n_602), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_602), .B(n_609), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_626), .Y(n_695) );
BUFx12f_ASAP7_75t_L g696 ( .A(n_651), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_637), .Y(n_697) );
INVx3_ASAP7_75t_L g698 ( .A(n_639), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_594), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_624), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_610), .B(n_612), .Y(n_701) );
AO21x2_ASAP7_75t_L g702 ( .A1(n_622), .A2(n_657), .B(n_655), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_605), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_662), .B(n_601), .Y(n_704) );
BUFx2_ASAP7_75t_L g705 ( .A(n_625), .Y(n_705) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_641), .Y(n_706) );
INVx2_ASAP7_75t_SL g707 ( .A(n_635), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_646), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_647), .A2(n_649), .B1(n_603), .B2(n_615), .Y(n_709) );
OR2x6_ASAP7_75t_L g710 ( .A(n_596), .B(n_599), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_663), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_683), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_675), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_676), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_684), .B(n_645), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_666), .B(n_650), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_669), .B(n_617), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_691), .B(n_656), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_695), .B(n_600), .Y(n_719) );
BUFx3_ASAP7_75t_L g720 ( .A(n_671), .Y(n_720) );
INVx2_ASAP7_75t_SL g721 ( .A(n_675), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_704), .B(n_618), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_672), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_691), .B(n_617), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_687), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_699), .B(n_654), .Y(n_726) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_664), .B(n_593), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_672), .B(n_591), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_705), .Y(n_729) );
INVx2_ASAP7_75t_SL g730 ( .A(n_675), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_702), .B(n_638), .Y(n_731) );
BUFx3_ASAP7_75t_L g732 ( .A(n_708), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_693), .B(n_608), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_678), .B(n_598), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_681), .B(n_613), .Y(n_735) );
BUFx3_ASAP7_75t_L g736 ( .A(n_673), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_694), .B(n_703), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_703), .B(n_701), .Y(n_738) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_679), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_738), .B(n_680), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_722), .B(n_668), .Y(n_741) );
AND2x2_ASAP7_75t_SL g742 ( .A(n_712), .B(n_729), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_738), .B(n_690), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_735), .B(n_702), .Y(n_744) );
CKINVDCx16_ASAP7_75t_R g745 ( .A(n_720), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_714), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_711), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_739), .B(n_686), .Y(n_748) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_727), .B(n_664), .Y(n_749) );
BUFx2_ASAP7_75t_L g750 ( .A(n_732), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_733), .B(n_688), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_716), .B(n_667), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_737), .B(n_706), .Y(n_753) );
INVx4_ASAP7_75t_L g754 ( .A(n_736), .Y(n_754) );
NOR2xp67_ASAP7_75t_L g755 ( .A(n_723), .B(n_682), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_732), .Y(n_756) );
AND2x4_ASAP7_75t_L g757 ( .A(n_719), .B(n_700), .Y(n_757) );
INVx4_ASAP7_75t_L g758 ( .A(n_736), .Y(n_758) );
NOR2xp33_ASAP7_75t_SL g759 ( .A(n_755), .B(n_682), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_746), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_747), .Y(n_761) );
NAND2x1_ASAP7_75t_L g762 ( .A(n_749), .B(n_727), .Y(n_762) );
OR2x2_ASAP7_75t_L g763 ( .A(n_753), .B(n_717), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_740), .B(n_674), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_743), .B(n_725), .Y(n_765) );
NAND2x1_ASAP7_75t_L g766 ( .A(n_749), .B(n_674), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_744), .B(n_731), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_751), .B(n_724), .Y(n_768) );
NAND2x1p5_ASAP7_75t_L g769 ( .A(n_754), .B(n_685), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_745), .B(n_689), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_752), .B(n_734), .Y(n_771) );
INVx2_ASAP7_75t_SL g772 ( .A(n_769), .Y(n_772) );
INVx2_ASAP7_75t_SL g773 ( .A(n_769), .Y(n_773) );
OAI22xp33_ASAP7_75t_L g774 ( .A1(n_766), .A2(n_689), .B1(n_754), .B2(n_758), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_765), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_760), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_761), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_760), .Y(n_778) );
OAI32xp33_ASAP7_75t_L g779 ( .A1(n_770), .A2(n_754), .A3(n_758), .B1(n_728), .B2(n_756), .Y(n_779) );
INVxp67_ASAP7_75t_L g780 ( .A(n_759), .Y(n_780) );
OAI221xp5_ASAP7_75t_SL g781 ( .A1(n_764), .A2(n_709), .B1(n_710), .B2(n_718), .C(n_715), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_771), .B(n_741), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_771), .B(n_741), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_777), .Y(n_784) );
AOI31xp33_ASAP7_75t_L g785 ( .A1(n_780), .A2(n_713), .A3(n_721), .B(n_730), .Y(n_785) );
O2A1O1Ixp33_ASAP7_75t_L g786 ( .A1(n_779), .A2(n_707), .B(n_677), .C(n_671), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_781), .A2(n_762), .B1(n_742), .B2(n_768), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_772), .A2(n_742), .B1(n_763), .B2(n_767), .Y(n_788) );
AOI222xp33_ASAP7_75t_L g789 ( .A1(n_787), .A2(n_775), .B1(n_774), .B2(n_779), .C1(n_782), .C2(n_783), .Y(n_789) );
AOI211xp5_ASAP7_75t_L g790 ( .A1(n_788), .A2(n_772), .B(n_773), .C(n_707), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_786), .B(n_692), .Y(n_791) );
AOI22x1_ASAP7_75t_L g792 ( .A1(n_785), .A2(n_692), .B1(n_696), .B2(n_750), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_784), .Y(n_793) );
OAI211xp5_ASAP7_75t_L g794 ( .A1(n_791), .A2(n_792), .B(n_789), .C(n_790), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_794), .B(n_793), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_795), .B(n_748), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_796), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_797), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_798), .A2(n_726), .B1(n_665), .B2(n_710), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g800 ( .A1(n_799), .A2(n_670), .B(n_698), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_800), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_801), .B(n_697), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_802), .A2(n_757), .B1(n_776), .B2(n_778), .Y(n_803) );
endmodule