module fake_jpeg_1786_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_48),
.Y(n_51)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_57),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_34),
.B1(n_40),
.B2(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_31),
.B1(n_38),
.B2(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_37),
.Y(n_57)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_66),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_32),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_53),
.Y(n_70)
);

AO22x1_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_29),
.B1(n_14),
.B2(n_16),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_53),
.B1(n_35),
.B2(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_77),
.B(n_39),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_62),
.B(n_35),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_33),
.Y(n_79)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_52),
.B(n_58),
.C(n_59),
.D(n_4),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_33),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AOI221xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_104)
);

OA21x2_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_93),
.B(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_91),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_74),
.B(n_8),
.Y(n_94)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_90),
.B1(n_70),
.B2(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_6),
.Y(n_93)
);

AOI21x1_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_104),
.B(n_10),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_70),
.B1(n_79),
.B2(n_9),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_99),
.B1(n_27),
.B2(n_13),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_19),
.B(n_25),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_7),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_109),
.Y(n_112)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_97),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_100),
.C(n_107),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_99),
.B1(n_101),
.B2(n_110),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_110),
.B(n_112),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_94),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_103),
.C(n_20),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_17),
.Y(n_121)
);


endmodule