module fake_jpeg_4686_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_31),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_58),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_2),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_69),
.A2(n_50),
.B1(n_55),
.B2(n_44),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_51),
.B1(n_53),
.B2(n_52),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_47),
.B1(n_59),
.B2(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_87),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_45),
.B1(n_61),
.B2(n_5),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_80),
.B(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_84),
.B1(n_89),
.B2(n_75),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_93),
.B1(n_92),
.B2(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_15),
.C(n_16),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_20),
.C(n_21),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_24),
.B(n_26),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_28),
.B(n_29),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_33),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_39),
.Y(n_106)
);


endmodule