module real_jpeg_33121_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI211xp5_ASAP7_75t_L g8 ( 
.A1(n_0),
.A2(n_9),
.B(n_10),
.C(n_34),
.Y(n_8)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx2_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_21),
.Y(n_32)
);

AND2x4_ASAP7_75t_SL g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_5),
.A2(n_6),
.B1(n_15),
.B2(n_21),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_11),
.A2(n_24),
.B1(n_28),
.B2(n_33),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_17),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_15),
.B(n_16),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_18),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_23),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AND2x4_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_40),
.B1(n_43),
.B2(n_46),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);


endmodule