module fake_jpeg_2482_n_610 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_610);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_610;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_58),
.B(n_61),
.Y(n_119)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_59),
.Y(n_141)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_R g68 ( 
.A(n_21),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_108),
.Y(n_149)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_84),
.Y(n_143)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_28),
.B(n_17),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_40),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_88),
.B(n_90),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_91),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g169 ( 
.A(n_93),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_94),
.B(n_96),
.Y(n_179)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_28),
.B(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_99),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_39),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_30),
.B(n_17),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_30),
.B(n_14),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_34),
.B(n_15),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_31),
.Y(n_105)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g109 ( 
.A(n_20),
.Y(n_109)
);

BUFx16f_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_39),
.B1(n_27),
.B2(n_53),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_116),
.A2(n_130),
.B1(n_135),
.B2(n_137),
.Y(n_195)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_49),
.CON(n_118),
.SN(n_118)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_118),
.B(n_23),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_64),
.A2(n_34),
.B1(n_39),
.B2(n_49),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_132),
.B(n_82),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_70),
.A2(n_55),
.B1(n_50),
.B2(n_45),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_72),
.A2(n_36),
.B1(n_50),
.B2(n_45),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_59),
.B(n_55),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_174),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_149),
.Y(n_223)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_151),
.Y(n_185)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_158),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_73),
.A2(n_38),
.B1(n_44),
.B2(n_43),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_43),
.B1(n_24),
.B2(n_35),
.Y(n_189)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_76),
.B(n_38),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_68),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_183),
.Y(n_262)
);

OR2x2_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_79),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_186),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_179),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_187),
.B(n_200),
.C(n_205),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_189),
.A2(n_204),
.B1(n_206),
.B2(n_217),
.Y(n_277)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_120),
.B(n_24),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_191),
.B(n_193),
.Y(n_245)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_192),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_44),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g274 ( 
.A(n_194),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_137),
.A2(n_36),
.B1(n_22),
.B2(n_52),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_196),
.Y(n_294)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_35),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_199),
.B(n_228),
.Y(n_300)
);

CKINVDCx12_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_78),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_203),
.B(n_220),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_116),
.A2(n_41),
.B1(n_77),
.B2(n_92),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_115),
.A2(n_41),
.B1(n_74),
.B2(n_91),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_207),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_209),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_119),
.B(n_110),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_211),
.B(n_221),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_124),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_143),
.A2(n_119),
.B(n_125),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_225),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_153),
.A2(n_36),
.B1(n_52),
.B2(n_42),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_141),
.B(n_95),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_143),
.B(n_85),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_163),
.A2(n_60),
.B1(n_69),
.B2(n_63),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_222),
.A2(n_224),
.B1(n_230),
.B2(n_241),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_128),
.A2(n_23),
.B1(n_42),
.B2(n_52),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_148),
.B(n_65),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_123),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_15),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_117),
.B(n_15),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_231),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_173),
.A2(n_42),
.B1(n_23),
.B2(n_112),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_141),
.B(n_13),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_138),
.B(n_12),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_234),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_127),
.A2(n_67),
.B(n_93),
.C(n_107),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_121),
.B(n_113),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_150),
.B(n_89),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_136),
.Y(n_235)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_235),
.Y(n_279)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_144),
.Y(n_239)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_243),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_133),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_144),
.Y(n_242)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

INVx3_ASAP7_75t_SL g243 ( 
.A(n_134),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_124),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_244)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_165),
.B1(n_172),
.B2(n_177),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_184),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_250),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_183),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_252),
.B(n_255),
.C(n_11),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_129),
.C(n_126),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_258),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_195),
.A2(n_142),
.B1(n_177),
.B2(n_172),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_263),
.A2(n_276),
.B1(n_288),
.B2(n_299),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_207),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_284),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_205),
.A2(n_155),
.B(n_169),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_269),
.A2(n_285),
.B(n_299),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_185),
.B(n_131),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_271),
.B(n_273),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_166),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_220),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_189),
.A2(n_142),
.B1(n_146),
.B2(n_156),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_213),
.B(n_156),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_198),
.B(n_146),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_233),
.A2(n_155),
.B(n_3),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_183),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_184),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_289),
.B(n_256),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_182),
.B(n_5),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_292),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_186),
.B(n_6),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_237),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_209),
.B(n_6),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_291),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_203),
.A2(n_7),
.B(n_8),
.Y(n_299)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_304),
.Y(n_367)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_307),
.Y(n_393)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_248),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_309),
.B(n_313),
.Y(n_398)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_236),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_314),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_188),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_248),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_282),
.B(n_249),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_317),
.Y(n_362)
);

AND2x2_ASAP7_75t_SL g316 ( 
.A(n_262),
.B(n_203),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_350),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_265),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g318 ( 
.A(n_254),
.B(n_194),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_318),
.B(n_324),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_319),
.A2(n_274),
.B1(n_295),
.B2(n_272),
.Y(n_383)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_263),
.A2(n_244),
.B1(n_235),
.B2(n_227),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_321),
.A2(n_323),
.B1(n_328),
.B2(n_336),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_276),
.A2(n_226),
.B1(n_190),
.B2(n_239),
.Y(n_323)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_252),
.B(n_269),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_270),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_331),
.Y(n_373)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_253),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_332),
.Y(n_391)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_220),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_348),
.B(n_292),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_347),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_294),
.A2(n_242),
.B1(n_208),
.B2(n_197),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_277),
.A2(n_240),
.B1(n_237),
.B2(n_188),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_337),
.A2(n_342),
.B1(n_344),
.B2(n_349),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_294),
.A2(n_202),
.B1(n_243),
.B2(n_214),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_338),
.A2(n_345),
.B1(n_274),
.B2(n_287),
.Y(n_384)
);

O2A1O1Ixp33_ASAP7_75t_SL g339 ( 
.A1(n_285),
.A2(n_213),
.B(n_212),
.C(n_219),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_339),
.A2(n_272),
.B(n_287),
.Y(n_386)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_247),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_340),
.B(n_343),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_282),
.B(n_219),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_346),
.Y(n_374)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_246),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

INVx13_ASAP7_75t_L g344 ( 
.A(n_253),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_280),
.A2(n_212),
.B1(n_181),
.B2(n_215),
.Y(n_345)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_259),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_181),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_280),
.B(n_11),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_261),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_351),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_290),
.B(n_9),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_260),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_262),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_356),
.C(n_360),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_316),
.B(n_255),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_383),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_268),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_324),
.C(n_302),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_363),
.B(n_379),
.C(n_380),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_353),
.A2(n_258),
.B(n_278),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_366),
.A2(n_378),
.B(n_392),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_319),
.A2(n_275),
.B1(n_251),
.B2(n_300),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_369),
.A2(n_372),
.B1(n_382),
.B2(n_390),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_245),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_385),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_319),
.A2(n_275),
.B1(n_286),
.B2(n_288),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_329),
.A2(n_281),
.B(n_293),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_293),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_308),
.B(n_260),
.C(n_295),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_335),
.A2(n_275),
.B1(n_286),
.B2(n_259),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_384),
.A2(n_394),
.B1(n_339),
.B2(n_331),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_267),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_386),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g404 ( 
.A(n_387),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_318),
.A2(n_246),
.B1(n_267),
.B2(n_11),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_329),
.A2(n_9),
.B(n_10),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_336),
.A2(n_10),
.B1(n_338),
.B2(n_345),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_305),
.B(n_306),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_397),
.B(n_340),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_322),
.B(n_330),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_399),
.B(n_348),
.Y(n_414)
);

INVx11_ASAP7_75t_L g400 ( 
.A(n_364),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_400),
.A2(n_377),
.B1(n_384),
.B2(n_366),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_399),
.B(n_371),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_408),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_330),
.Y(n_405)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_405),
.B(n_420),
.C(n_421),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_368),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_398),
.Y(n_409)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_409),
.Y(n_456)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_410),
.Y(n_459)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

INVx13_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_413),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_419),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_361),
.B(n_322),
.Y(n_415)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_415),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_429),
.Y(n_443)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_418),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_361),
.B(n_348),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_325),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_375),
.B(n_343),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_424),
.Y(n_449)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_388),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_375),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_363),
.B(n_332),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_355),
.C(n_360),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_311),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_428),
.Y(n_452)
);

INVx13_ASAP7_75t_L g427 ( 
.A(n_367),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_427),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_320),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_369),
.B(n_326),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_430),
.B(n_431),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_359),
.B(n_304),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_433),
.A2(n_436),
.B1(n_372),
.B2(n_382),
.Y(n_464)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_437),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_381),
.A2(n_321),
.B1(n_312),
.B2(n_323),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_374),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_370),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_367),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_356),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_441),
.B(n_445),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_403),
.A2(n_365),
.B(n_386),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_444),
.A2(n_446),
.B(n_417),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_354),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_434),
.A2(n_417),
.B(n_378),
.Y(n_446)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_448),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_354),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_451),
.B(n_462),
.Y(n_497)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_457),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_405),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_460),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_357),
.Y(n_460)
);

OAI32xp33_ASAP7_75t_L g461 ( 
.A1(n_424),
.A2(n_391),
.A3(n_359),
.B1(n_396),
.B2(n_389),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_379),
.C(n_358),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_432),
.C(n_421),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_464),
.A2(n_465),
.B1(n_469),
.B2(n_410),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_406),
.A2(n_381),
.B1(n_392),
.B2(n_396),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_409),
.B(n_370),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_466),
.B(n_472),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_434),
.A2(n_383),
.B(n_389),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_468),
.A2(n_417),
.B(n_408),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_406),
.A2(n_393),
.B1(n_342),
.B2(n_349),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_422),
.Y(n_472)
);

XNOR2x2_ASAP7_75t_SL g473 ( 
.A(n_407),
.B(n_327),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_473),
.B(n_426),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_401),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_476),
.B(n_479),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_477),
.B(n_452),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_478),
.A2(n_450),
.B(n_447),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_453),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_480),
.A2(n_473),
.B(n_469),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_464),
.A2(n_430),
.B1(n_402),
.B2(n_407),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_481),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_440),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_483),
.B(n_494),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_465),
.A2(n_436),
.B1(n_415),
.B2(n_428),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_484),
.A2(n_452),
.B1(n_440),
.B2(n_447),
.Y(n_516)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_485),
.Y(n_508)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_456),
.Y(n_486)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_486),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_487),
.Y(n_532)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_442),
.Y(n_489)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_489),
.Y(n_521)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_492),
.Y(n_526)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_443),
.Y(n_493)
);

BUFx4f_ASAP7_75t_SL g515 ( 
.A(n_493),
.Y(n_515)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_449),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_437),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_496),
.Y(n_512)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_449),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_500),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_463),
.B(n_414),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_471),
.A2(n_404),
.B1(n_438),
.B2(n_419),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_501),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_462),
.B(n_435),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_505),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_441),
.B(n_412),
.C(n_429),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_504),
.B(n_445),
.C(n_459),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_451),
.B(n_423),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_506),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_507),
.B(n_488),
.Y(n_539)
);

NOR2x1_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_459),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_SL g549 ( 
.A(n_509),
.B(n_522),
.C(n_524),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_516),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_504),
.B(n_444),
.C(n_468),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_529),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_446),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_520),
.B(n_523),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_491),
.B(n_497),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_503),
.A2(n_474),
.B(n_470),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_525),
.A2(n_481),
.B(n_467),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_484),
.A2(n_470),
.B1(n_455),
.B2(n_439),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_527),
.A2(n_490),
.B1(n_418),
.B2(n_431),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_498),
.B(n_439),
.C(n_467),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_482),
.B(n_474),
.Y(n_531)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_531),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_507),
.B(n_502),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_533),
.B(n_538),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_511),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_534),
.B(n_537),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_528),
.B(n_497),
.C(n_505),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_536),
.B(n_539),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_500),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_480),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_515),
.B(n_499),
.Y(n_541)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_541),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_477),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_542),
.B(n_546),
.Y(n_563)
);

OA21x2_ASAP7_75t_SL g543 ( 
.A1(n_510),
.A2(n_475),
.B(n_499),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_543),
.B(n_515),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_514),
.B(n_501),
.Y(n_546)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_547),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_548),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_508),
.Y(n_550)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_550),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_515),
.B(n_346),
.Y(n_551)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_551),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_528),
.B(n_490),
.C(n_393),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_532),
.C(n_521),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_549),
.A2(n_509),
.B(n_530),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_559),
.B(n_524),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_550),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_562),
.B(n_568),
.Y(n_572)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_564),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_535),
.B(n_518),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_569),
.Y(n_581)
);

MAJx2_ASAP7_75t_L g567 ( 
.A(n_546),
.B(n_530),
.C(n_519),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_567),
.B(n_539),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_540),
.B(n_529),
.Y(n_568)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_548),
.Y(n_570)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_570),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_552),
.A2(n_513),
.B1(n_526),
.B2(n_506),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_571),
.B(n_527),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_573),
.B(n_575),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_555),
.B(n_544),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_566),
.B(n_533),
.C(n_536),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_576),
.B(n_579),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_577),
.A2(n_557),
.B(n_571),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_560),
.B(n_553),
.C(n_542),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_580),
.B(n_567),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_569),
.B(n_512),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_582),
.B(n_583),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_561),
.B(n_522),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_513),
.C(n_545),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_584),
.B(n_585),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_556),
.B(n_565),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_554),
.C(n_557),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_587),
.Y(n_598)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_588),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_574),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_593),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_581),
.B(n_559),
.C(n_563),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_SL g596 ( 
.A1(n_590),
.A2(n_572),
.B(n_578),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_596),
.B(n_589),
.Y(n_602)
);

AOI322xp5_ASAP7_75t_L g597 ( 
.A1(n_592),
.A2(n_558),
.A3(n_545),
.B1(n_506),
.B2(n_584),
.C1(n_517),
.C2(n_427),
.Y(n_597)
);

OAI321xp33_ASAP7_75t_L g601 ( 
.A1(n_597),
.A2(n_594),
.A3(n_592),
.B1(n_400),
.B2(n_413),
.C(n_427),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_558),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_599),
.A2(n_579),
.B(n_576),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_601),
.B(n_602),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_603),
.B(n_598),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_604),
.A2(n_600),
.B(n_605),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_606),
.A2(n_595),
.B1(n_563),
.B2(n_400),
.Y(n_607)
);

NOR4xp25_ASAP7_75t_L g608 ( 
.A(n_607),
.B(n_516),
.C(n_538),
.D(n_413),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_608),
.B(n_344),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_609),
.A2(n_310),
.B(n_307),
.Y(n_610)
);


endmodule