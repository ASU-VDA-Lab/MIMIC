module real_jpeg_12237_n_13 (n_46, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_45, n_6, n_44, n_7, n_3, n_10, n_9, n_13);

input n_46;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_45;
input n_6;
input n_44;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_17;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_31;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_14;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_1),
.C(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_2),
.A2(n_6),
.B(n_16),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_6),
.C(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_29),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_5),
.C(n_16),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_7),
.A2(n_16),
.B(n_44),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_16),
.C(n_46),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_9),
.A2(n_11),
.B(n_16),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_9),
.B(n_11),
.C(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_18),
.B(n_19),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_10),
.B(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_33),
.B(n_34),
.Y(n_32)
);

NOR3xp33_ASAP7_75t_L g35 ( 
.A(n_10),
.B(n_33),
.C(n_34),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_38),
.B(n_39),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_20),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_17),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B(n_42),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_37),
.B(n_40),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_36),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_35),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_31),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_45),
.Y(n_30)
);


endmodule