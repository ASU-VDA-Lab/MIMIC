module fake_jpeg_1394_n_197 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_47),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_74),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_60),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_52),
.B1(n_58),
.B2(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_57),
.B1(n_63),
.B2(n_58),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_53),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_64),
.B1(n_62),
.B2(n_59),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_76),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_59),
.B1(n_49),
.B2(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_49),
.B1(n_64),
.B2(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_96),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_89),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_88),
.B1(n_89),
.B2(n_77),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_103),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_107),
.B1(n_105),
.B2(n_104),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NAND2x1_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_62),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_61),
.B1(n_70),
.B2(n_76),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_75),
.B1(n_73),
.B2(n_53),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_117),
.B(n_29),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_118),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_54),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_13),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_68),
.B1(n_88),
.B2(n_51),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_126),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_22),
.C(n_46),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_15),
.C(n_17),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

AO221x1_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.C(n_40),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_132),
.C(n_137),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_103),
.B(n_11),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_115),
.B1(n_20),
.B2(n_19),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_136),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_141),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_14),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_15),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_147),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_144),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_17),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_18),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_18),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_124),
.C(n_39),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_143),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_156),
.B1(n_158),
.B2(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_165),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_128),
.B1(n_138),
.B2(n_132),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_41),
.C(n_42),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_161),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_168),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_135),
.B(n_138),
.Y(n_168)
);

OAI322xp33_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_174),
.A3(n_177),
.B1(n_149),
.B2(n_154),
.C1(n_153),
.C2(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_133),
.B1(n_134),
.B2(n_48),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_172),
.A2(n_151),
.B1(n_156),
.B2(n_158),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_134),
.B(n_43),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_45),
.Y(n_174)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_134),
.B1(n_166),
.B2(n_153),
.C(n_163),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_181),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_157),
.C(n_161),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_176),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_175),
.B1(n_172),
.B2(n_173),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_188),
.B1(n_184),
.B2(n_183),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_186),
.A2(n_180),
.B(n_181),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_189),
.B(n_169),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_185),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_178),
.B1(n_192),
.B2(n_191),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_196),
.Y(n_197)
);


endmodule