module fake_jpeg_18430_n_209 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_165;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_30),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_12),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_19),
.B1(n_22),
.B2(n_18),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_27),
.B1(n_25),
.B2(n_37),
.Y(n_69)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_44),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_18),
.B1(n_13),
.B2(n_22),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_27),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_13),
.B1(n_22),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_27),
.CON(n_52),
.SN(n_52)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_17),
.B1(n_16),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_59),
.B1(n_64),
.B2(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_55),
.B(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_73),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_17),
.B1(n_16),
.B2(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_20),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_35),
.B1(n_31),
.B2(n_21),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_35),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_37),
.B(n_28),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_37),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_77),
.B(n_88),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_47),
.B(n_50),
.C(n_40),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_43),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_44),
.B1(n_41),
.B2(n_50),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_50),
.B1(n_41),
.B2(n_44),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_91),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_87),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_107),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_69),
.B1(n_72),
.B2(n_71),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_105),
.B1(n_97),
.B2(n_75),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_118),
.B(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_66),
.C(n_63),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_95),
.C(n_80),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_114),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

AO21x2_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_77),
.B(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_121),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_90),
.B(n_94),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_90),
.B(n_94),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_136),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_81),
.B(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_129),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_116),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_107),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_138),
.Y(n_152)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_111),
.C(n_118),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_79),
.B(n_75),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_73),
.B(n_57),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_109),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_27),
.B(n_24),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_147),
.C(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

OA21x2_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_27),
.B(n_24),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_117),
.C(n_101),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_151),
.B1(n_153),
.B2(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_114),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_149),
.A2(n_154),
.B1(n_122),
.B2(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_156),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_127),
.B1(n_120),
.B2(n_124),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_150),
.B(n_121),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_145),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_162),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_108),
.B1(n_120),
.B2(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_161),
.B1(n_141),
.B2(n_140),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_120),
.B1(n_131),
.B2(n_108),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_131),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_167),
.C(n_152),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_172),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_170),
.A2(n_164),
.B1(n_65),
.B2(n_5),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_165),
.B(n_78),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

BUFx4f_ASAP7_75t_SL g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_25),
.B(n_65),
.C(n_78),
.D(n_4),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_0),
.B(n_2),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_2),
.B(n_3),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_166),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_161),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_177),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_191),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_178),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_180),
.B(n_179),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_186),
.B(n_189),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_6),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_3),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_197),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_201),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

AOI321xp33_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_206),
.A3(n_198),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_194),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_11),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_208),
.A2(n_6),
.B(n_10),
.Y(n_209)
);


endmodule