module real_jpeg_41_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_3),
.B(n_11),
.Y(n_10)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_9),
.B1(n_15),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_5),
.A2(n_9),
.B1(n_14),
.B2(n_15),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_19),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_12),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_18),
.Y(n_17)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_9),
.A2(n_15),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_12)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_13),
.B1(n_17),
.B2(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);


endmodule