module fake_jpeg_11568_n_426 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_426);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_65),
.Y(n_106)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_57),
.Y(n_123)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_61),
.Y(n_95)
);

AND2x4_ASAP7_75t_SL g62 ( 
.A(n_34),
.B(n_0),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_66),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_31),
.B(n_8),
.Y(n_65)
);

INVx2_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_70),
.Y(n_116)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_68),
.Y(n_98)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_44),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_0),
.B(n_1),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_80),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_87),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_31),
.B(n_41),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_96),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_39),
.B1(n_33),
.B2(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_97),
.B(n_111),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_53),
.A2(n_39),
.B1(n_20),
.B2(n_33),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_127),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_33),
.B1(n_38),
.B2(n_25),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_38),
.B1(n_36),
.B2(n_42),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_66),
.B(n_41),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_58),
.A2(n_42),
.B1(n_40),
.B2(n_35),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_120),
.B1(n_78),
.B2(n_49),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_40),
.B1(n_35),
.B2(n_29),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_61),
.A2(n_42),
.B1(n_29),
.B2(n_27),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_62),
.B(n_10),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_10),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_144),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_48),
.B1(n_57),
.B2(n_54),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_143),
.A2(n_150),
.B1(n_164),
.B2(n_167),
.Y(n_195)
);

BUFx4f_ASAP7_75t_SL g144 ( 
.A(n_102),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_147),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_55),
.B1(n_56),
.B2(n_69),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_154),
.Y(n_176)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_85),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_85),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_100),
.B(n_1),
.Y(n_158)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_81),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_2),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_91),
.Y(n_163)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_97),
.A2(n_64),
.B1(n_73),
.B2(n_63),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_96),
.B(n_73),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_172),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_110),
.A2(n_63),
.B1(n_12),
.B2(n_4),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_12),
.B1(n_17),
.B2(n_5),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_168),
.A2(n_169),
.B1(n_114),
.B2(n_95),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_105),
.A2(n_123),
.B1(n_128),
.B2(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_123),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_18),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_114),
.B(n_119),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_155),
.B(n_163),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_92),
.C(n_94),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_190),
.C(n_158),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_101),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_124),
.C(n_95),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_108),
.C(n_13),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_151),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_164),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_170),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_201),
.B(n_182),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_205),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_193),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_207),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_148),
.B1(n_139),
.B2(n_170),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_220),
.B1(n_190),
.B2(n_192),
.Y(n_238)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_135),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_224),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_216),
.B(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_222),
.A2(n_223),
.B(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_175),
.B(n_135),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_192),
.B(n_183),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_141),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_228),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_149),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_173),
.B(n_180),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_230),
.A2(n_205),
.B(n_214),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_195),
.B1(n_189),
.B2(n_197),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_231),
.A2(n_235),
.B1(n_250),
.B2(n_249),
.Y(n_271)
);

AOI22x1_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_195),
.B1(n_167),
.B2(n_143),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_238),
.B(n_220),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_203),
.B1(n_208),
.B2(n_227),
.Y(n_235)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_161),
.A3(n_168),
.B1(n_142),
.B2(n_153),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_179),
.Y(n_281)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_246),
.B(n_183),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_137),
.B1(n_136),
.B2(n_140),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_177),
.B1(n_136),
.B2(n_140),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_177),
.B1(n_188),
.B2(n_213),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_179),
.C(n_196),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_224),
.C(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_257),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_262),
.C(n_280),
.Y(n_289)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_206),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_261),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_215),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_265),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_207),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_238),
.A2(n_220),
.B(n_202),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_276),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_270),
.B1(n_279),
.B2(n_284),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_218),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_233),
.A2(n_225),
.B1(n_219),
.B2(n_210),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_271),
.A2(n_275),
.B1(n_281),
.B2(n_236),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_245),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_231),
.A2(n_209),
.B1(n_222),
.B2(n_223),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_234),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_255),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_232),
.A2(n_254),
.B1(n_235),
.B2(n_248),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_217),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_232),
.A2(n_200),
.B(n_191),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_286),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_243),
.B1(n_244),
.B2(n_196),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_241),
.A2(n_200),
.B(n_191),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_237),
.B1(n_251),
.B2(n_252),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_287),
.A2(n_299),
.B1(n_281),
.B2(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_242),
.C(n_251),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_297),
.C(n_256),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_252),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_304),
.Y(n_317)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_296),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_250),
.C(n_166),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_236),
.B1(n_213),
.B2(n_177),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_298),
.A2(n_107),
.B1(n_145),
.B2(n_93),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_280),
.B(n_159),
.CI(n_144),
.CON(n_302),
.SN(n_302)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_302),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_171),
.Y(n_304)
);

XOR2x2_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_98),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_306),
.A2(n_276),
.B(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_286),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_314),
.Y(n_354)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_274),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_316),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_261),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_322),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_284),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_320),
.B(n_332),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_273),
.B1(n_269),
.B2(n_263),
.Y(n_321)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_321),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_257),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_293),
.B(n_269),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_323),
.B(n_330),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_327),
.C(n_331),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_300),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_326),
.A2(n_309),
.B(n_329),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_275),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_295),
.A2(n_272),
.B1(n_181),
.B2(n_188),
.Y(n_328)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_290),
.B(n_272),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_98),
.C(n_89),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_301),
.B(n_308),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_291),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_313),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_181),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_334),
.B(n_335),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_88),
.C(n_89),
.Y(n_335)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_336),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_309),
.B(n_306),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_338),
.A2(n_340),
.B(n_346),
.Y(n_358)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

AO221x1_ASAP7_75t_L g340 ( 
.A1(n_325),
.A2(n_294),
.B1(n_311),
.B2(n_303),
.C(n_312),
.Y(n_340)
);

INVx13_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_318),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_327),
.A2(n_288),
.B1(n_302),
.B2(n_300),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_12),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_17),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_349),
.B(n_8),
.Y(n_369)
);

OA21x2_ASAP7_75t_L g355 ( 
.A1(n_328),
.A2(n_88),
.B(n_144),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_SL g365 ( 
.A1(n_355),
.A2(n_144),
.B(n_159),
.C(n_107),
.Y(n_365)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_352),
.B(n_330),
.C(n_345),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_359),
.B(n_351),
.Y(n_386)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_352),
.B(n_345),
.C(n_322),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_373),
.Y(n_377)
);

OAI221xp5_ASAP7_75t_L g362 ( 
.A1(n_354),
.A2(n_317),
.B1(n_323),
.B2(n_331),
.C(n_6),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_362),
.A2(n_366),
.B1(n_350),
.B2(n_342),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_357),
.Y(n_364)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

AOI21x1_ASAP7_75t_L g381 ( 
.A1(n_365),
.A2(n_355),
.B(n_338),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_337),
.A2(n_317),
.B1(n_131),
.B2(n_128),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_357),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_367),
.B(n_346),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_14),
.C(n_16),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_371),
.C(n_341),
.Y(n_387)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_104),
.C(n_119),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_121),
.C(n_8),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_7),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_374),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_383),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_SL g380 ( 
.A(n_361),
.B(n_348),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_384),
.Y(n_394)
);

AOI21x1_ASAP7_75t_SL g393 ( 
.A1(n_381),
.A2(n_365),
.B(n_363),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_388),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_341),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_386),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_387),
.B(n_368),
.C(n_355),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_342),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_351),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_121),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_373),
.C(n_353),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_397),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_376),
.A2(n_340),
.B(n_353),
.Y(n_391)
);

OAI21x1_ASAP7_75t_L g410 ( 
.A1(n_391),
.A2(n_393),
.B(n_398),
.Y(n_410)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_365),
.C(n_344),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_380),
.A2(n_363),
.B(n_365),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_363),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_5),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_387),
.Y(n_401)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_401),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_381),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_403),
.B(n_404),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_399),
.B(n_14),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_407),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_6),
.B(n_15),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_390),
.C(n_15),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_6),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_409),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_402),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_411),
.A2(n_15),
.B(n_18),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_401),
.A2(n_393),
.B(n_389),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_414),
.A2(n_406),
.B(n_410),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_3),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_418),
.A2(n_419),
.B(n_420),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_417),
.B(n_18),
.C(n_2),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_421),
.Y(n_422)
);

OAI321xp33_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_412),
.A3(n_414),
.B1(n_415),
.B2(n_413),
.C(n_3),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_424),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_422),
.Y(n_426)
);


endmodule