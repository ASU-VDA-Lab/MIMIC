module real_aes_6580_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_0), .B(n_84), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g457 ( .A(n_0), .Y(n_457) );
INVx1_ASAP7_75t_L g508 ( .A(n_1), .Y(n_508) );
INVx1_ASAP7_75t_L g203 ( .A(n_2), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_3), .A2(n_77), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_3), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_4), .A2(n_38), .B1(n_159), .B2(n_524), .Y(n_534) );
AOI21xp33_ASAP7_75t_L g183 ( .A1(n_5), .A2(n_140), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_6), .B(n_133), .Y(n_499) );
AND2x6_ASAP7_75t_L g145 ( .A(n_7), .B(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_8), .A2(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_9), .B(n_39), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_10), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g190 ( .A(n_11), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_12), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g503 ( .A(n_13), .Y(n_503) );
INVx1_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
INVx1_ASAP7_75t_L g248 ( .A(n_15), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_16), .B(n_171), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_17), .B(n_134), .Y(n_480) );
AO32x2_ASAP7_75t_L g532 ( .A1(n_18), .A2(n_133), .A3(n_168), .B1(n_486), .B2(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_19), .B(n_159), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_20), .B(n_154), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_21), .B(n_134), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_22), .A2(n_50), .B1(n_159), .B2(n_524), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_23), .B(n_140), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_24), .A2(n_74), .B1(n_159), .B2(n_171), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_25), .B(n_159), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_26), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_27), .A2(n_246), .B(n_247), .C(n_249), .Y(n_245) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_28), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_29), .B(n_192), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_30), .B(n_188), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_31), .A2(n_42), .B1(n_751), .B2(n_752), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_31), .Y(n_751) );
INVx1_ASAP7_75t_L g177 ( .A(n_32), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_33), .B(n_192), .Y(n_547) );
INVx2_ASAP7_75t_L g143 ( .A(n_34), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_35), .B(n_159), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_36), .B(n_192), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_37), .A2(n_145), .B(n_149), .C(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_39), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g175 ( .A(n_40), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_41), .B(n_188), .Y(n_258) );
CKINVDCx14_ASAP7_75t_R g752 ( .A(n_42), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_43), .B(n_159), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_44), .A2(n_85), .B1(n_221), .B2(n_524), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_45), .B(n_159), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_46), .B(n_159), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_47), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_48), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_49), .B(n_140), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_51), .A2(n_60), .B1(n_159), .B2(n_171), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_52), .A2(n_149), .B1(n_171), .B2(n_173), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_53), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_54), .B(n_159), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_55), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_56), .B(n_159), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_57), .A2(n_158), .B(n_187), .C(n_189), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_58), .Y(n_262) );
INVx1_ASAP7_75t_L g185 ( .A(n_59), .Y(n_185) );
INVx1_ASAP7_75t_L g146 ( .A(n_61), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_62), .B(n_159), .Y(n_509) );
INVx1_ASAP7_75t_L g137 ( .A(n_63), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_64), .Y(n_118) );
AO32x2_ASAP7_75t_L g527 ( .A1(n_65), .A2(n_133), .A3(n_228), .B1(n_486), .B2(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g566 ( .A(n_66), .Y(n_566) );
INVx1_ASAP7_75t_L g542 ( .A(n_67), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_SL g153 ( .A1(n_68), .A2(n_154), .B(n_155), .C(n_158), .Y(n_153) );
INVxp67_ASAP7_75t_L g156 ( .A(n_69), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_70), .B(n_171), .Y(n_543) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_72), .Y(n_181) );
INVx1_ASAP7_75t_L g255 ( .A(n_73), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_75), .A2(n_145), .B(n_149), .C(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_76), .B(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_77), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_78), .B(n_171), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_79), .B(n_204), .Y(n_217) );
INVx2_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_81), .B(n_154), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_82), .B(n_171), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_83), .A2(n_145), .B(n_149), .C(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g454 ( .A(n_84), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g467 ( .A(n_84), .B(n_456), .Y(n_467) );
INVx2_ASAP7_75t_L g471 ( .A(n_84), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_86), .A2(n_100), .B1(n_171), .B2(n_172), .Y(n_483) );
AOI222xp33_ASAP7_75t_L g463 ( .A1(n_87), .A2(n_464), .B1(n_750), .B2(n_753), .C1(n_755), .C2(n_756), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_88), .B(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_89), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_90), .A2(n_145), .B(n_149), .C(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_91), .Y(n_238) );
INVx1_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_93), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_94), .B(n_204), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_95), .B(n_171), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_96), .B(n_133), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_97), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_98), .A2(n_140), .B(n_147), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_99), .A2(n_102), .B1(n_105), .B2(n_113), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_462), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g760 ( .A(n_117), .Y(n_760) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_451), .B(n_459), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_125), .B2(n_450), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g450 ( .A(n_125), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_125), .A2(n_465), .B1(n_468), .B2(n_472), .Y(n_464) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_387), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_317), .C(n_348), .D(n_367), .Y(n_126) );
NAND4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_275), .C(n_290), .D(n_308), .Y(n_127) );
AOI222xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_210), .B1(n_251), .B2(n_263), .C1(n_268), .C2(n_270), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_193), .Y(n_129) );
INVx1_ASAP7_75t_L g331 ( .A(n_130), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_164), .Y(n_130) );
AND2x2_ASAP7_75t_L g194 ( .A(n_131), .B(n_182), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_131), .B(n_197), .Y(n_360) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g267 ( .A(n_132), .B(n_166), .Y(n_267) );
AND2x2_ASAP7_75t_L g276 ( .A(n_132), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g302 ( .A(n_132), .Y(n_302) );
AND2x2_ASAP7_75t_L g323 ( .A(n_132), .B(n_166), .Y(n_323) );
BUFx2_ASAP7_75t_L g346 ( .A(n_132), .Y(n_346) );
AND2x2_ASAP7_75t_L g370 ( .A(n_132), .B(n_167), .Y(n_370) );
AND2x2_ASAP7_75t_L g434 ( .A(n_132), .B(n_182), .Y(n_434) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B(n_161), .Y(n_132) );
INVx4_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_133), .A2(n_491), .B(n_499), .Y(n_490) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_135), .B(n_136), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g242 ( .A(n_140), .Y(n_242) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_141), .B(n_145), .Y(n_179) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g498 ( .A(n_142), .Y(n_498) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g150 ( .A(n_143), .Y(n_150) );
INVx1_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
INVx1_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
INVx1_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
INVx3_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_144), .Y(n_188) );
INVx4_ASAP7_75t_SL g160 ( .A(n_145), .Y(n_160) );
BUFx3_ASAP7_75t_L g486 ( .A(n_145), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_145), .A2(n_492), .B(n_495), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_145), .A2(n_502), .B(n_506), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_145), .A2(n_517), .B(n_521), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_145), .A2(n_541), .B(n_544), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B(n_153), .C(n_160), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_148), .A2(n_160), .B(n_185), .C(n_186), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_148), .A2(n_160), .B(n_244), .C(n_245), .Y(n_243) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx3_ASAP7_75t_L g221 ( .A(n_150), .Y(n_221) );
INVx1_ASAP7_75t_L g524 ( .A(n_150), .Y(n_524) );
INVx1_ASAP7_75t_L g520 ( .A(n_154), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_157), .B(n_190), .Y(n_189) );
INVx5_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
OAI22xp5_ASAP7_75t_SL g528 ( .A1(n_157), .A2(n_188), .B1(n_529), .B2(n_530), .Y(n_528) );
O2A1O1Ixp5_ASAP7_75t_SL g541 ( .A1(n_158), .A2(n_204), .B(n_542), .C(n_543), .Y(n_541) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_159), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g169 ( .A1(n_160), .A2(n_170), .B1(n_178), .B2(n_179), .Y(n_169) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_162), .A2(n_183), .B(n_191), .Y(n_182) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g223 ( .A(n_163), .B(n_224), .Y(n_223) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_163), .B(n_482), .C(n_486), .Y(n_481) );
AO21x1_ASAP7_75t_L g574 ( .A1(n_163), .A2(n_482), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g335 ( .A(n_164), .B(n_266), .Y(n_335) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_165), .B(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_182), .Y(n_165) );
OR2x2_ASAP7_75t_L g295 ( .A(n_166), .B(n_198), .Y(n_295) );
AND2x2_ASAP7_75t_L g307 ( .A(n_166), .B(n_266), .Y(n_307) );
BUFx2_ASAP7_75t_L g439 ( .A(n_166), .Y(n_439) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OR2x2_ASAP7_75t_L g196 ( .A(n_167), .B(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g289 ( .A(n_167), .B(n_198), .Y(n_289) );
AND2x2_ASAP7_75t_L g342 ( .A(n_167), .B(n_182), .Y(n_342) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_167), .Y(n_378) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_180), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_168), .B(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_168), .A2(n_199), .B(n_207), .Y(n_198) );
INVx2_ASAP7_75t_L g222 ( .A(n_168), .Y(n_222) );
INVx2_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_173) );
INVx2_ASAP7_75t_L g176 ( .A(n_174), .Y(n_176) );
INVx4_ASAP7_75t_L g246 ( .A(n_174), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_179), .A2(n_200), .B(n_201), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_179), .A2(n_255), .B(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g265 ( .A(n_182), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_SL g277 ( .A(n_182), .Y(n_277) );
INVx2_ASAP7_75t_L g288 ( .A(n_182), .Y(n_288) );
BUFx2_ASAP7_75t_L g312 ( .A(n_182), .Y(n_312) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_182), .B(n_370), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_187), .A2(n_522), .B(n_523), .Y(n_521) );
O2A1O1Ixp5_ASAP7_75t_L g565 ( .A1(n_187), .A2(n_507), .B(n_566), .C(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx4_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_188), .A2(n_483), .B1(n_484), .B2(n_485), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_188), .A2(n_484), .B1(n_534), .B2(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g209 ( .A(n_192), .Y(n_209) );
INVx2_ASAP7_75t_L g228 ( .A(n_192), .Y(n_228) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_192), .A2(n_241), .B(n_250), .Y(n_240) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_192), .A2(n_516), .B(n_525), .Y(n_515) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_192), .A2(n_540), .B(n_547), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AOI332xp33_ASAP7_75t_L g290 ( .A1(n_194), .A2(n_291), .A3(n_295), .B1(n_296), .B2(n_300), .B3(n_303), .C1(n_304), .C2(n_306), .Y(n_290) );
NAND2x1_ASAP7_75t_L g375 ( .A(n_194), .B(n_266), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_194), .B(n_280), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_SL g308 ( .A1(n_195), .A2(n_309), .B(n_312), .C(n_313), .Y(n_308) );
AND2x2_ASAP7_75t_L g447 ( .A(n_195), .B(n_288), .Y(n_447) );
INVx3_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g344 ( .A(n_196), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g349 ( .A(n_196), .B(n_346), .Y(n_349) );
INVx1_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
AND2x2_ASAP7_75t_L g383 ( .A(n_197), .B(n_342), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_197), .B(n_323), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_197), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_197), .B(n_301), .Y(n_409) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g266 ( .A(n_198), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .C(n_206), .Y(n_202) );
INVx2_ASAP7_75t_L g484 ( .A(n_204), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_204), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_204), .A2(n_563), .B(n_564), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_206), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_209), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_209), .B(n_262), .Y(n_261) );
OAI31xp33_ASAP7_75t_L g448 ( .A1(n_210), .A2(n_369), .A3(n_376), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_225), .Y(n_210) );
AND2x2_ASAP7_75t_L g251 ( .A(n_211), .B(n_252), .Y(n_251) );
NAND2x1_ASAP7_75t_SL g271 ( .A(n_211), .B(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_211), .Y(n_358) );
AND2x2_ASAP7_75t_L g363 ( .A(n_211), .B(n_274), .Y(n_363) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_212), .A2(n_276), .B(n_278), .C(n_281), .Y(n_275) );
OR2x2_ASAP7_75t_L g292 ( .A(n_212), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g305 ( .A(n_212), .Y(n_305) );
AND2x2_ASAP7_75t_L g311 ( .A(n_212), .B(n_253), .Y(n_311) );
INVx2_ASAP7_75t_L g329 ( .A(n_212), .Y(n_329) );
AND2x2_ASAP7_75t_L g340 ( .A(n_212), .B(n_294), .Y(n_340) );
AND2x2_ASAP7_75t_L g372 ( .A(n_212), .B(n_330), .Y(n_372) );
AND2x2_ASAP7_75t_L g376 ( .A(n_212), .B(n_299), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_212), .B(n_225), .Y(n_381) );
AND2x2_ASAP7_75t_L g415 ( .A(n_212), .B(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_212), .B(n_318), .Y(n_449) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
AOI21xp5_ASAP7_75t_SL g213 ( .A1(n_214), .A2(n_215), .B(n_222), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_219), .A2(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
INVx1_ASAP7_75t_L g260 ( .A(n_222), .Y(n_260) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_222), .A2(n_501), .B(n_510), .Y(n_500) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_222), .A2(n_561), .B(n_568), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_225), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g357 ( .A(n_225), .Y(n_357) );
AND2x2_ASAP7_75t_L g419 ( .A(n_225), .B(n_340), .Y(n_419) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
OR2x2_ASAP7_75t_L g273 ( .A(n_226), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g283 ( .A(n_226), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_226), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g391 ( .A(n_226), .Y(n_391) );
AND2x2_ASAP7_75t_L g408 ( .A(n_226), .B(n_253), .Y(n_408) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g299 ( .A(n_227), .B(n_239), .Y(n_299) );
AND2x2_ASAP7_75t_L g328 ( .A(n_227), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g339 ( .A(n_227), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_227), .B(n_294), .Y(n_430) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_235), .Y(n_231) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g252 ( .A(n_240), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g274 ( .A(n_240), .Y(n_274) );
AND2x2_ASAP7_75t_L g330 ( .A(n_240), .B(n_294), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_246), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g505 ( .A(n_246), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_246), .A2(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g432 ( .A(n_251), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_252), .Y(n_436) );
INVx2_ASAP7_75t_L g294 ( .A(n_253), .Y(n_294) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_260), .B(n_261), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_265), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_265), .B(n_370), .Y(n_428) );
OR2x2_ASAP7_75t_L g269 ( .A(n_266), .B(n_267), .Y(n_269) );
INVx1_ASAP7_75t_SL g321 ( .A(n_266), .Y(n_321) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_272), .A2(n_325), .B1(n_327), .B2(n_331), .C(n_332), .Y(n_324) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g352 ( .A(n_273), .B(n_316), .Y(n_352) );
INVx2_ASAP7_75t_L g284 ( .A(n_274), .Y(n_284) );
INVx1_ASAP7_75t_L g310 ( .A(n_274), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_274), .B(n_294), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_274), .B(n_297), .Y(n_404) );
INVx1_ASAP7_75t_L g412 ( .A(n_274), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_276), .B(n_280), .Y(n_326) );
AND2x4_ASAP7_75t_L g301 ( .A(n_277), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g414 ( .A(n_280), .B(n_370), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_283), .B(n_315), .Y(n_314) );
INVxp67_ASAP7_75t_L g422 ( .A(n_284), .Y(n_422) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g322 ( .A(n_288), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g394 ( .A(n_288), .B(n_370), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_288), .B(n_307), .Y(n_400) );
AOI322xp5_ASAP7_75t_L g354 ( .A1(n_289), .A2(n_323), .A3(n_330), .B1(n_355), .B2(n_358), .C1(n_359), .C2(n_361), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_289), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g420 ( .A(n_292), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g366 ( .A(n_293), .Y(n_366) );
INVx2_ASAP7_75t_L g297 ( .A(n_294), .Y(n_297) );
INVx1_ASAP7_75t_L g356 ( .A(n_294), .Y(n_356) );
CKINVDCx16_ASAP7_75t_R g303 ( .A(n_295), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g392 ( .A(n_297), .B(n_305), .Y(n_392) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_299), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g347 ( .A(n_299), .B(n_340), .Y(n_347) );
AND2x2_ASAP7_75t_L g351 ( .A(n_299), .B(n_311), .Y(n_351) );
OAI21xp33_ASAP7_75t_SL g361 ( .A1(n_300), .A2(n_362), .B(n_364), .Y(n_361) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_300), .A2(n_432), .B1(n_433), .B2(n_435), .Y(n_431) );
INVx3_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g306 ( .A(n_301), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_301), .B(n_321), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_303), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g443 ( .A(n_310), .Y(n_443) );
INVx4_ASAP7_75t_L g316 ( .A(n_311), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_311), .B(n_338), .Y(n_386) );
INVx1_ASAP7_75t_SL g398 ( .A(n_312), .Y(n_398) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp67_ASAP7_75t_L g411 ( .A(n_316), .B(n_412), .Y(n_411) );
OAI211xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_319), .B(n_324), .C(n_341), .Y(n_317) );
OAI221xp5_ASAP7_75t_SL g437 ( .A1(n_319), .A2(n_357), .B1(n_436), .B2(n_438), .C(n_440), .Y(n_437) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_321), .B(n_434), .Y(n_433) );
OAI31xp33_ASAP7_75t_L g413 ( .A1(n_322), .A2(n_399), .A3(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g353 ( .A(n_323), .Y(n_353) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g403 ( .A(n_328), .Y(n_403) );
AND2x2_ASAP7_75t_L g416 ( .A(n_330), .B(n_339), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B(n_336), .Y(n_332) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_340), .B(n_443), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI221xp5_ASAP7_75t_SL g348 ( .A1(n_349), .A2(n_350), .B1(n_352), .B2(n_353), .C(n_354), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_349), .A2(n_418), .B(n_420), .C(n_423), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_352), .B(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g379 ( .A(n_360), .Y(n_379) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g365 ( .A(n_363), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g407 ( .A(n_363), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B(n_373), .C(n_382), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g444 ( .A1(n_371), .A2(n_381), .B1(n_445), .B2(n_446), .C(n_448), .Y(n_444) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B1(n_377), .B2(n_380), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_384), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_SL g445 ( .A(n_384), .Y(n_445) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR4xp25_ASAP7_75t_L g387 ( .A(n_388), .B(n_417), .C(n_437), .D(n_444), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_393), .B(n_395), .C(n_413), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .B(n_401), .C(n_405), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g424 ( .A(n_402), .Y(n_424) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
OR2x2_ASAP7_75t_L g435 ( .A(n_403), .B(n_436), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_427), .B2(n_429), .C(n_431), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_434), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22x1_ASAP7_75t_SL g753 ( .A1(n_450), .A2(n_470), .B1(n_473), .B2(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_454), .Y(n_461) );
NOR2x2_ASAP7_75t_L g758 ( .A(n_455), .B(n_471), .Y(n_758) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g470 ( .A(n_456), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_459), .B(n_463), .C(n_759), .Y(n_462) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g754 ( .A(n_466), .Y(n_754) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_475), .B(n_684), .Y(n_474) );
NOR5xp2_ASAP7_75t_L g475 ( .A(n_476), .B(n_597), .C(n_643), .D(n_656), .E(n_668), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_511), .B(n_551), .C(n_578), .Y(n_476) );
INVx1_ASAP7_75t_SL g679 ( .A(n_477), .Y(n_679) );
OR2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_487), .Y(n_477) );
AND2x2_ASAP7_75t_L g603 ( .A(n_478), .B(n_488), .Y(n_603) );
AND2x2_ASAP7_75t_L g631 ( .A(n_478), .B(n_577), .Y(n_631) );
AND2x2_ASAP7_75t_L g639 ( .A(n_478), .B(n_582), .Y(n_639) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g569 ( .A(n_479), .B(n_489), .Y(n_569) );
INVx2_ASAP7_75t_L g581 ( .A(n_479), .Y(n_581) );
AND2x2_ASAP7_75t_L g706 ( .A(n_479), .B(n_648), .Y(n_706) );
OR2x2_ASAP7_75t_L g708 ( .A(n_479), .B(n_709), .Y(n_708) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g575 ( .A(n_480), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_484), .A2(n_496), .B(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_484), .A2(n_507), .B(n_508), .C(n_509), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_486), .A2(n_562), .B(n_565), .Y(n_561) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g619 ( .A(n_488), .B(n_591), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_488), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g733 ( .A(n_488), .B(n_573), .Y(n_733) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_500), .Y(n_488) );
AND2x2_ASAP7_75t_L g576 ( .A(n_489), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g623 ( .A(n_489), .Y(n_623) );
AND2x2_ASAP7_75t_L g648 ( .A(n_489), .B(n_560), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_489), .B(n_681), .Y(n_718) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g582 ( .A(n_490), .B(n_560), .Y(n_582) );
AND2x2_ASAP7_75t_L g596 ( .A(n_490), .B(n_559), .Y(n_596) );
AND2x2_ASAP7_75t_L g613 ( .A(n_490), .B(n_500), .Y(n_613) );
AND2x2_ASAP7_75t_L g670 ( .A(n_490), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_490), .B(n_577), .Y(n_683) );
AND2x2_ASAP7_75t_L g735 ( .A(n_490), .B(n_660), .Y(n_735) );
INVx2_ASAP7_75t_L g507 ( .A(n_498), .Y(n_507) );
AND2x2_ASAP7_75t_L g558 ( .A(n_500), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g577 ( .A(n_500), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_500), .B(n_560), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_536), .B(n_548), .Y(n_511) );
INVx1_ASAP7_75t_SL g667 ( .A(n_512), .Y(n_667) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_526), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_SL g555 ( .A(n_514), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g550 ( .A(n_515), .Y(n_550) );
INVx1_ASAP7_75t_L g587 ( .A(n_515), .Y(n_587) );
AND2x2_ASAP7_75t_L g608 ( .A(n_515), .B(n_531), .Y(n_608) );
AND2x2_ASAP7_75t_L g642 ( .A(n_515), .B(n_532), .Y(n_642) );
OR2x2_ASAP7_75t_L g661 ( .A(n_515), .B(n_538), .Y(n_661) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_515), .Y(n_675) );
AND2x2_ASAP7_75t_L g688 ( .A(n_515), .B(n_689), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_526), .A2(n_610), .B1(n_611), .B2(n_620), .Y(n_609) );
AND2x2_ASAP7_75t_L g693 ( .A(n_526), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
INVx1_ASAP7_75t_L g554 ( .A(n_527), .Y(n_554) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_527), .Y(n_591) );
INVx1_ASAP7_75t_L g602 ( .A(n_527), .Y(n_602) );
AND2x2_ASAP7_75t_L g617 ( .A(n_527), .B(n_532), .Y(n_617) );
OR2x2_ASAP7_75t_L g571 ( .A(n_531), .B(n_556), .Y(n_571) );
AND2x2_ASAP7_75t_L g601 ( .A(n_531), .B(n_602), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_531), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g549 ( .A(n_532), .B(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g658 ( .A(n_532), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_536), .B(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g636 ( .A(n_537), .B(n_602), .Y(n_636) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g548 ( .A(n_538), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g556 ( .A(n_539), .Y(n_556) );
OR2x2_ASAP7_75t_L g586 ( .A(n_539), .B(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_539), .Y(n_641) );
AOI32xp33_ASAP7_75t_L g678 ( .A1(n_548), .A2(n_608), .A3(n_679), .B1(n_680), .B2(n_682), .Y(n_678) );
AND2x2_ASAP7_75t_L g604 ( .A(n_549), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_549), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_549), .B(n_636), .Y(n_722) );
INVx1_ASAP7_75t_L g727 ( .A(n_549), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_557), .B1(n_570), .B2(n_572), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
AND2x2_ASAP7_75t_L g657 ( .A(n_553), .B(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_554), .B(n_556), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_555), .A2(n_579), .B1(n_583), .B2(n_593), .Y(n_578) );
AND2x2_ASAP7_75t_L g600 ( .A(n_555), .B(n_601), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g651 ( .A1(n_555), .A2(n_569), .B(n_617), .C(n_652), .Y(n_651) );
OAI332xp33_ASAP7_75t_L g656 ( .A1(n_555), .A2(n_657), .A3(n_659), .B1(n_661), .B2(n_662), .B3(n_664), .C1(n_665), .C2(n_667), .Y(n_656) );
INVx2_ASAP7_75t_L g697 ( .A(n_555), .Y(n_697) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_556), .Y(n_615) );
INVx1_ASAP7_75t_L g690 ( .A(n_556), .Y(n_690) );
AND2x2_ASAP7_75t_L g744 ( .A(n_556), .B(n_608), .Y(n_744) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_569), .Y(n_557) );
AND2x2_ASAP7_75t_L g624 ( .A(n_559), .B(n_574), .Y(n_624) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g573 ( .A(n_560), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g672 ( .A(n_560), .B(n_574), .Y(n_672) );
INVx1_ASAP7_75t_L g681 ( .A(n_560), .Y(n_681) );
INVx1_ASAP7_75t_L g655 ( .A(n_569), .Y(n_655) );
INVxp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g739 ( .A(n_571), .B(n_591), .Y(n_739) );
INVx1_ASAP7_75t_SL g650 ( .A(n_572), .Y(n_650) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
AND2x2_ASAP7_75t_L g677 ( .A(n_573), .B(n_635), .Y(n_677) );
INVx1_ASAP7_75t_L g696 ( .A(n_573), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_573), .B(n_663), .Y(n_698) );
INVx1_ASAP7_75t_L g595 ( .A(n_574), .Y(n_595) );
AND2x2_ASAP7_75t_L g599 ( .A(n_576), .B(n_580), .Y(n_599) );
AND2x2_ASAP7_75t_L g666 ( .A(n_576), .B(n_624), .Y(n_666) );
INVx2_ASAP7_75t_L g709 ( .A(n_576), .Y(n_709) );
INVx2_ASAP7_75t_L g592 ( .A(n_577), .Y(n_592) );
AND2x2_ASAP7_75t_L g594 ( .A(n_577), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g610 ( .A(n_580), .Y(n_610) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_581), .B(n_654), .Y(n_660) );
OR2x2_ASAP7_75t_L g724 ( .A(n_581), .B(n_683), .Y(n_724) );
INVx1_ASAP7_75t_L g748 ( .A(n_581), .Y(n_748) );
INVx1_ASAP7_75t_L g704 ( .A(n_582), .Y(n_704) );
AND2x2_ASAP7_75t_L g749 ( .A(n_582), .B(n_592), .Y(n_749) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_586), .A2(n_612), .B1(n_614), .B2(n_618), .Y(n_611) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI322xp33_ASAP7_75t_SL g695 ( .A1(n_589), .A2(n_696), .A3(n_697), .B1(n_698), .B2(n_699), .C1(n_702), .C2(n_704), .Y(n_695) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
AND2x2_ASAP7_75t_L g692 ( .A(n_590), .B(n_608), .Y(n_692) );
OR2x2_ASAP7_75t_L g726 ( .A(n_590), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g729 ( .A(n_590), .B(n_661), .Y(n_729) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g674 ( .A(n_591), .B(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g730 ( .A(n_591), .B(n_661), .Y(n_730) );
INVx3_ASAP7_75t_L g663 ( .A(n_592), .Y(n_663) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx1_ASAP7_75t_L g719 ( .A(n_594), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g598 ( .A1(n_596), .A2(n_599), .B1(n_600), .B2(n_603), .C1(n_604), .C2(n_606), .Y(n_598) );
INVx1_ASAP7_75t_L g629 ( .A(n_596), .Y(n_629) );
NAND3xp33_ASAP7_75t_SL g597 ( .A(n_598), .B(n_609), .C(n_626), .Y(n_597) );
AND2x2_ASAP7_75t_L g714 ( .A(n_601), .B(n_615), .Y(n_714) );
BUFx2_ASAP7_75t_L g605 ( .A(n_602), .Y(n_605) );
INVx1_ASAP7_75t_L g646 ( .A(n_602), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_603), .A2(n_639), .B1(n_692), .B2(n_693), .C(n_695), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_605), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_608), .Y(n_632) );
AND2x2_ASAP7_75t_L g645 ( .A(n_608), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_613), .B(n_624), .Y(n_625) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g620 ( .A1(n_615), .A2(n_621), .B(n_625), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_615), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g712 ( .A(n_617), .B(n_694), .Y(n_712) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g635 ( .A(n_623), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_624), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g741 ( .A(n_624), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_632), .B1(n_633), .B2(n_636), .C(n_637), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_628), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g737 ( .A(n_636), .B(n_642), .Y(n_737) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OAI31xp33_ASAP7_75t_SL g705 ( .A1(n_640), .A2(n_679), .A3(n_706), .B(n_707), .Y(n_705) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g694 ( .A(n_641), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_642), .B(n_646), .Y(n_745) );
OAI221xp5_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_647), .B1(n_649), .B2(n_650), .C(n_651), .Y(n_643) );
INVx1_ASAP7_75t_L g649 ( .A(n_645), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_648), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g664 ( .A(n_657), .Y(n_664) );
INVx2_ASAP7_75t_L g700 ( .A(n_658), .Y(n_700) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g686 ( .A(n_663), .B(n_672), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_663), .A2(n_680), .B(n_737), .C(n_738), .Y(n_736) );
OAI221xp5_ASAP7_75t_SL g668 ( .A1(n_664), .A2(n_669), .B1(n_673), .B2(n_676), .C(n_678), .Y(n_668) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_L g731 ( .A1(n_667), .A2(n_732), .B(n_734), .C(n_736), .Y(n_731) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_670), .A2(n_721), .B1(n_723), .B2(n_725), .C(n_728), .Y(n_720) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
NOR4xp25_ASAP7_75t_L g684 ( .A(n_685), .B(n_710), .C(n_731), .D(n_742), .Y(n_684) );
OAI211xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_687), .B(n_691), .C(n_705), .Y(n_685) );
INVx1_ASAP7_75t_SL g740 ( .A(n_692), .Y(n_740) );
OR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_SL g703 ( .A(n_701), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_708), .A2(n_717), .B1(n_729), .B2(n_730), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_713), .B(n_715), .C(n_720), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI31xp33_ASAP7_75t_L g742 ( .A1(n_713), .A2(n_743), .A3(n_745), .B(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g755 ( .A(n_750), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
endmodule