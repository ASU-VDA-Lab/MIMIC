module fake_ariane_701_n_76 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_32, n_28, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_33, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_76);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_32;
input n_28;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_33;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_76;

wire n_56;
wire n_60;
wire n_48;
wire n_64;
wire n_38;
wire n_47;
wire n_58;
wire n_37;
wire n_65;
wire n_75;
wire n_67;
wire n_45;
wire n_69;
wire n_52;
wire n_74;
wire n_73;
wire n_40;
wire n_53;
wire n_61;
wire n_66;
wire n_71;
wire n_43;
wire n_49;
wire n_41;
wire n_50;
wire n_55;
wire n_62;
wire n_51;
wire n_46;
wire n_36;
wire n_68;
wire n_72;
wire n_44;
wire n_39;
wire n_63;
wire n_59;
wire n_42;
wire n_57;
wire n_70;
wire n_35;
wire n_54;

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_28),
.Y(n_39)
);

NOR2xp67_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_26),
.A2(n_18),
.B1(n_10),
.B2(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_4),
.C(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

OAI21x1_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_35),
.B(n_47),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_49),
.Y(n_60)
);

OAI21x1_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_48),
.B(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_42),
.B(n_41),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_54),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_40),
.C(n_37),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

OAI221xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_57),
.B1(n_69),
.B2(n_71),
.C(n_55),
.Y(n_73)
);

NAND4xp25_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_39),
.C(n_46),
.D(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_14),
.A3(n_20),
.B1(n_27),
.B2(n_29),
.C1(n_30),
.C2(n_31),
.Y(n_76)
);


endmodule