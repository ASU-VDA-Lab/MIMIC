module fake_jpeg_13178_n_185 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_73),
.Y(n_85)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_47),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_69),
.B1(n_65),
.B2(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_95),
.B1(n_97),
.B2(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_52),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_53),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_66),
.B1(n_62),
.B2(n_61),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_57),
.B1(n_45),
.B2(n_59),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_109),
.B1(n_116),
.B2(n_70),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_50),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_54),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_59),
.B(n_58),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_116),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_58),
.B1(n_54),
.B2(n_55),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_1),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_1),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_2),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_112),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_13),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_141),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_3),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_139),
.B(n_142),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_70),
.C(n_49),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_127),
.C(n_128),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_5),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_122),
.B(n_137),
.C(n_138),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_44),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_155),
.Y(n_170)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_149),
.B(n_22),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_43),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_122),
.Y(n_153)
);

CKINVDCx11_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_157),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_14),
.B(n_18),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_19),
.B(n_21),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_150),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_159),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_169),
.C(n_24),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_23),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_39),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_151),
.B1(n_160),
.B2(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_174),
.Y(n_176)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_144),
.B(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_173),
.Y(n_177)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_168),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_172),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_176),
.B(n_170),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_163),
.B(n_164),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_163),
.B(n_175),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_25),
.C(n_27),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_184),
.Y(n_185)
);


endmodule