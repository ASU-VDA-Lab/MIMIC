module fake_jpeg_28915_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx12f_ASAP7_75t_SL g40 ( 
.A(n_21),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_42),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_24),
.B1(n_22),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_50),
.A2(n_41),
.B1(n_33),
.B2(n_32),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_46),
.B1(n_22),
.B2(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_52),
.A2(n_62),
.B1(n_63),
.B2(n_21),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_36),
.B1(n_29),
.B2(n_22),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_33),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_35),
.B1(n_23),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_66),
.B1(n_69),
.B2(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_17),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_46),
.B1(n_24),
.B2(n_37),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_35),
.B1(n_23),
.B2(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_35),
.B1(n_23),
.B2(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_71),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_17),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_38),
.A2(n_44),
.B1(n_41),
.B2(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_51),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_79),
.Y(n_124)
);

AOI22x1_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_39),
.B1(n_44),
.B2(n_38),
.Y(n_79)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_85),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_44),
.B1(n_26),
.B2(n_18),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_88),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_62),
.B(n_67),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_19),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_19),
.CI(n_28),
.CON(n_93),
.SN(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_93),
.A2(n_9),
.B(n_15),
.C(n_14),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_49),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_61),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_68),
.B1(n_65),
.B2(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_109),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_63),
.A2(n_18),
.B1(n_41),
.B2(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_20),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_114),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_53),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_123),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_52),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_118),
.B(n_126),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_129),
.B1(n_138),
.B2(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_75),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_72),
.C(n_64),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_103),
.C(n_87),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_47),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_50),
.B1(n_64),
.B2(n_48),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_86),
.A2(n_48),
.B1(n_76),
.B2(n_21),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_139),
.B1(n_141),
.B2(n_104),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_48),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_137),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_21),
.B1(n_20),
.B2(n_2),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_79),
.A2(n_20),
.B1(n_9),
.B2(n_10),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_20),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_0),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_12),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_147),
.B(n_13),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_149),
.B1(n_154),
.B2(n_159),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_79),
.B1(n_78),
.B2(n_93),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_82),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_112),
.B(n_83),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_175),
.B(n_128),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_77),
.B1(n_80),
.B2(n_83),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_80),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_164),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_124),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_14),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_124),
.A2(n_111),
.B1(n_110),
.B2(n_90),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_179),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_119),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_99),
.B(n_94),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_99),
.C(n_94),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_126),
.C(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_118),
.A2(n_87),
.B1(n_90),
.B2(n_81),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g210 ( 
.A1(n_180),
.A2(n_191),
.B(n_194),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_195),
.C(n_145),
.Y(n_233)
);

OA21x2_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_144),
.B(n_129),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_119),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_202),
.Y(n_215)
);

AOI22x1_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_134),
.B1(n_147),
.B2(n_127),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_146),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_175),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_136),
.B(n_132),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_207),
.B(n_186),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_149),
.A2(n_132),
.B(n_120),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_0),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_165),
.A2(n_132),
.B(n_145),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_161),
.B(n_170),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_179),
.B1(n_154),
.B2(n_153),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_186),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_194),
.B1(n_182),
.B2(n_198),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_148),
.Y(n_213)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_177),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_183),
.C(n_195),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_171),
.B1(n_156),
.B2(n_151),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_193),
.B(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_164),
.Y(n_219)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_169),
.B(n_168),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_225),
.B(n_229),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_206),
.B1(n_208),
.B2(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_172),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_198),
.B(n_161),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_188),
.B(n_9),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_8),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_230),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_145),
.B(n_1),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_181),
.B(n_10),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_231),
.A2(n_190),
.B1(n_189),
.B2(n_199),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_185),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_220),
.B1(n_210),
.B2(n_218),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_5),
.C(n_14),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_239),
.C(n_242),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_191),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_252),
.B(n_221),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_191),
.B1(n_181),
.B2(n_196),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_220),
.B1(n_210),
.B2(n_218),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_204),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_222),
.C(n_215),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_244),
.C(n_254),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_203),
.C(n_196),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_190),
.B1(n_189),
.B2(n_203),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_228),
.B1(n_223),
.B2(n_213),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_232),
.C(n_228),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_211),
.B1(n_216),
.B2(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_269),
.Y(n_275)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_263),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_246),
.B1(n_263),
.B2(n_256),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_230),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_266),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_224),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_226),
.C(n_210),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_271),
.C(n_251),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_227),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_270),
.B(n_5),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_226),
.B1(n_199),
.B2(n_234),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_6),
.B(n_15),
.Y(n_270)
);

NOR3xp33_ASAP7_75t_SL g272 ( 
.A(n_270),
.B(n_251),
.C(n_239),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_277),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_12),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_242),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_281),
.B1(n_269),
.B2(n_262),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_238),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_260),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_249),
.B1(n_253),
.B2(n_247),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_257),
.A2(n_240),
.B1(n_252),
.B2(n_6),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_259),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_293),
.B1(n_276),
.B2(n_281),
.Y(n_295)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_288),
.B(n_292),
.Y(n_301)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_278),
.B1(n_277),
.B2(n_280),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_262),
.B(n_271),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_273),
.B(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_4),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_296),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_275),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_300),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_284),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_290),
.B1(n_294),
.B2(n_12),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_279),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_302),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_299),
.A3(n_301),
.B1(n_298),
.B2(n_302),
.C1(n_16),
.C2(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_297),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_310),
.A3(n_307),
.B1(n_306),
.B2(n_16),
.C1(n_294),
.C2(n_3),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_305),
.B(n_307),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_309),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_16),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_312),
.B1(n_1),
.B2(n_3),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_0),
.Y(n_315)
);


endmodule