module real_jpeg_32553_n_17 (n_8, n_0, n_141, n_2, n_139, n_142, n_143, n_10, n_137, n_9, n_12, n_147, n_146, n_6, n_11, n_14, n_138, n_7, n_3, n_145, n_144, n_5, n_4, n_1, n_140, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_141;
input n_2;
input n_139;
input n_142;
input n_143;
input n_10;
input n_137;
input n_9;
input n_12;
input n_147;
input n_146;
input n_6;
input n_11;
input n_14;
input n_138;
input n_7;
input n_3;
input n_145;
input n_144;
input n_5;
input n_4;
input n_1;
input n_140;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AND2x2_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_1),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_1),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g88 ( 
.A1(n_2),
.A2(n_9),
.B1(n_89),
.B2(n_93),
.C(n_95),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_3),
.A2(n_55),
.A3(n_57),
.B1(n_64),
.B2(n_127),
.C1(n_129),
.C2(n_147),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_5),
.B(n_118),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_7),
.B(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_9),
.B(n_89),
.C(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_13),
.B(n_40),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_14),
.B(n_73),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g123 ( 
.A(n_14),
.B(n_124),
.CON(n_123),
.SN(n_123)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_16),
.B(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_26),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_37),
.B(n_133),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_29),
.B(n_36),
.Y(n_134)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_45),
.B(n_132),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_42),
.B(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI31xp67_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_78),
.A3(n_116),
.B(n_121),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_63),
.C(n_72),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_48),
.A2(n_122),
.B(n_126),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_72),
.C(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_138),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OA21x2_ASAP7_75t_SL g122 ( 
.A1(n_63),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_109),
.C(n_110),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_99),
.B(n_108),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_88),
.B1(n_97),
.B2(n_98),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_143),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_107),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_137),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_139),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_140),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_141),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_142),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_144),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_145),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_146),
.Y(n_119)
);


endmodule