module real_aes_6674_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_1170;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1175;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_792;
wire n_673;
wire n_1067;
wire n_518;
wire n_635;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_1110;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_852;
wire n_1113;
wire n_766;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_1123;
wire n_549;
wire n_491;
wire n_694;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1166;
wire n_1137;
wire n_448;
wire n_556;
wire n_545;
wire n_752;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_638;
wire n_564;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_892;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_994;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_875;
wire n_467;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_1182;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_1180;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_1082;
wire n_468;
wire n_746;
wire n_1025;
wire n_532;
wire n_656;
wire n_755;
wire n_1168;
wire n_1148;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_725;
wire n_455;
wire n_504;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_1135;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_745;
wire n_722;
wire n_867;
wire n_1167;
wire n_1100;
wire n_1174;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_1112;
wire n_437;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_1041;
wire n_501;
wire n_1111;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_756;
wire n_1073;
wire n_404;
wire n_728;
wire n_713;
wire n_598;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_563;
wire n_785;
wire n_997;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1158;
wire n_1157;
wire n_1132;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_1056;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_1155;
wire n_1165;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_982;
wire n_717;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_1150;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_1143;
wire n_929;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_719;
wire n_566;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_1156;
wire n_1159;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_1176;
wire n_483;
wire n_611;
wire n_640;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1097;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_1101;
wire n_447;
wire n_1102;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_0), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_1), .A2(n_362), .B1(n_494), .B2(n_756), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g931 ( .A1(n_2), .A2(n_138), .B1(n_445), .B2(n_830), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_3), .A2(n_100), .B1(n_530), .B2(n_851), .Y(n_1013) );
AO22x2_ASAP7_75t_L g421 ( .A1(n_4), .A2(n_230), .B1(n_422), .B2(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g1124 ( .A(n_4), .Y(n_1124) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_5), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_6), .A2(n_156), .B1(n_517), .B2(n_578), .Y(n_825) );
AOI222xp33_ASAP7_75t_L g935 ( .A1(n_7), .A2(n_336), .B1(n_349), .B2(n_458), .C1(n_637), .C2(n_638), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_8), .Y(n_960) );
CKINVDCx20_ASAP7_75t_R g1149 ( .A(n_9), .Y(n_1149) );
INVx1_ASAP7_75t_L g818 ( .A(n_10), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_11), .A2(n_130), .B1(n_533), .B2(n_622), .Y(n_884) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_12), .A2(n_118), .B1(n_651), .B2(n_652), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_13), .A2(n_206), .B1(n_514), .B2(n_787), .C(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g802 ( .A(n_14), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_15), .A2(n_293), .B1(n_637), .B2(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g809 ( .A(n_16), .Y(n_809) );
INVx1_ASAP7_75t_L g1042 ( .A(n_17), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_18), .A2(n_328), .B1(n_576), .B2(n_581), .Y(n_1139) );
AOI22xp5_ASAP7_75t_SL g840 ( .A1(n_19), .A2(n_201), .B1(n_679), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_20), .A2(n_267), .B1(n_516), .B2(n_586), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g1016 ( .A1(n_21), .A2(n_216), .B1(n_585), .B2(n_586), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_22), .A2(n_159), .B1(n_673), .B2(n_781), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_23), .A2(n_110), .B1(n_513), .B2(n_684), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_24), .A2(n_331), .B1(n_888), .B2(n_1085), .Y(n_1084) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_25), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g1015 ( .A1(n_26), .A2(n_141), .B1(n_479), .B2(n_779), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_27), .A2(n_255), .B1(n_439), .B2(n_445), .Y(n_438) );
AO22x2_ASAP7_75t_L g425 ( .A1(n_28), .A2(n_117), .B1(n_422), .B2(n_426), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_29), .A2(n_81), .B1(n_439), .B2(n_610), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_30), .A2(n_277), .B1(n_517), .B2(n_574), .Y(n_751) );
AOI222xp33_ASAP7_75t_L g834 ( .A1(n_31), .A2(n_200), .B1(n_308), .B2(n_466), .C1(n_610), .C2(n_662), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_32), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_33), .A2(n_322), .B1(n_500), .B2(n_503), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_34), .B(n_1012), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_35), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_36), .A2(n_73), .B1(n_574), .B2(n_576), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_37), .A2(n_266), .B1(n_781), .B2(n_807), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_38), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g991 ( .A(n_39), .Y(n_991) );
CKINVDCx20_ASAP7_75t_R g1067 ( .A(n_40), .Y(n_1067) );
AOI22xp33_ASAP7_75t_SL g646 ( .A1(n_41), .A2(n_119), .B1(n_582), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_42), .A2(n_381), .B1(n_673), .B2(n_674), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_43), .A2(n_182), .B1(n_576), .B2(n_890), .Y(n_889) );
AOI22xp33_ASAP7_75t_SL g771 ( .A1(n_44), .A2(n_131), .B1(n_610), .B2(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_45), .B(n_556), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_46), .A2(n_76), .B1(n_488), .B2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_47), .A2(n_97), .B1(n_574), .B2(n_758), .Y(n_1106) );
CKINVDCx20_ASAP7_75t_R g1138 ( .A(n_48), .Y(n_1138) );
INVx1_ASAP7_75t_L g795 ( .A(n_49), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_50), .A2(n_146), .B1(n_513), .B2(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g618 ( .A(n_51), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_52), .A2(n_86), .B1(n_585), .B2(n_679), .Y(n_885) );
AOI22x1_ASAP7_75t_L g1047 ( .A1(n_53), .A2(n_1048), .B1(n_1073), .B2(n_1074), .Y(n_1047) );
CKINVDCx20_ASAP7_75t_R g1073 ( .A(n_53), .Y(n_1073) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_54), .A2(n_122), .B1(n_682), .B2(n_683), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_55), .A2(n_289), .B1(n_599), .B2(n_787), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_56), .Y(n_949) );
AO22x1_ASAP7_75t_L g971 ( .A1(n_57), .A2(n_972), .B1(n_999), .B2(n_1000), .Y(n_971) );
INVx1_ASAP7_75t_L g999 ( .A(n_57), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_58), .A2(n_95), .B1(n_484), .B2(n_927), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_59), .A2(n_321), .B1(n_473), .B2(n_625), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_60), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_61), .A2(n_193), .B1(n_439), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_62), .A2(n_179), .B1(n_585), .B2(n_993), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_63), .A2(n_305), .B1(n_812), .B2(n_906), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_64), .A2(n_83), .B1(n_523), .B2(n_1090), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_65), .A2(n_383), .B1(n_484), .B2(n_488), .Y(n_483) );
INVx1_ASAP7_75t_L g759 ( .A(n_66), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_67), .B(n_523), .Y(n_930) );
AOI22xp33_ASAP7_75t_SL g1018 ( .A1(n_68), .A2(n_396), .B1(n_844), .B2(n_890), .Y(n_1018) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_69), .A2(n_166), .B1(n_777), .B2(n_779), .Y(n_776) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_70), .A2(n_234), .B1(n_503), .B2(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_71), .A2(n_307), .B1(n_500), .B2(n_758), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_72), .A2(n_343), .B1(n_493), .B2(n_496), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_74), .A2(n_390), .B1(n_439), .B2(n_610), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_75), .Y(n_1032) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_77), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_78), .A2(n_209), .B1(n_493), .B2(n_888), .Y(n_887) );
CKINVDCx20_ASAP7_75t_R g945 ( .A(n_79), .Y(n_945) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_80), .A2(n_264), .B1(n_582), .B2(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_82), .A2(n_286), .B1(n_445), .B2(n_772), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_84), .A2(n_208), .B1(n_585), .B2(n_586), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_85), .A2(n_258), .B1(n_574), .B2(n_673), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_87), .A2(n_144), .B1(n_496), .B2(n_779), .Y(n_1174) );
AO22x2_ASAP7_75t_L g429 ( .A1(n_88), .A2(n_265), .B1(n_422), .B2(n_423), .Y(n_429) );
INVx1_ASAP7_75t_L g1121 ( .A(n_88), .Y(n_1121) );
CKINVDCx20_ASAP7_75t_R g1132 ( .A(n_89), .Y(n_1132) );
CKINVDCx20_ASAP7_75t_R g1051 ( .A(n_90), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_91), .A2(n_149), .B1(n_451), .B2(n_851), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_92), .A2(n_241), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_93), .A2(n_105), .B1(n_533), .B2(n_576), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_94), .A2(n_225), .B1(n_851), .B2(n_852), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g1064 ( .A(n_96), .Y(n_1064) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_98), .A2(n_279), .B1(n_441), .B2(n_538), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_99), .A2(n_195), .B1(n_522), .B2(n_526), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_101), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_102), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_103), .A2(n_387), .B1(n_627), .B2(n_830), .Y(n_829) );
AOI222xp33_ASAP7_75t_L g1108 ( .A1(n_104), .A2(n_112), .B1(n_185), .B2(n_550), .C1(n_638), .C2(n_644), .Y(n_1108) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_106), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_107), .A2(n_413), .B1(n_506), .B2(n_507), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_107), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_108), .A2(n_269), .B1(n_503), .B2(n_571), .Y(n_570) );
XOR2x2_ASAP7_75t_L g899 ( .A(n_109), .B(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g855 ( .A(n_111), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g1162 ( .A(n_113), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_114), .A2(n_285), .B1(n_647), .B2(n_675), .Y(n_933) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_115), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_116), .A2(n_274), .B1(n_498), .B2(n_756), .Y(n_839) );
INVx1_ASAP7_75t_L g1125 ( .A(n_117), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_120), .A2(n_268), .B1(n_845), .B2(n_1056), .Y(n_1055) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_121), .A2(n_311), .B1(n_844), .B2(n_845), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_123), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_124), .Y(n_1068) );
XOR2x2_ASAP7_75t_L g631 ( .A(n_125), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_126), .B(n_912), .Y(n_911) );
CKINVDCx20_ASAP7_75t_R g1166 ( .A(n_127), .Y(n_1166) );
CKINVDCx20_ASAP7_75t_R g975 ( .A(n_128), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_129), .A2(n_217), .B1(n_493), .B2(n_1171), .Y(n_1170) );
AO22x1_ASAP7_75t_L g1077 ( .A1(n_132), .A2(n_1078), .B1(n_1079), .B2(n_1093), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g1093 ( .A(n_132), .Y(n_1093) );
CKINVDCx20_ASAP7_75t_R g1063 ( .A(n_133), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_134), .A2(n_151), .B1(n_519), .B2(n_678), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g1161 ( .A(n_135), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_136), .B(n_910), .Y(n_909) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_137), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_139), .A2(n_363), .B1(n_475), .B2(n_494), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_140), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_142), .Y(n_1072) );
OAI22xp5_ASAP7_75t_SL g864 ( .A1(n_143), .A2(n_865), .B1(n_866), .B2(n_892), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_143), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_145), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_147), .A2(n_360), .B1(n_516), .B2(n_518), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_148), .A2(n_163), .B1(n_484), .B2(n_679), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_150), .A2(n_373), .B1(n_686), .B2(n_787), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_152), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g1145 ( .A(n_153), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_154), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_155), .A2(n_207), .B1(n_538), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_157), .A2(n_313), .B1(n_533), .B2(n_684), .Y(n_925) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_158), .A2(n_355), .B1(n_686), .B2(n_688), .Y(n_685) );
AND2x6_ASAP7_75t_L g401 ( .A(n_160), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_160), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_161), .A2(n_292), .B1(n_518), .B2(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_162), .A2(n_344), .B1(n_466), .B2(n_627), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_164), .A2(n_270), .B1(n_556), .B2(n_815), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g1152 ( .A(n_165), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_167), .A2(n_348), .B1(n_679), .B2(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_168), .A2(n_334), .B1(n_488), .B2(n_601), .Y(n_721) );
AOI222xp33_ASAP7_75t_L g626 ( .A1(n_169), .A2(n_244), .B1(n_263), .B2(n_460), .C1(n_556), .C2(n_627), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g936 ( .A(n_170), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_171), .A2(n_320), .B1(n_513), .B2(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g628 ( .A(n_172), .Y(n_628) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_173), .A2(n_351), .B1(n_804), .B2(n_847), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g1058 ( .A(n_174), .Y(n_1058) );
INVx1_ASAP7_75t_L g998 ( .A(n_175), .Y(n_998) );
INVx1_ASAP7_75t_L g817 ( .A(n_176), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_177), .A2(n_326), .B1(n_514), .B2(n_847), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_178), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_180), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_181), .A2(n_399), .B(n_407), .C(n_1126), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_183), .A2(n_259), .B1(n_585), .B2(n_586), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_184), .A2(n_251), .B1(n_536), .B2(n_601), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_186), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_187), .A2(n_365), .B1(n_675), .B2(n_1041), .Y(n_1040) );
AO22x2_ASAP7_75t_L g431 ( .A1(n_188), .A2(n_252), .B1(n_422), .B2(n_426), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g1122 ( .A(n_188), .B(n_1123), .Y(n_1122) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_189), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_190), .A2(n_223), .B1(n_518), .B2(n_921), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g929 ( .A(n_191), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_192), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_194), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_196), .A2(n_385), .B1(n_535), .B2(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g1007 ( .A(n_197), .Y(n_1007) );
XOR2xp5_ASAP7_75t_L g1127 ( .A(n_198), .B(n_1128), .Y(n_1127) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_199), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g1092 ( .A1(n_202), .A2(n_342), .B1(n_350), .B2(n_465), .C1(n_538), .C2(n_550), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_203), .A2(n_257), .B1(n_501), .B2(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_204), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_205), .A2(n_357), .B1(n_677), .B2(n_679), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_210), .A2(n_283), .B1(n_608), .B2(n_670), .Y(n_669) );
XOR2x2_ASAP7_75t_L g1095 ( .A(n_211), .B(n_1096), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_212), .A2(n_317), .B1(n_526), .B2(n_745), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_213), .Y(n_835) );
OA22x2_ASAP7_75t_L g791 ( .A1(n_214), .A2(n_792), .B1(n_793), .B2(n_820), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_214), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g994 ( .A1(n_215), .A2(n_303), .B1(n_513), .B2(n_571), .C(n_995), .Y(n_994) );
INVx1_ASAP7_75t_L g620 ( .A(n_218), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_219), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_220), .A2(n_312), .B1(n_745), .B2(n_747), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_221), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_222), .B(n_665), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_224), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_226), .A2(n_273), .B1(n_494), .B2(n_678), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_227), .B(n_526), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_228), .A2(n_302), .B1(n_582), .B2(n_1103), .Y(n_1102) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_229), .A2(n_249), .B1(n_530), .B2(n_666), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_231), .A2(n_325), .B1(n_445), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_232), .A2(n_291), .B1(n_479), .B2(n_753), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_233), .A2(n_304), .B1(n_439), .B2(n_644), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_235), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g1101 ( .A1(n_236), .A2(n_384), .B1(n_519), .B2(n_756), .Y(n_1101) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_237), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_238), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_239), .Y(n_965) );
INVx1_ASAP7_75t_L g613 ( .A(n_240), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_242), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_243), .A2(n_347), .B1(n_627), .B2(n_830), .Y(n_1099) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_245), .A2(n_364), .B1(n_376), .B2(n_460), .C1(n_465), .C2(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_246), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_247), .A2(n_395), .B1(n_522), .B2(n_670), .Y(n_773) );
AND2x2_ASAP7_75t_L g405 ( .A(n_248), .B(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_250), .A2(n_287), .B1(n_666), .B2(n_906), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_253), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g1134 ( .A(n_254), .Y(n_1134) );
XNOR2xp5_ASAP7_75t_L g760 ( .A(n_256), .B(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_260), .A2(n_309), .B1(n_466), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_261), .A2(n_380), .B1(n_571), .B2(n_581), .Y(n_1081) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_262), .Y(n_551) );
INVx1_ASAP7_75t_L g1033 ( .A(n_271), .Y(n_1033) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_272), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_275), .A2(n_300), .B1(n_682), .B2(n_847), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_276), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_278), .A2(n_540), .B1(n_587), .B2(n_588), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_278), .Y(n_587) );
INVx1_ASAP7_75t_L g796 ( .A(n_280), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_281), .A2(n_393), .B1(n_578), .B2(n_654), .Y(n_653) );
XOR2x2_ASAP7_75t_L g1003 ( .A(n_282), .B(n_1004), .Y(n_1003) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_284), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_288), .A2(n_345), .B1(n_688), .B2(n_725), .Y(n_1175) );
INVx1_ASAP7_75t_L g422 ( .A(n_290), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_290), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_294), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_295), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_296), .A2(n_382), .B1(n_585), .B2(n_586), .Y(n_1135) );
AOI22xp5_ASAP7_75t_L g1157 ( .A1(n_297), .A2(n_1158), .B1(n_1176), .B2(n_1177), .Y(n_1157) );
CKINVDCx20_ASAP7_75t_R g1176 ( .A(n_297), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_298), .A2(n_353), .B1(n_652), .B2(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_299), .B(n_523), .Y(n_642) );
INVx1_ASAP7_75t_L g819 ( .A(n_301), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_306), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_310), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g1142 ( .A(n_314), .Y(n_1142) );
INVx1_ASAP7_75t_L g810 ( .A(n_315), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g1165 ( .A(n_316), .Y(n_1165) );
INVx1_ASAP7_75t_L g996 ( .A(n_318), .Y(n_996) );
OA22x2_ASAP7_75t_L g656 ( .A1(n_319), .A2(n_657), .B1(n_658), .B2(n_690), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_319), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_323), .A2(n_391), .B1(n_523), .B2(n_528), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_324), .A2(n_366), .B1(n_689), .B2(n_725), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_327), .Y(n_720) );
INVx1_ASAP7_75t_L g406 ( .A(n_329), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g1137 ( .A(n_330), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_332), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g402 ( .A(n_333), .Y(n_402) );
INVx1_ASAP7_75t_L g858 ( .A(n_335), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g1071 ( .A(n_337), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g904 ( .A(n_338), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_339), .A2(n_346), .B1(n_503), .B2(n_756), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_340), .Y(n_1029) );
INVx1_ASAP7_75t_L g623 ( .A(n_341), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_352), .A2(n_375), .B1(n_601), .B2(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g976 ( .A(n_354), .Y(n_976) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_356), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g1059 ( .A(n_358), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_359), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_361), .Y(n_558) );
INVx1_ASAP7_75t_L g604 ( .A(n_367), .Y(n_604) );
CKINVDCx20_ASAP7_75t_R g1151 ( .A(n_368), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_369), .B(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_370), .B(n_465), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_371), .B(n_526), .Y(n_641) );
XOR2x2_ASAP7_75t_L g509 ( .A(n_372), .B(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_374), .A2(n_698), .B1(n_727), .B2(n_728), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_374), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g1146 ( .A(n_377), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_378), .B(n_607), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_379), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_386), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_388), .Y(n_988) );
CKINVDCx20_ASAP7_75t_R g1167 ( .A(n_389), .Y(n_1167) );
INVx1_ASAP7_75t_L g805 ( .A(n_392), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_394), .A2(n_940), .B1(n_966), .B2(n_967), .Y(n_939) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_394), .Y(n_966) );
CKINVDCx20_ASAP7_75t_R g1027 ( .A(n_397), .Y(n_1027) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_402), .Y(n_1117) );
OAI21xp5_ASAP7_75t_L g1182 ( .A1(n_403), .A2(n_1116), .B(n_1183), .Y(n_1182) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_861), .B1(n_1111), .B2(n_1112), .C(n_1113), .Y(n_407) );
INVx1_ASAP7_75t_L g1112 ( .A(n_408), .Y(n_1112) );
XNOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_732), .Y(n_408) );
XNOR2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_593), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_508), .B1(n_591), .B2(n_592), .Y(n_410) );
INVx1_ASAP7_75t_L g591 ( .A(n_411), .Y(n_591) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g507 ( .A(n_413), .Y(n_507) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_470), .Y(n_413) );
NOR2xp33_ASAP7_75t_SL g414 ( .A(n_415), .B(n_449), .Y(n_414) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_432), .B1(n_433), .B2(n_437), .C(n_438), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_416), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g808 ( .A1(n_416), .A2(n_433), .B1(n_809), .B2(n_810), .C(n_811), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_416), .A2(n_1063), .B1(n_1064), .B2(n_1065), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_416), .A2(n_1065), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
OAI221xp5_ASAP7_75t_L g1160 ( .A1(n_416), .A2(n_545), .B1(n_1161), .B2(n_1162), .C(n_1163), .Y(n_1160) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g870 ( .A(n_417), .Y(n_870) );
INVx2_ASAP7_75t_L g957 ( .A(n_417), .Y(n_957) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_418), .Y(n_702) );
BUFx3_ASAP7_75t_L g1026 ( .A(n_418), .Y(n_1026) );
OR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_427), .Y(n_418) );
INVx2_ASAP7_75t_L g476 ( .A(n_419), .Y(n_476) );
OR2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_425), .Y(n_419) );
AND2x2_ASAP7_75t_L g436 ( .A(n_420), .B(n_425), .Y(n_436) );
AND2x2_ASAP7_75t_L g481 ( .A(n_420), .B(n_455), .Y(n_481) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g444 ( .A(n_421), .B(n_431), .Y(n_444) );
AND2x2_ASAP7_75t_L g448 ( .A(n_421), .B(n_425), .Y(n_448) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_424), .Y(n_426) );
INVx1_ASAP7_75t_L g443 ( .A(n_425), .Y(n_443) );
INVx2_ASAP7_75t_L g455 ( .A(n_425), .Y(n_455) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_428), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g480 ( .A(n_428), .B(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g525 ( .A(n_428), .B(n_476), .Y(n_525) );
AND2x6_ASAP7_75t_L g528 ( .A(n_428), .B(n_436), .Y(n_528) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g447 ( .A(n_429), .Y(n_447) );
INVx1_ASAP7_75t_L g454 ( .A(n_429), .Y(n_454) );
INVx1_ASAP7_75t_L g462 ( .A(n_429), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_429), .B(n_431), .Y(n_490) );
AND2x2_ASAP7_75t_L g461 ( .A(n_430), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g487 ( .A(n_431), .B(n_447), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_433), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_433), .A2(n_1025), .B1(n_1026), .B2(n_1027), .Y(n_1024) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g977 ( .A(n_434), .Y(n_977) );
INVx2_ASAP7_75t_L g1065 ( .A(n_434), .Y(n_1065) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g547 ( .A(n_435), .Y(n_547) );
AND2x2_ASAP7_75t_L g486 ( .A(n_436), .B(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_L g498 ( .A(n_436), .B(n_461), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g990 ( .A(n_436), .B(n_487), .Y(n_990) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g812 ( .A(n_440), .Y(n_812) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g772 ( .A(n_441), .Y(n_772) );
BUFx3_ASAP7_75t_L g830 ( .A(n_441), .Y(n_830) );
BUFx2_ASAP7_75t_L g851 ( .A(n_441), .Y(n_851) );
AND2x4_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x6_ASAP7_75t_L g489 ( .A(n_443), .B(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g452 ( .A(n_444), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g467 ( .A(n_444), .B(n_468), .Y(n_467) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_444), .B(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_SL g530 ( .A(n_445), .Y(n_530) );
BUFx3_ASAP7_75t_L g610 ( .A(n_445), .Y(n_610) );
BUFx2_ASAP7_75t_SL g644 ( .A(n_445), .Y(n_644) );
BUFx6f_ASAP7_75t_L g852 ( .A(n_445), .Y(n_852) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g567 ( .A(n_446), .Y(n_567) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x6_ASAP7_75t_L g460 ( .A(n_448), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g566 ( .A(n_448), .Y(n_566) );
OAI222xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_456), .B1(n_457), .B2(n_463), .C1(n_464), .C2(n_469), .Y(n_449) );
OAI222xp33_ASAP7_75t_L g1164 ( .A1(n_450), .A2(n_740), .B1(n_1147), .B2(n_1165), .C1(n_1166), .C2(n_1167), .Y(n_1164) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx4f_ASAP7_75t_SL g538 ( .A(n_452), .Y(n_538) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_452), .Y(n_627) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_452), .Y(n_766) );
BUFx2_ASAP7_75t_L g857 ( .A(n_452), .Y(n_857) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g468 ( .A(n_454), .Y(n_468) );
INVx1_ASAP7_75t_L g561 ( .A(n_455), .Y(n_561) );
OAI221xp5_ASAP7_75t_SL g872 ( .A1(n_457), .A2(n_873), .B1(n_874), .B2(n_875), .C(n_876), .Y(n_872) );
OAI21xp5_ASAP7_75t_SL g1006 ( .A1(n_457), .A2(n_1007), .B(n_1008), .Y(n_1006) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx4_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI222xp33_ASAP7_75t_L g813 ( .A1(n_459), .A2(n_464), .B1(n_814), .B2(n_817), .C1(n_818), .C2(n_819), .Y(n_813) );
BUFx2_ASAP7_75t_L g854 ( .A(n_459), .Y(n_854) );
INVx4_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_460), .Y(n_550) );
BUFx3_ASAP7_75t_L g662 ( .A(n_460), .Y(n_662) );
INVx2_ASAP7_75t_L g740 ( .A(n_460), .Y(n_740) );
INVx2_ASAP7_75t_SL g903 ( .A(n_460), .Y(n_903) );
AND2x6_ASAP7_75t_L g475 ( .A(n_461), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g495 ( .A(n_461), .B(n_481), .Y(n_495) );
OAI222xp33_ASAP7_75t_L g1066 ( .A1(n_464), .A2(n_552), .B1(n_707), .B2(n_1067), .C1(n_1068), .C2(n_1069), .Y(n_1066) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx4f_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g639 ( .A(n_466), .Y(n_639) );
BUFx12f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_467), .Y(n_666) );
INVx1_ASAP7_75t_L g768 ( .A(n_467), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_491), .Y(n_470) );
OAI221xp5_ASAP7_75t_SL g471 ( .A1(n_472), .A2(n_477), .B1(n_478), .B2(n_482), .C(n_483), .Y(n_471) );
OAI221xp5_ASAP7_75t_SL g1136 ( .A1(n_472), .A2(n_1052), .B1(n_1137), .B2(n_1138), .C(n_1139), .Y(n_1136) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g535 ( .A(n_474), .Y(n_535) );
INVx2_ASAP7_75t_SL g781 ( .A(n_474), .Y(n_781) );
INVx2_ASAP7_75t_L g845 ( .A(n_474), .Y(n_845) );
HB1xp67_ASAP7_75t_L g1086 ( .A(n_474), .Y(n_1086) );
INVx11_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx11_ASAP7_75t_L g575 ( .A(n_475), .Y(n_575) );
INVx4_ASAP7_75t_L g514 ( .A(n_478), .Y(n_514) );
INVx3_ASAP7_75t_L g599 ( .A(n_478), .Y(n_599) );
OAI221xp5_ASAP7_75t_SL g717 ( .A1(n_478), .A2(n_718), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_717) );
OAI221xp5_ASAP7_75t_SL g794 ( .A1(n_478), .A2(n_778), .B1(n_795), .B2(n_796), .C(n_797), .Y(n_794) );
INVx4_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g583 ( .A(n_480), .Y(n_583) );
BUFx3_ASAP7_75t_L g675 ( .A(n_480), .Y(n_675) );
BUFx3_ASAP7_75t_L g888 ( .A(n_480), .Y(n_888) );
BUFx3_ASAP7_75t_L g921 ( .A(n_480), .Y(n_921) );
AND2x2_ASAP7_75t_L g502 ( .A(n_481), .B(n_487), .Y(n_502) );
AND2x4_ASAP7_75t_L g504 ( .A(n_481), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_481), .B(n_487), .Y(n_616) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx5_ASAP7_75t_L g517 ( .A(n_485), .Y(n_517) );
BUFx3_ASAP7_75t_L g602 ( .A(n_485), .Y(n_602) );
INVx2_ASAP7_75t_L g678 ( .A(n_485), .Y(n_678) );
INVx4_ASAP7_75t_L g800 ( .A(n_485), .Y(n_800) );
INVx1_ASAP7_75t_L g953 ( .A(n_485), .Y(n_953) );
INVx8_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx6_ASAP7_75t_SL g519 ( .A(n_489), .Y(n_519) );
INVx1_ASAP7_75t_SL g783 ( .A(n_489), .Y(n_783) );
INVx1_ASAP7_75t_L g505 ( .A(n_490), .Y(n_505) );
NAND2xp33_ASAP7_75t_SL g491 ( .A(n_492), .B(n_499), .Y(n_491) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx3_ASAP7_75t_L g581 ( .A(n_494), .Y(n_581) );
INVx3_ASAP7_75t_L g778 ( .A(n_494), .Y(n_778) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_494), .Y(n_844) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_SL g513 ( .A(n_495), .Y(n_513) );
BUFx2_ASAP7_75t_SL g647 ( .A(n_495), .Y(n_647) );
INVx2_ASAP7_75t_L g687 ( .A(n_495), .Y(n_687) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g536 ( .A(n_497), .Y(n_536) );
INVx3_ASAP7_75t_L g625 ( .A(n_497), .Y(n_625) );
INVx2_ASAP7_75t_L g804 ( .A(n_497), .Y(n_804) );
INVx6_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx3_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
BUFx3_ASAP7_75t_L g673 ( .A(n_498), .Y(n_673) );
BUFx3_ASAP7_75t_L g758 ( .A(n_498), .Y(n_758) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g572 ( .A(n_501), .Y(n_572) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx3_ASAP7_75t_L g651 ( .A(n_502), .Y(n_651) );
BUFx3_ASAP7_75t_L g684 ( .A(n_502), .Y(n_684) );
BUFx3_ASAP7_75t_L g756 ( .A(n_502), .Y(n_756) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_503), .Y(n_1056) );
INVx2_ASAP7_75t_L g1133 ( .A(n_503), .Y(n_1133) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx3_ASAP7_75t_L g533 ( .A(n_504), .Y(n_533) );
BUFx2_ASAP7_75t_SL g652 ( .A(n_504), .Y(n_652) );
BUFx3_ASAP7_75t_L g689 ( .A(n_504), .Y(n_689) );
BUFx3_ASAP7_75t_L g787 ( .A(n_504), .Y(n_787) );
BUFx2_ASAP7_75t_SL g847 ( .A(n_504), .Y(n_847) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_504), .Y(n_1041) );
INVx1_ASAP7_75t_L g1104 ( .A(n_504), .Y(n_1104) );
AND2x2_ASAP7_75t_L g753 ( .A(n_505), .B(n_561), .Y(n_753) );
INVx3_ASAP7_75t_L g592 ( .A(n_508), .Y(n_592) );
OA22x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_539), .B1(n_589), .B2(n_590), .Y(n_508) );
INVx1_ASAP7_75t_L g590 ( .A(n_509), .Y(n_590) );
XNOR2xp5_ASAP7_75t_L g696 ( .A(n_509), .B(n_631), .Y(n_696) );
NAND4xp75_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .C(n_531), .D(n_537), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g718 ( .A(n_513), .Y(n_718) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g585 ( .A(n_517), .Y(n_585) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g586 ( .A(n_519), .Y(n_586) );
BUFx2_ASAP7_75t_L g679 ( .A(n_519), .Y(n_679) );
BUFx2_ASAP7_75t_L g927 ( .A(n_519), .Y(n_927) );
BUFx4f_ASAP7_75t_SL g993 ( .A(n_519), .Y(n_993) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_521), .B(n_529), .Y(n_520) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_523), .Y(n_910) );
INVx5_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g608 ( .A(n_524), .Y(n_608) );
INVx2_ASAP7_75t_L g745 ( .A(n_524), .Y(n_745) );
INVx2_ASAP7_75t_L g1012 ( .A(n_524), .Y(n_1012) );
INVx4_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_SL g670 ( .A(n_527), .Y(n_670) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
BUFx4f_ASAP7_75t_L g747 ( .A(n_528), .Y(n_747) );
BUFx2_ASAP7_75t_L g912 ( .A(n_528), .Y(n_912) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_528), .Y(n_1090) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
INVxp67_ASAP7_75t_L g617 ( .A(n_533), .Y(n_617) );
INVx1_ASAP7_75t_L g552 ( .A(n_538), .Y(n_552) );
INVx1_ASAP7_75t_L g705 ( .A(n_538), .Y(n_705) );
INVx1_ASAP7_75t_L g589 ( .A(n_539), .Y(n_589) );
INVx2_ASAP7_75t_L g588 ( .A(n_540), .Y(n_588) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_568), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .C(n_557), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_545), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_545), .A2(n_869), .B1(n_870), .B2(n_871), .Y(n_868) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g605 ( .A(n_547), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_551), .B1(n_552), .B2(n_553), .C(n_554), .Y(n_548) );
OAI21xp5_ASAP7_75t_SL g634 ( .A1(n_549), .A2(n_635), .B(n_636), .Y(n_634) );
OAI222xp33_ASAP7_75t_L g763 ( .A1(n_549), .A2(n_764), .B1(n_765), .B2(n_767), .C1(n_768), .C2(n_769), .Y(n_763) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g707 ( .A(n_550), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g959 ( .A1(n_552), .A2(n_903), .B1(n_960), .B2(n_961), .C(n_962), .Y(n_959) );
BUFx4f_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_562), .B2(n_563), .Y(n_557) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx4_ASAP7_75t_L g714 ( .A(n_560), .Y(n_714) );
BUFx3_ASAP7_75t_L g879 ( .A(n_560), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_563), .A2(n_712), .B1(n_713), .B2(n_715), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_563), .A2(n_713), .B1(n_964), .B2(n_965), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_563), .A2(n_713), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_563), .A2(n_713), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g881 ( .A(n_564), .Y(n_881) );
CKINVDCx16_ASAP7_75t_R g564 ( .A(n_565), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_565), .A2(n_879), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
OR2x6_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_579), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx4_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx3_ASAP7_75t_L g622 ( .A(n_575), .Y(n_622) );
INVx2_ASAP7_75t_SL g654 ( .A(n_575), .Y(n_654) );
INVx4_ASAP7_75t_L g682 ( .A(n_575), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g801 ( .A1(n_575), .A2(n_802), .B1(n_803), .B2(n_805), .C(n_806), .Y(n_801) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_584), .Y(n_579) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g1171 ( .A(n_583), .Y(n_1171) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_693), .B1(n_730), .B2(n_731), .Y(n_593) );
INVx1_ASAP7_75t_L g730 ( .A(n_594), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_629), .B1(n_630), .B2(n_692), .Y(n_594) );
INVx2_ASAP7_75t_L g692 ( .A(n_595), .Y(n_692) );
XOR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_628), .Y(n_595) );
NAND4xp75_ASAP7_75t_L g596 ( .A(n_597), .B(n_603), .C(n_611), .D(n_626), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OA211x2_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B(n_606), .C(n_609), .Y(n_603) );
OA211x2_ASAP7_75t_L g928 ( .A1(n_605), .A2(n_929), .B(n_930), .C(n_931), .Y(n_928) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_619), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_617), .B2(n_618), .Y(n_612) );
OAI221xp5_ASAP7_75t_SL g947 ( .A1(n_614), .A2(n_948), .B1(n_949), .B2(n_950), .C(n_951), .Y(n_947) );
OAI221xp5_ASAP7_75t_SL g1057 ( .A1(n_614), .A2(n_803), .B1(n_1058), .B2(n_1059), .C(n_1060), .Y(n_1057) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g1131 ( .A(n_615), .Y(n_1131) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_623), .B2(n_624), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_627), .Y(n_637) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_655), .B1(n_656), .B2(n_691), .Y(n_630) );
INVx1_ASAP7_75t_L g691 ( .A(n_631), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_645), .C(n_649), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_640), .Y(n_633) );
INVx2_ASAP7_75t_SL g874 ( .A(n_637), .Y(n_874) );
INVx2_ASAP7_75t_SL g980 ( .A(n_637), .Y(n_980) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .C(n_643), .Y(n_640) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
INVx1_ASAP7_75t_L g726 ( .A(n_651), .Y(n_726) );
BUFx4f_ASAP7_75t_SL g807 ( .A(n_651), .Y(n_807) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g690 ( .A(n_658), .Y(n_690) );
NAND3x1_ASAP7_75t_L g658 ( .A(n_659), .B(n_671), .C(n_680), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_667), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_663), .B(n_664), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g978 ( .A1(n_661), .A2(n_979), .B1(n_980), .B2(n_981), .C(n_982), .Y(n_978) );
OAI21xp33_ASAP7_75t_L g1028 ( .A1(n_661), .A2(n_1029), .B(n_1030), .Y(n_1028) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g709 ( .A(n_666), .Y(n_709) );
BUFx3_ASAP7_75t_L g1148 ( .A(n_666), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_676), .Y(n_671) );
INVx1_ASAP7_75t_L g948 ( .A(n_673), .Y(n_948) );
INVx1_ASAP7_75t_L g944 ( .A(n_674), .Y(n_944) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_685), .Y(n_680) );
INVx1_ASAP7_75t_L g997 ( .A(n_682), .Y(n_997) );
BUFx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g731 ( .A(n_693), .Y(n_731) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_729), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g729 ( .A(n_697), .Y(n_729) );
INVx1_ASAP7_75t_L g728 ( .A(n_698), .Y(n_728) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_716), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_704), .C(n_711), .Y(n_699) );
OAI222xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_708), .C1(n_709), .C2(n_710), .Y(n_704) );
OAI222xp33_ASAP7_75t_L g1144 ( .A1(n_707), .A2(n_874), .B1(n_1145), .B2(n_1146), .C1(n_1147), .C2(n_1149), .Y(n_1144) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_713), .A2(n_881), .B1(n_984), .B2(n_985), .Y(n_983) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_722), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_789), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OA22x2_ASAP7_75t_SL g734 ( .A1(n_735), .A2(n_736), .B1(n_760), .B2(n_788), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
XOR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_759), .Y(n_736) );
NAND2x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_749), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
OAI21xp5_ASAP7_75t_SL g739 ( .A1(n_740), .A2(n_741), .B(n_742), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .C(n_748), .Y(n_743) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_754), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
INVx1_ASAP7_75t_L g891 ( .A(n_756), .Y(n_891) );
INVx1_ASAP7_75t_L g788 ( .A(n_760), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_774), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_770), .Y(n_762) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx4_ASAP7_75t_L g816 ( .A(n_766), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_784), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_782), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI221xp5_ASAP7_75t_SL g942 ( .A1(n_778), .A2(n_943), .B1(n_944), .B2(n_945), .C(n_946), .Y(n_942) );
OAI221xp5_ASAP7_75t_SL g1050 ( .A1(n_778), .A2(n_1051), .B1(n_1052), .B2(n_1054), .C(n_1055), .Y(n_1050) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_821), .B1(n_859), .B2(n_860), .Y(n_790) );
INVx1_ASAP7_75t_L g859 ( .A(n_791), .Y(n_859) );
INVx1_ASAP7_75t_L g820 ( .A(n_793), .Y(n_820) );
OR4x1_ASAP7_75t_L g793 ( .A(n_794), .B(n_801), .C(n_808), .D(n_813), .Y(n_793) );
INVx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
BUFx6f_ASAP7_75t_L g841 ( .A(n_800), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_803), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_995) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx3_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g860 ( .A(n_821), .Y(n_860) );
XNOR2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_836), .Y(n_821) );
XOR2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_835), .Y(n_822) );
NAND4xp75_ASAP7_75t_L g823 ( .A(n_824), .B(n_827), .C(n_831), .D(n_834), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
AND2x2_ASAP7_75t_SL g827 ( .A(n_828), .B(n_829), .Y(n_827) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
XOR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_858), .Y(n_836) );
NOR4xp75_ASAP7_75t_L g837 ( .A(n_838), .B(n_842), .C(n_848), .D(n_853), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g838 ( .A(n_839), .B(n_840), .Y(n_838) );
NAND2x1_ASAP7_75t_L g842 ( .A(n_843), .B(n_846), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx1_ASAP7_75t_SL g907 ( .A(n_852), .Y(n_907) );
OAI21xp5_ASAP7_75t_SL g853 ( .A1(n_854), .A2(n_855), .B(n_856), .Y(n_853) );
INVx1_ASAP7_75t_L g1111 ( .A(n_861), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_893), .B2(n_1110), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
BUFx2_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_SL g865 ( .A(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_882), .Y(n_866) );
NOR3xp33_ASAP7_75t_L g867 ( .A(n_868), .B(n_872), .C(n_877), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_870), .A2(n_975), .B1(n_976), .B2(n_977), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B1(n_880), .B2(n_881), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_886), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_889), .Y(n_886) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g1110 ( .A(n_893), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_895), .B1(n_1044), .B2(n_1045), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_897), .B1(n_968), .B2(n_969), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
XNOR2xp5_ASAP7_75t_L g897 ( .A(n_898), .B(n_939), .Y(n_897) );
AO22x2_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_922), .B1(n_937), .B2(n_938), .Y(n_898) );
INVx2_ASAP7_75t_L g937 ( .A(n_899), .Y(n_937) );
XOR2x2_ASAP7_75t_L g1094 ( .A(n_899), .B(n_1095), .Y(n_1094) );
NAND2xp5_ASAP7_75t_SL g900 ( .A(n_901), .B(n_914), .Y(n_900) );
NOR2xp33_ASAP7_75t_SL g901 ( .A(n_902), .B(n_908), .Y(n_901) );
OAI21xp5_ASAP7_75t_SL g902 ( .A1(n_903), .A2(n_904), .B(n_905), .Y(n_902) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
NAND3xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_911), .C(n_913), .Y(n_908) );
NOR2x1_ASAP7_75t_L g914 ( .A(n_915), .B(n_918), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_921), .Y(n_1053) );
INVx3_ASAP7_75t_SL g938 ( .A(n_922), .Y(n_938) );
XOR2x2_ASAP7_75t_L g922 ( .A(n_923), .B(n_936), .Y(n_922) );
NAND4xp75_ASAP7_75t_L g923 ( .A(n_924), .B(n_928), .C(n_932), .D(n_935), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_925), .B(n_926), .Y(n_924) );
AND2x2_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .Y(n_932) );
INVx2_ASAP7_75t_L g967 ( .A(n_940), .Y(n_967) );
AND2x2_ASAP7_75t_SL g940 ( .A(n_941), .B(n_954), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_942), .B(n_947), .Y(n_941) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
NOR3xp33_ASAP7_75t_L g954 ( .A(n_955), .B(n_959), .C(n_963), .Y(n_954) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g969 ( .A1(n_970), .A2(n_971), .B1(n_1001), .B2(n_1002), .Y(n_969) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g1000 ( .A(n_972), .Y(n_1000) );
AND3x1_ASAP7_75t_L g972 ( .A(n_973), .B(n_986), .C(n_994), .Y(n_972) );
NOR3xp33_ASAP7_75t_L g973 ( .A(n_974), .B(n_978), .C(n_983), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_989), .B1(n_991), .B2(n_992), .Y(n_987) );
BUFx2_ASAP7_75t_R g989 ( .A(n_990), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g992 ( .A(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_1003), .A2(n_1020), .B1(n_1021), .B2(n_1043), .Y(n_1002) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1003), .Y(n_1043) );
NAND3x2_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1014), .C(n_1017), .Y(n_1004) );
NOR2x1_ASAP7_75t_SL g1005 ( .A(n_1006), .B(n_1009), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .C(n_1013), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_1021), .Y(n_1020) );
XOR2x2_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1042), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1034), .Y(n_1022) );
NOR3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1028), .C(n_1031), .Y(n_1023) );
NOR2xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1038), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1045 ( .A1(n_1046), .A2(n_1047), .B1(n_1075), .B2(n_1109), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1048), .Y(n_1074) );
AND2x2_ASAP7_75t_SL g1048 ( .A(n_1049), .B(n_1061), .Y(n_1048) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1057), .Y(n_1049) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
NOR3xp33_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1066), .C(n_1070), .Y(n_1061) );
INVx2_ASAP7_75t_L g1109 ( .A(n_1075), .Y(n_1109) );
XNOR2x1_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1094), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_SL g1078 ( .A(n_1079), .Y(n_1078) );
NAND4xp75_ASAP7_75t_SL g1079 ( .A(n_1080), .B(n_1083), .C(n_1088), .D(n_1092), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1087), .Y(n_1083) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
AND2x2_ASAP7_75t_SL g1088 ( .A(n_1089), .B(n_1091), .Y(n_1088) );
NAND4xp75_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1100), .C(n_1105), .D(n_1108), .Y(n_1096) );
AND2x2_ASAP7_75t_SL g1097 ( .A(n_1098), .B(n_1099), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1102), .Y(n_1100) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1107), .Y(n_1105) );
INVx1_ASAP7_75t_SL g1113 ( .A(n_1114), .Y(n_1113) );
NOR2x1_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1119), .Y(n_1114) );
OR2x2_ASAP7_75t_SL g1180 ( .A(n_1115), .B(n_1120), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1118), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1116), .B(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1117), .B(n_1154), .Y(n_1183) );
CKINVDCx16_ASAP7_75t_R g1154 ( .A(n_1118), .Y(n_1154) );
CKINVDCx20_ASAP7_75t_R g1119 ( .A(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1122), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1125), .Y(n_1123) );
OAI222xp33_ASAP7_75t_L g1126 ( .A1(n_1127), .A2(n_1153), .B1(n_1155), .B2(n_1176), .C1(n_1178), .C2(n_1181), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1140), .Y(n_1128) );
NOR2xp33_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1136), .Y(n_1129) );
OAI221xp5_ASAP7_75t_SL g1130 ( .A1(n_1131), .A2(n_1132), .B1(n_1133), .B2(n_1134), .C(n_1135), .Y(n_1130) );
NOR3xp33_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1144), .C(n_1150), .Y(n_1140) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_SL g1177 ( .A(n_1158), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1159), .B(n_1168), .Y(n_1158) );
NOR2xp33_ASAP7_75t_SL g1159 ( .A(n_1160), .B(n_1164), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1173), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1172), .Y(n_1169) );
NAND2xp5_ASAP7_75t_SL g1173 ( .A(n_1174), .B(n_1175), .Y(n_1173) );
CKINVDCx20_ASAP7_75t_R g1178 ( .A(n_1179), .Y(n_1178) );
CKINVDCx20_ASAP7_75t_R g1179 ( .A(n_1180), .Y(n_1179) );
CKINVDCx20_ASAP7_75t_R g1181 ( .A(n_1182), .Y(n_1181) );
endmodule