module fake_jpeg_11420_n_552 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_552);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx8_ASAP7_75t_SL g42 ( 
.A(n_13),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_55),
.B(n_100),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_61),
.B(n_67),
.Y(n_129)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g117 ( 
.A(n_69),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_16),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_76),
.B(n_98),
.Y(n_171)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_24),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_93),
.Y(n_119)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g157 ( 
.A(n_85),
.Y(n_157)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_24),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_33),
.B(n_16),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_25),
.B(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_33),
.B(n_15),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_101),
.B(n_103),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_14),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_107),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_114),
.B(n_136),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_25),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_123),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_83),
.B1(n_75),
.B2(n_19),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_127),
.A2(n_172),
.B1(n_84),
.B2(n_70),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

BUFx16f_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_81),
.A2(n_19),
.B1(n_41),
.B2(n_32),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_36),
.B(n_39),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_25),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_69),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_140),
.B(n_150),
.Y(n_213)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_49),
.Y(n_150)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

BUFx2_ASAP7_75t_SL g221 ( 
.A(n_153),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_49),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_162),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_79),
.B(n_52),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_161),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_52),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_60),
.B(n_38),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_60),
.B(n_38),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_170),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_19),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_56),
.A2(n_41),
.B1(n_37),
.B2(n_27),
.Y(n_172)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_40),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_177),
.B(n_181),
.C(n_204),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_208),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_68),
.C(n_90),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_126),
.A2(n_88),
.B1(n_72),
.B2(n_96),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_182),
.A2(n_186),
.B1(n_191),
.B2(n_194),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_28),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_183),
.B(n_199),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_111),
.A2(n_82),
.B1(n_74),
.B2(n_71),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_185),
.A2(n_230),
.B1(n_145),
.B2(n_159),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_126),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_186)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_188),
.Y(n_241)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_143),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_192),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_193),
.A2(n_195),
.B1(n_184),
.B2(n_204),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_59),
.B1(n_37),
.B2(n_40),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_113),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_203),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_119),
.A2(n_0),
.B(n_1),
.Y(n_198)
);

AO22x1_ASAP7_75t_L g261 ( 
.A1(n_198),
.A2(n_164),
.B1(n_12),
.B2(n_13),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_129),
.B(n_0),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_1),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_225),
.Y(n_255)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_202),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_153),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_51),
.C(n_14),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_205),
.Y(n_285)
);

CKINVDCx12_ASAP7_75t_R g206 ( 
.A(n_157),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_206),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_207),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_1),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_128),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_209),
.B(n_219),
.Y(n_280)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_152),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_117),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_134),
.B(n_3),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_215),
.B(n_223),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_115),
.Y(n_216)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_151),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_218),
.A2(n_222),
.B1(n_234),
.B2(n_11),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_116),
.B(n_3),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_120),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_160),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_6),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_108),
.Y(n_224)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_111),
.B(n_7),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_146),
.B(n_8),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_233),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_125),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_116),
.Y(n_231)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_122),
.Y(n_232)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_146),
.B(n_10),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_160),
.A2(n_173),
.B1(n_124),
.B2(n_154),
.Y(n_234)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_110),
.B(n_13),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_173),
.B(n_154),
.Y(n_252)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_132),
.Y(n_236)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_242),
.B(n_261),
.Y(n_326)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_183),
.B(n_117),
.C(n_109),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_248),
.B(n_228),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_252),
.B(n_273),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_179),
.B(n_115),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_256),
.B(n_281),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_259),
.A2(n_282),
.B1(n_232),
.B2(n_202),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_193),
.A2(n_167),
.B1(n_159),
.B2(n_155),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_263),
.A2(n_236),
.B1(n_188),
.B2(n_175),
.Y(n_300)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_265),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_199),
.B(n_109),
.CI(n_137),
.CON(n_269),
.SN(n_269)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_288),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_164),
.B(n_109),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_271),
.A2(n_201),
.B(n_174),
.Y(n_334)
);

OA22x2_ASAP7_75t_L g273 ( 
.A1(n_178),
.A2(n_139),
.B1(n_155),
.B2(n_145),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_187),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_211),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

FAx1_ASAP7_75t_L g276 ( 
.A(n_198),
.B(n_130),
.CI(n_124),
.CON(n_276),
.SN(n_276)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_205),
.Y(n_307)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_278),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_213),
.B(n_147),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_185),
.A2(n_139),
.B1(n_132),
.B2(n_141),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_181),
.A2(n_167),
.B1(n_141),
.B2(n_130),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_283),
.A2(n_287),
.B1(n_290),
.B2(n_177),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_209),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_225),
.A2(n_11),
.B1(n_12),
.B2(n_229),
.Y(n_290)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_293),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_238),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_294),
.B(n_296),
.Y(n_342)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_257),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_259),
.A2(n_233),
.B1(n_212),
.B2(n_200),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_298),
.A2(n_303),
.B1(n_314),
.B2(n_317),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_180),
.Y(n_299)
);

A2O1A1O1Ixp25_ASAP7_75t_L g365 ( 
.A1(n_299),
.A2(n_328),
.B(n_247),
.C(n_253),
.D(n_228),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_300),
.A2(n_325),
.B1(n_264),
.B2(n_285),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_265),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_302),
.B(n_318),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_266),
.A2(n_226),
.B1(n_190),
.B2(n_176),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_219),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_311),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_307),
.A2(n_334),
.B(n_250),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_268),
.B(n_209),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_255),
.B(n_219),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_255),
.B(n_175),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_315),
.B(n_324),
.Y(n_360)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_316),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_254),
.A2(n_189),
.B1(n_175),
.B2(n_197),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_246),
.B(n_208),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_243),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_319),
.B(n_320),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_260),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

BUFx16f_ASAP7_75t_L g322 ( 
.A(n_258),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_322),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_246),
.A2(n_230),
.B1(n_208),
.B2(n_231),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_323),
.A2(n_335),
.B1(n_317),
.B2(n_327),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_177),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_228),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_260),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_249),
.Y(n_371)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_245),
.Y(n_331)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_241),
.Y(n_332)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_245),
.Y(n_333)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_L g335 ( 
.A1(n_282),
.A2(n_227),
.B1(n_217),
.B2(n_207),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_251),
.Y(n_345)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_338),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_348),
.C(n_351),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_273),
.B1(n_283),
.B2(n_239),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_347),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_280),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_349),
.B(n_368),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_280),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_325),
.A2(n_251),
.B1(n_252),
.B2(n_271),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_359),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_306),
.B(n_248),
.C(n_239),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_373),
.C(n_324),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_327),
.A2(n_239),
.B1(n_273),
.B2(n_269),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_355),
.A2(n_300),
.B1(n_312),
.B2(n_291),
.Y(n_402)
);

NOR2x1_ASAP7_75t_R g359 ( 
.A(n_301),
.B(n_269),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_307),
.A2(n_261),
.B(n_273),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_361),
.A2(n_377),
.B(n_309),
.Y(n_393)
);

AOI32xp33_ASAP7_75t_L g364 ( 
.A1(n_299),
.A2(n_237),
.A3(n_240),
.B1(n_247),
.B2(n_272),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_297),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_365),
.B(n_294),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_285),
.B(n_262),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_370),
.A2(n_376),
.B(n_379),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_371),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_311),
.B(n_249),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_298),
.B(n_250),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_378),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_309),
.A2(n_262),
.B1(n_241),
.B2(n_279),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_326),
.B(n_244),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_328),
.A2(n_244),
.B(n_267),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_371),
.Y(n_380)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_386),
.C(n_387),
.Y(n_443)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_342),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_333),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_391),
.Y(n_435)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_331),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_312),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_394),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_393),
.A2(n_402),
.B1(n_406),
.B2(n_410),
.Y(n_438)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_372),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_396),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_357),
.Y(n_396)
);

INVx13_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g442 ( 
.A(n_397),
.Y(n_442)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_409),
.Y(n_433)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_399),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_345),
.C(n_348),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_340),
.B(n_303),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_401),
.B(n_407),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_376),
.A2(n_313),
.B(n_337),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_403),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_343),
.A2(n_335),
.B1(n_291),
.B2(n_292),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_292),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_375),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_343),
.A2(n_313),
.B1(n_332),
.B2(n_293),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_375),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_412),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_353),
.A2(n_305),
.B(n_338),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_339),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_352),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_357),
.B(n_304),
.Y(n_414)
);

NOR2x1_ASAP7_75t_L g422 ( 
.A(n_414),
.B(n_392),
.Y(n_422)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_352),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_SL g418 ( 
.A(n_390),
.B(n_400),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_431),
.Y(n_452)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_419),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_423),
.C(n_426),
.Y(n_448)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_422),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_383),
.B(n_359),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_390),
.B(n_354),
.C(n_351),
.Y(n_426)
);

HAxp5_ASAP7_75t_SL g427 ( 
.A(n_403),
.B(n_365),
.CON(n_427),
.SN(n_427)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_427),
.A2(n_393),
.B(n_401),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_381),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_430),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_373),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_413),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_432),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_355),
.C(n_379),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_434),
.B(n_444),
.C(n_408),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_322),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_439),
.A2(n_346),
.B1(n_369),
.B2(n_321),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_383),
.B(n_349),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_441),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_388),
.B(n_361),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_370),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_408),
.A2(n_358),
.B1(n_341),
.B2(n_369),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_445),
.A2(n_404),
.B1(n_380),
.B2(n_411),
.Y(n_450)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_408),
.B1(n_405),
.B2(n_402),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_447),
.A2(n_453),
.B1(n_438),
.B2(n_445),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_450),
.A2(n_455),
.B1(n_424),
.B2(n_416),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_425),
.Y(n_451)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_451),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_436),
.A2(n_408),
.B1(n_410),
.B2(n_412),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_382),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_454),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_438),
.A2(n_404),
.B1(n_414),
.B2(n_382),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_468),
.Y(n_488)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_423),
.A2(n_396),
.B(n_385),
.C(n_386),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_464),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_395),
.C(n_385),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_466),
.C(n_471),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_463),
.A2(n_472),
.B(n_305),
.Y(n_485)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_465),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_418),
.B(n_389),
.C(n_384),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_467),
.A2(n_470),
.B1(n_424),
.B2(n_428),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_420),
.B(n_409),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_420),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_398),
.C(n_394),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_444),
.A2(n_415),
.B(n_406),
.Y(n_472)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_474),
.Y(n_506)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_475),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_466),
.A2(n_434),
.B(n_443),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_476),
.B(n_481),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_452),
.B(n_426),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_SL g511 ( 
.A(n_478),
.B(n_490),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_479),
.A2(n_464),
.B1(n_470),
.B2(n_459),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_455),
.A2(n_437),
.B1(n_440),
.B2(n_427),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_480),
.A2(n_468),
.B1(n_457),
.B2(n_454),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_449),
.B(n_422),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_450),
.A2(n_442),
.B1(n_425),
.B2(n_428),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_485),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_441),
.C(n_346),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_487),
.C(n_492),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_458),
.B(n_322),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_484),
.B(n_461),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_341),
.C(n_362),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_358),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_399),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_451),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_448),
.B(n_399),
.C(n_295),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_472),
.A2(n_429),
.B(n_397),
.Y(n_493)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_473),
.Y(n_495)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_495),
.Y(n_514)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_489),
.Y(n_498)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_498),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_491),
.B(n_456),
.C(n_462),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_502),
.C(n_507),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_474),
.A2(n_463),
.B(n_459),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_501),
.A2(n_485),
.B(n_397),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_477),
.B(n_462),
.C(n_467),
.Y(n_502)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_503),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_505),
.A2(n_482),
.B1(n_494),
.B2(n_493),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_453),
.C(n_447),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_508),
.A2(n_486),
.B1(n_479),
.B2(n_494),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_488),
.Y(n_515)
);

XNOR2x1_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_490),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_515),
.Y(n_529)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_513),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_522),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_495),
.A2(n_469),
.B1(n_480),
.B2(n_461),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_518),
.B(n_521),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_488),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_519),
.B(n_520),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_483),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_487),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_502),
.B(n_492),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_524),
.A2(n_509),
.B(n_501),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_513),
.A2(n_497),
.B1(n_506),
.B2(n_505),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_526),
.A2(n_523),
.B1(n_429),
.B2(n_310),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_517),
.A2(n_507),
.B(n_509),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_530),
.A2(n_515),
.B(n_516),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_496),
.C(n_500),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_519),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_517),
.B(n_506),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_534),
.A2(n_535),
.B(n_511),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_536),
.B(n_533),
.C(n_529),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_531),
.A2(n_514),
.B(n_525),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_537),
.A2(n_538),
.B1(n_540),
.B2(n_541),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_539),
.A2(n_528),
.B(n_527),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_527),
.A2(n_512),
.B(n_478),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_542),
.A2(n_544),
.B(n_529),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_545),
.B(n_546),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_543),
.A2(n_535),
.B(n_532),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_526),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_548),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_549),
.B(n_329),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_316),
.C(n_207),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_11),
.Y(n_552)
);


endmodule