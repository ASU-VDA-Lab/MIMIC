module real_aes_7493_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_283;
wire n_252;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
INVx1_ASAP7_75t_L g486 ( .A(n_1), .Y(n_486) );
INVx1_ASAP7_75t_L g199 ( .A(n_2), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_3), .A2(n_102), .B1(n_113), .B2(n_753), .Y(n_101) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_4), .A2(n_38), .B1(n_171), .B2(n_495), .Y(n_494) );
AOI21xp33_ASAP7_75t_L g210 ( .A1(n_5), .A2(n_128), .B(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_6), .B(n_158), .Y(n_478) );
AND2x6_ASAP7_75t_L g133 ( .A(n_7), .B(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_8), .A2(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_9), .B(n_39), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_10), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g216 ( .A(n_11), .Y(n_216) );
INVx1_ASAP7_75t_L g154 ( .A(n_12), .Y(n_154) );
INVx1_ASAP7_75t_L g482 ( .A(n_13), .Y(n_482) );
INVx1_ASAP7_75t_L g187 ( .A(n_14), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_15), .B(n_202), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_16), .B(n_150), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_17), .A2(n_42), .B1(n_724), .B2(n_725), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_17), .Y(n_725) );
AO32x2_ASAP7_75t_L g492 ( .A1(n_18), .A2(n_149), .A3(n_158), .B1(n_464), .B2(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_19), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_20), .B(n_171), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_21), .B(n_144), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_22), .B(n_150), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_23), .A2(n_50), .B1(n_171), .B2(n_495), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g127 ( .A(n_24), .B(n_128), .Y(n_127) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_25), .A2(n_76), .B1(n_171), .B2(n_202), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_26), .B(n_171), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_27), .B(n_209), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_28), .A2(n_184), .B(n_186), .C(n_188), .Y(n_183) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_29), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_30), .B(n_162), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_31), .B(n_169), .Y(n_200) );
INVx1_ASAP7_75t_L g226 ( .A(n_32), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_33), .B(n_162), .Y(n_508) );
INVx2_ASAP7_75t_L g131 ( .A(n_34), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_35), .B(n_171), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_36), .B(n_162), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_37), .A2(n_133), .B(n_136), .C(n_139), .Y(n_135) );
INVx1_ASAP7_75t_L g224 ( .A(n_40), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_41), .B(n_169), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_42), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_43), .B(n_171), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_44), .A2(n_86), .B1(n_147), .B2(n_495), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_45), .B(n_171), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_46), .B(n_171), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_47), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_48), .B(n_462), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_49), .B(n_128), .Y(n_172) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_51), .A2(n_60), .B1(n_171), .B2(n_202), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_52), .A2(n_136), .B1(n_202), .B2(n_223), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_53), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_54), .B(n_171), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_55), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_56), .B(n_171), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_57), .A2(n_214), .B(n_215), .C(n_217), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_58), .Y(n_264) );
INVx1_ASAP7_75t_L g212 ( .A(n_59), .Y(n_212) );
INVx1_ASAP7_75t_L g134 ( .A(n_61), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_62), .B(n_171), .Y(n_487) );
INVx1_ASAP7_75t_L g153 ( .A(n_63), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_64), .Y(n_738) );
AO32x2_ASAP7_75t_L g528 ( .A1(n_65), .A2(n_158), .A3(n_161), .B1(n_464), .B2(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g460 ( .A(n_66), .Y(n_460) );
INVx1_ASAP7_75t_L g503 ( .A(n_67), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_68), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_SL g234 ( .A1(n_69), .A2(n_144), .B(n_217), .C(n_235), .Y(n_234) );
INVxp67_ASAP7_75t_L g236 ( .A(n_70), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_71), .B(n_202), .Y(n_504) );
INVx1_ASAP7_75t_L g106 ( .A(n_72), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_73), .Y(n_229) );
INVx1_ASAP7_75t_L g257 ( .A(n_74), .Y(n_257) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_75), .A2(n_88), .B1(n_744), .B2(n_745), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_75), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_77), .A2(n_133), .B(n_136), .C(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_78), .B(n_495), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_79), .B(n_202), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_80), .B(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g151 ( .A(n_81), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_82), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_83), .B(n_202), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_84), .A2(n_133), .B(n_136), .C(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g108 ( .A(n_85), .B(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g119 ( .A(n_85), .B(n_110), .Y(n_119) );
INVx2_ASAP7_75t_L g447 ( .A(n_85), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_87), .A2(n_100), .B1(n_202), .B2(n_203), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_88), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_89), .B(n_162), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_90), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_91), .A2(n_133), .B(n_136), .C(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_92), .Y(n_174) );
INVx1_ASAP7_75t_L g233 ( .A(n_93), .Y(n_233) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_94), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_95), .B(n_141), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_96), .B(n_202), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_97), .B(n_158), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_98), .B(n_106), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_99), .A2(n_128), .B(n_232), .Y(n_231) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g754 ( .A(n_103), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g746 ( .A(n_108), .Y(n_746) );
INVx1_ASAP7_75t_SL g752 ( .A(n_108), .Y(n_752) );
NOR2x2_ASAP7_75t_L g734 ( .A(n_109), .B(n_447), .Y(n_734) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g446 ( .A(n_110), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AO221x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_736), .B1(n_739), .B2(n_747), .C(n_749), .Y(n_113) );
OAI222xp33_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_723), .B1(n_726), .B2(n_730), .C1(n_731), .C2(n_735), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_120), .B1(n_444), .B2(n_448), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_119), .A2(n_444), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_120), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g741 ( .A1(n_120), .A2(n_728), .B1(n_742), .B2(n_743), .Y(n_741) );
AND2x2_ASAP7_75t_SL g120 ( .A(n_121), .B(n_413), .Y(n_120) );
NOR3xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_306), .C(n_379), .Y(n_121) );
OAI211xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_191), .B(n_238), .C(n_290), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_159), .Y(n_124) );
AND2x2_ASAP7_75t_L g254 ( .A(n_125), .B(n_255), .Y(n_254) );
INVx3_ASAP7_75t_L g273 ( .A(n_125), .Y(n_273) );
INVx2_ASAP7_75t_L g288 ( .A(n_125), .Y(n_288) );
INVx1_ASAP7_75t_L g318 ( .A(n_125), .Y(n_318) );
AND2x2_ASAP7_75t_L g368 ( .A(n_125), .B(n_289), .Y(n_368) );
AOI32xp33_ASAP7_75t_L g395 ( .A1(n_125), .A2(n_323), .A3(n_396), .B1(n_398), .B2(n_399), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_125), .B(n_244), .Y(n_401) );
AND2x2_ASAP7_75t_L g428 ( .A(n_125), .B(n_271), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_125), .B(n_437), .Y(n_436) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_155), .Y(n_125) );
AOI21xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_135), .B(n_148), .Y(n_126) );
BUFx2_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_133), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_129), .B(n_133), .Y(n_196) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
INVx1_ASAP7_75t_L g462 ( .A(n_130), .Y(n_462) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx1_ASAP7_75t_L g203 ( .A(n_131), .Y(n_203) );
INVx1_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
INVx3_ASAP7_75t_L g142 ( .A(n_132), .Y(n_142) );
INVx1_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_132), .Y(n_185) );
INVx4_ASAP7_75t_SL g189 ( .A(n_133), .Y(n_189) );
BUFx3_ASAP7_75t_L g464 ( .A(n_133), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_133), .A2(n_471), .B(n_474), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_133), .A2(n_481), .B(n_485), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_133), .A2(n_502), .B(n_505), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_133), .A2(n_511), .B(n_515), .Y(n_510) );
INVx5_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx3_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_137), .Y(n_171) );
INVx1_ASAP7_75t_L g495 ( .A(n_137), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_143), .B(n_145), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_141), .A2(n_199), .B(n_200), .C(n_201), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_141), .A2(n_457), .B(n_458), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_141), .A2(n_472), .B(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g477 ( .A(n_141), .Y(n_477) );
O2A1O1Ixp5_ASAP7_75t_SL g502 ( .A1(n_141), .A2(n_217), .B(n_503), .C(n_504), .Y(n_502) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_142), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_142), .B(n_236), .Y(n_235) );
OAI22xp5_ASAP7_75t_SL g529 ( .A1(n_142), .A2(n_169), .B1(n_530), .B2(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g514 ( .A(n_144), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_145), .A2(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
INVx1_ASAP7_75t_L g262 ( .A(n_148), .Y(n_262) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_148), .A2(n_455), .B(n_465), .Y(n_454) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_148), .A2(n_480), .B(n_488), .Y(n_479) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_149), .A2(n_194), .B(n_204), .Y(n_193) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_149), .A2(n_221), .B(n_228), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_149), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x2_ASAP7_75t_SL g162 ( .A(n_151), .B(n_152), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx3_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
AO21x1_ASAP7_75t_L g540 ( .A1(n_157), .A2(n_541), .B(n_544), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_157), .B(n_464), .C(n_541), .Y(n_565) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_158), .A2(n_231), .B(n_237), .Y(n_230) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_158), .A2(n_470), .B(n_478), .Y(n_469) );
AND2x2_ASAP7_75t_L g317 ( .A(n_159), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g339 ( .A(n_159), .Y(n_339) );
AND2x2_ASAP7_75t_L g424 ( .A(n_159), .B(n_254), .Y(n_424) );
AND2x2_ASAP7_75t_L g427 ( .A(n_159), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_176), .Y(n_159) );
INVx2_ASAP7_75t_L g246 ( .A(n_160), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_160), .B(n_271), .Y(n_277) );
AND2x2_ASAP7_75t_L g287 ( .A(n_160), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g323 ( .A(n_160), .Y(n_323) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_173), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g175 ( .A(n_162), .Y(n_175) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_162), .A2(n_178), .B(n_190), .Y(n_177) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_162), .A2(n_501), .B(n_508), .Y(n_500) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_162), .A2(n_510), .B(n_518), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_172), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_170), .Y(n_165) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_169), .A2(n_477), .B1(n_494), .B2(n_496), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_169), .A2(n_477), .B1(n_542), .B2(n_543), .Y(n_541) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx3_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_175), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_175), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g265 ( .A(n_176), .B(n_246), .Y(n_265) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g247 ( .A(n_177), .Y(n_247) );
AND2x2_ASAP7_75t_L g289 ( .A(n_177), .B(n_271), .Y(n_289) );
AND2x2_ASAP7_75t_L g358 ( .A(n_177), .B(n_255), .Y(n_358) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .C(n_189), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_182), .A2(n_189), .B(n_212), .C(n_213), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_182), .A2(n_189), .B(n_233), .C(n_234), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_184), .B(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g484 ( .A(n_184), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_184), .A2(n_506), .B(n_507), .Y(n_505) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g223 ( .A1(n_185), .A2(n_224), .B1(n_225), .B2(n_226), .Y(n_223) );
INVx2_ASAP7_75t_L g225 ( .A(n_185), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g221 ( .A1(n_189), .A2(n_196), .B1(n_222), .B2(n_227), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_206), .Y(n_191) );
OR2x2_ASAP7_75t_L g252 ( .A(n_192), .B(n_220), .Y(n_252) );
INVx1_ASAP7_75t_L g331 ( .A(n_192), .Y(n_331) );
AND2x2_ASAP7_75t_L g345 ( .A(n_192), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_192), .B(n_219), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_192), .B(n_343), .Y(n_397) );
AND2x2_ASAP7_75t_L g405 ( .A(n_192), .B(n_406), .Y(n_405) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g242 ( .A(n_193), .Y(n_242) );
AND2x2_ASAP7_75t_L g312 ( .A(n_193), .B(n_220), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_196), .A2(n_257), .B(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_201), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_206), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g439 ( .A(n_206), .Y(n_439) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_219), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_207), .B(n_283), .Y(n_305) );
OR2x2_ASAP7_75t_L g334 ( .A(n_207), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g366 ( .A(n_207), .B(n_346), .Y(n_366) );
INVx1_ASAP7_75t_SL g386 ( .A(n_207), .Y(n_386) );
AND2x2_ASAP7_75t_L g390 ( .A(n_207), .B(n_251), .Y(n_390) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_208), .B(n_219), .Y(n_243) );
AND2x2_ASAP7_75t_L g250 ( .A(n_208), .B(n_230), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_208), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g293 ( .A(n_208), .B(n_275), .Y(n_293) );
INVx1_ASAP7_75t_SL g300 ( .A(n_208), .Y(n_300) );
BUFx2_ASAP7_75t_L g311 ( .A(n_208), .Y(n_311) );
AND2x2_ASAP7_75t_L g327 ( .A(n_208), .B(n_242), .Y(n_327) );
AND2x2_ASAP7_75t_L g342 ( .A(n_208), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g406 ( .A(n_208), .B(n_220), .Y(n_406) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_218), .Y(n_208) );
O2A1O1Ixp5_ASAP7_75t_L g459 ( .A1(n_214), .A2(n_460), .B(n_461), .C(n_463), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_214), .A2(n_516), .B(n_517), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_219), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g330 ( .A(n_219), .B(n_331), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_219), .A2(n_348), .B1(n_351), .B2(n_354), .C(n_359), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_219), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_230), .Y(n_219) );
INVx3_ASAP7_75t_L g275 ( .A(n_220), .Y(n_275) );
BUFx2_ASAP7_75t_L g285 ( .A(n_230), .Y(n_285) );
AND2x2_ASAP7_75t_L g299 ( .A(n_230), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g316 ( .A(n_230), .Y(n_316) );
OR2x2_ASAP7_75t_L g335 ( .A(n_230), .B(n_275), .Y(n_335) );
INVx3_ASAP7_75t_L g343 ( .A(n_230), .Y(n_343) );
AND2x2_ASAP7_75t_L g346 ( .A(n_230), .B(n_275), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_244), .B1(n_248), .B2(n_253), .C(n_266), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_243), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_241), .B(n_315), .Y(n_440) );
OR2x2_ASAP7_75t_L g443 ( .A(n_241), .B(n_274), .Y(n_443) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
OAI221xp5_ASAP7_75t_SL g266 ( .A1(n_242), .A2(n_267), .B1(n_274), .B2(n_276), .C(n_279), .Y(n_266) );
AND2x2_ASAP7_75t_L g283 ( .A(n_242), .B(n_275), .Y(n_283) );
AND2x2_ASAP7_75t_L g291 ( .A(n_242), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_242), .B(n_299), .Y(n_298) );
NAND2x1_ASAP7_75t_L g341 ( .A(n_242), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g393 ( .A(n_242), .B(n_335), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_244), .A2(n_353), .B1(n_382), .B2(n_384), .Y(n_381) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AOI322xp5_ASAP7_75t_L g290 ( .A1(n_245), .A2(n_254), .A3(n_291), .B1(n_294), .B2(n_297), .C1(n_301), .C2(n_304), .Y(n_290) );
OR2x2_ASAP7_75t_L g302 ( .A(n_245), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_246), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g281 ( .A(n_246), .B(n_255), .Y(n_281) );
INVx1_ASAP7_75t_L g296 ( .A(n_246), .Y(n_296) );
AND2x2_ASAP7_75t_L g362 ( .A(n_246), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g272 ( .A(n_247), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g363 ( .A(n_247), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_247), .B(n_271), .Y(n_437) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_251), .B(n_386), .Y(n_385) );
INVx3_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g337 ( .A(n_252), .B(n_284), .Y(n_337) );
OR2x2_ASAP7_75t_L g434 ( .A(n_252), .B(n_285), .Y(n_434) );
INVx1_ASAP7_75t_L g415 ( .A(n_253), .Y(n_415) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_265), .Y(n_253) );
INVx4_ASAP7_75t_L g303 ( .A(n_254), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_254), .B(n_322), .Y(n_328) );
INVx2_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_262), .B(n_263), .Y(n_255) );
INVx1_ASAP7_75t_L g353 ( .A(n_265), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_265), .B(n_325), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g340 ( .A1(n_267), .A2(n_341), .B(n_344), .Y(n_340) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g325 ( .A(n_271), .Y(n_325) );
INVx1_ASAP7_75t_L g352 ( .A(n_271), .Y(n_352) );
INVx1_ASAP7_75t_L g278 ( .A(n_272), .Y(n_278) );
AND2x2_ASAP7_75t_L g280 ( .A(n_272), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g376 ( .A(n_273), .B(n_362), .Y(n_376) );
AND2x2_ASAP7_75t_L g398 ( .A(n_273), .B(n_358), .Y(n_398) );
BUFx2_ASAP7_75t_L g350 ( .A(n_275), .Y(n_350) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AOI32xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_282), .A3(n_283), .B1(n_284), .B2(n_286), .Y(n_279) );
INVx1_ASAP7_75t_L g360 ( .A(n_280), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_280), .A2(n_408), .B1(n_409), .B2(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_283), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_283), .B(n_342), .Y(n_383) );
AND2x2_ASAP7_75t_L g430 ( .A(n_283), .B(n_315), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_284), .B(n_331), .Y(n_378) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g431 ( .A(n_286), .Y(n_431) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g356 ( .A(n_287), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_289), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g403 ( .A(n_289), .B(n_323), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_289), .B(n_318), .Y(n_410) );
INVx1_ASAP7_75t_SL g392 ( .A(n_291), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_292), .B(n_343), .Y(n_370) );
NOR4xp25_ASAP7_75t_L g416 ( .A(n_292), .B(n_315), .C(n_417), .D(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_293), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVxp67_ASAP7_75t_L g373 ( .A(n_296), .Y(n_373) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI21xp33_ASAP7_75t_L g423 ( .A1(n_299), .A2(n_390), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g315 ( .A(n_300), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g364 ( .A(n_303), .Y(n_364) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND4xp25_ASAP7_75t_SL g306 ( .A(n_307), .B(n_332), .C(n_347), .D(n_367), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_313), .B(n_317), .C(n_319), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g399 ( .A(n_312), .B(n_342), .Y(n_399) );
AND2x2_ASAP7_75t_L g408 ( .A(n_312), .B(n_386), .Y(n_408) );
INVx3_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_315), .B(n_350), .Y(n_412) );
AND2x2_ASAP7_75t_L g324 ( .A(n_318), .B(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_326), .B1(n_328), .B2(n_329), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
AND2x2_ASAP7_75t_L g422 ( .A(n_322), .B(n_368), .Y(n_422) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_324), .B(n_373), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_325), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_336), .B(n_338), .C(n_340), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_333), .A2(n_368), .B1(n_369), .B2(n_371), .C(n_374), .Y(n_367) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_341), .A2(n_426), .B1(n_429), .B2(n_431), .C(n_432), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_342), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_350), .B(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g380 ( .A(n_352), .Y(n_380) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_355), .A2(n_375), .B1(n_377), .B2(n_378), .Y(n_374) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI21xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B(n_365), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_364), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_375), .A2(n_401), .B1(n_439), .B2(n_440), .C(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g420 ( .A(n_377), .Y(n_420) );
OAI211xp5_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_381), .B(n_387), .C(n_407), .Y(n_379) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI211xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_391), .C(n_400), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_394), .C(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g419 ( .A(n_397), .Y(n_419) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_398), .A2(n_424), .B(n_442), .Y(n_441) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_404), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g433 ( .A1(n_410), .A2(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_425), .C(n_438), .Y(n_413) );
OAI211xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B(n_421), .C(n_423), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
CKINVDCx14_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g729 ( .A(n_448), .Y(n_729) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_651), .C(n_700), .Y(n_449) );
NAND5xp2_ASAP7_75t_L g450 ( .A(n_451), .B(n_566), .C(n_594), .D(n_624), .E(n_638), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_489), .B1(n_519), .B2(n_524), .C(n_533), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_466), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_453), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g546 ( .A(n_454), .Y(n_546) );
AND2x2_ASAP7_75t_L g554 ( .A(n_454), .B(n_469), .Y(n_554) );
AND2x2_ASAP7_75t_L g577 ( .A(n_454), .B(n_468), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_454), .B(n_479), .Y(n_592) );
OR2x2_ASAP7_75t_L g601 ( .A(n_454), .B(n_540), .Y(n_601) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_454), .Y(n_604) );
AND2x2_ASAP7_75t_L g712 ( .A(n_454), .B(n_540), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_459), .B(n_464), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_461), .A2(n_477), .B(n_486), .C(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_466), .B(n_604), .Y(n_660) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
OAI311xp33_ASAP7_75t_L g602 ( .A1(n_467), .A2(n_603), .A3(n_604), .B1(n_605), .C1(n_620), .Y(n_602) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_479), .Y(n_467) );
AND2x2_ASAP7_75t_L g563 ( .A(n_468), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g570 ( .A(n_468), .Y(n_570) );
AND2x2_ASAP7_75t_L g691 ( .A(n_468), .B(n_523), .Y(n_691) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_469), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g547 ( .A(n_469), .B(n_479), .Y(n_547) );
AND2x2_ASAP7_75t_L g599 ( .A(n_469), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g613 ( .A(n_469), .B(n_546), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_477), .Y(n_474) );
INVx2_ASAP7_75t_L g523 ( .A(n_479), .Y(n_523) );
AND2x2_ASAP7_75t_L g562 ( .A(n_479), .B(n_546), .Y(n_562) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_497), .Y(n_489) );
OR2x2_ASAP7_75t_L g657 ( .A(n_490), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_490), .B(n_663), .Y(n_674) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_491), .B(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g532 ( .A(n_492), .Y(n_532) );
AND2x2_ASAP7_75t_L g598 ( .A(n_492), .B(n_528), .Y(n_598) );
AND2x2_ASAP7_75t_L g609 ( .A(n_492), .B(n_509), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_492), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_497), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_497), .B(n_559), .Y(n_603) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g590 ( .A(n_498), .B(n_549), .Y(n_590) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_509), .Y(n_498) );
INVx2_ASAP7_75t_L g526 ( .A(n_499), .Y(n_526) );
AND2x2_ASAP7_75t_L g617 ( .A(n_499), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g536 ( .A(n_500), .Y(n_536) );
OR2x2_ASAP7_75t_L g634 ( .A(n_500), .B(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_500), .Y(n_697) );
AND2x2_ASAP7_75t_L g537 ( .A(n_509), .B(n_532), .Y(n_537) );
INVx1_ASAP7_75t_L g557 ( .A(n_509), .Y(n_557) );
AND2x2_ASAP7_75t_L g578 ( .A(n_509), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g619 ( .A(n_509), .Y(n_619) );
INVx1_ASAP7_75t_L g635 ( .A(n_509), .Y(n_635) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_509), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_514), .Y(n_511) );
INVxp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_521), .B(n_623), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_521), .A2(n_608), .B1(n_657), .B2(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
OAI211xp5_ASAP7_75t_SL g700 ( .A1(n_522), .A2(n_701), .B(n_703), .C(n_721), .Y(n_700) );
INVx2_ASAP7_75t_L g553 ( .A(n_523), .Y(n_553) );
AND2x2_ASAP7_75t_L g611 ( .A(n_523), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g622 ( .A(n_523), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_524), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
AND2x2_ASAP7_75t_L g595 ( .A(n_525), .B(n_559), .Y(n_595) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g627 ( .A(n_526), .B(n_618), .Y(n_627) );
AND2x2_ASAP7_75t_L g646 ( .A(n_526), .B(n_560), .Y(n_646) );
AND2x4_ASAP7_75t_L g582 ( .A(n_527), .B(n_556), .Y(n_582) );
AND2x2_ASAP7_75t_L g720 ( .A(n_527), .B(n_696), .Y(n_720) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .Y(n_527) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_528), .Y(n_549) );
INVx1_ASAP7_75t_L g560 ( .A(n_528), .Y(n_560) );
INVx1_ASAP7_75t_L g659 ( .A(n_528), .Y(n_659) );
OR2x2_ASAP7_75t_L g550 ( .A(n_532), .B(n_536), .Y(n_550) );
AND2x2_ASAP7_75t_L g559 ( .A(n_532), .B(n_560), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g579 ( .A(n_532), .B(n_580), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_538), .B1(n_548), .B2(n_551), .C(n_555), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_535), .A2(n_556), .B(n_558), .C(n_561), .Y(n_555) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g580 ( .A(n_536), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_536), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_SL g663 ( .A(n_536), .B(n_557), .Y(n_663) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_536), .Y(n_670) );
AND2x2_ASAP7_75t_L g588 ( .A(n_537), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g625 ( .A(n_537), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_547), .Y(n_538) );
INVx2_ASAP7_75t_L g616 ( .A(n_539), .Y(n_616) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_539), .A2(n_549), .B1(n_666), .B2(n_668), .C1(n_669), .C2(n_671), .Y(n_665) );
AND2x2_ASAP7_75t_L g722 ( .A(n_539), .B(n_691), .Y(n_722) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_546), .Y(n_539) );
INVx1_ASAP7_75t_L g612 ( .A(n_540), .Y(n_612) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g564 ( .A(n_545), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g650 ( .A(n_547), .B(n_584), .Y(n_650) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_548), .A2(n_662), .B(n_664), .Y(n_661) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g589 ( .A(n_549), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_549), .B(n_556), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_549), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx3_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
OR2x2_ASAP7_75t_L g667 ( .A(n_553), .B(n_589), .Y(n_667) );
AND2x2_ASAP7_75t_L g583 ( .A(n_554), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g621 ( .A(n_554), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_554), .B(n_615), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_554), .B(n_611), .Y(n_637) );
AND2x2_ASAP7_75t_L g641 ( .A(n_554), .B(n_623), .Y(n_641) );
INVxp67_ASAP7_75t_L g573 ( .A(n_556), .Y(n_573) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_558), .A2(n_631), .B1(n_636), .B2(n_637), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_558), .B(n_663), .Y(n_693) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g679 ( .A(n_559), .B(n_670), .Y(n_679) );
AND2x2_ASAP7_75t_L g708 ( .A(n_559), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g713 ( .A(n_559), .B(n_663), .Y(n_713) );
INVx1_ASAP7_75t_L g626 ( .A(n_560), .Y(n_626) );
BUFx2_ASAP7_75t_L g632 ( .A(n_560), .Y(n_632) );
INVx1_ASAP7_75t_L g717 ( .A(n_561), .Y(n_717) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_562), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g593 ( .A(n_563), .Y(n_593) );
NOR2x1_ASAP7_75t_L g569 ( .A(n_564), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g576 ( .A(n_564), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g585 ( .A(n_564), .Y(n_585) );
INVx3_ASAP7_75t_L g623 ( .A(n_564), .Y(n_623) );
OR2x2_ASAP7_75t_L g689 ( .A(n_564), .B(n_690), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_571), .B(n_574), .C(n_586), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_567), .A2(n_704), .B1(n_711), .B2(n_713), .C(n_714), .Y(n_703) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_575), .B(n_581), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_577), .B(n_615), .Y(n_629) );
AND2x2_ASAP7_75t_L g671 ( .A(n_577), .B(n_611), .Y(n_671) );
INVx1_ASAP7_75t_SL g684 ( .A(n_578), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_578), .B(n_632), .Y(n_687) );
INVx1_ASAP7_75t_L g705 ( .A(n_579), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_583), .A2(n_673), .B1(n_675), .B2(n_679), .C(n_680), .Y(n_672) );
AND2x2_ASAP7_75t_L g699 ( .A(n_584), .B(n_691), .Y(n_699) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g683 ( .A(n_585), .Y(n_683) );
AOI21xp33_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_590), .B(n_591), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g654 ( .A(n_589), .B(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g640 ( .A(n_590), .Y(n_640) );
INVx1_ASAP7_75t_L g668 ( .A(n_591), .Y(n_668) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_599), .C(n_602), .Y(n_594) );
OAI31xp33_ASAP7_75t_L g721 ( .A1(n_595), .A2(n_633), .A3(n_720), .B(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g695 ( .A(n_598), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g716 ( .A(n_598), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_600), .B(n_615), .Y(n_643) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g718 ( .A(n_601), .B(n_615), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_610), .B1(n_614), .B2(n_617), .Y(n_605) );
NAND2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_609), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g645 ( .A(n_609), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g648 ( .A(n_609), .B(n_632), .Y(n_648) );
AND2x2_ASAP7_75t_L g702 ( .A(n_609), .B(n_697), .Y(n_702) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g677 ( .A(n_613), .Y(n_677) );
NOR2xp67_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OAI32xp33_ASAP7_75t_L g680 ( .A1(n_615), .A2(n_649), .A3(n_681), .B1(n_683), .B2(n_684), .Y(n_680) );
INVx1_ASAP7_75t_L g655 ( .A(n_618), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_618), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g678 ( .A(n_622), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_628), .C(n_630), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_626), .B(n_663), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_627), .A2(n_639), .B1(n_640), .B2(n_641), .C(n_642), .Y(n_638) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g639 ( .A(n_637), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B1(n_647), .B2(n_649), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND4xp25_ASAP7_75t_SL g704 ( .A(n_647), .B(n_705), .C(n_706), .D(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NAND4xp25_ASAP7_75t_SL g651 ( .A(n_652), .B(n_665), .C(n_672), .D(n_685), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B(n_660), .C(n_661), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g682 ( .A(n_658), .Y(n_682) );
INVx2_ASAP7_75t_L g706 ( .A(n_663), .Y(n_706) );
OR2x2_ASAP7_75t_L g715 ( .A(n_670), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_692), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g711 ( .A(n_691), .B(n_712), .Y(n_711) );
AOI21xp33_ASAP7_75t_SL g692 ( .A1(n_693), .A2(n_694), .B(n_698), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
CKINVDCx16_ASAP7_75t_R g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g730 ( .A(n_723), .Y(n_730) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g748 ( .A(n_737), .Y(n_748) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_741), .B(n_746), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx3_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
endmodule