module fake_netlist_6_2754_n_2249 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2249);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2249;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_343;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_811;
wire n_683;
wire n_527;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_374;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g230 ( 
.A(n_51),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_127),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_99),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_154),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_11),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_3),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_163),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_196),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_92),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_75),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_3),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_124),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_114),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_105),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_30),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_54),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_194),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_55),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_198),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_197),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_161),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_51),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_125),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_119),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_8),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_150),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_100),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_180),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_96),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_167),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_184),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_188),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_126),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_116),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_113),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_98),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_143),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_56),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_72),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_11),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_219),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_65),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_120),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_136),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_133),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_187),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_166),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_66),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_28),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_228),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_215),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_21),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_141),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_201),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_15),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_27),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_176),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_227),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_7),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_203),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_151),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_213),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_22),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_89),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_142),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_204),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_190),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_72),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_24),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_5),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_131),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_24),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_36),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_128),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_68),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_206),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_172),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_101),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_115),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_217),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_71),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_108),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_73),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_224),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_43),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_66),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_186),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_153),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_156),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_37),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_28),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_169),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_10),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_159),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_57),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_56),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_69),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_175),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_210),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_55),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_199),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_57),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_111),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_26),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_84),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_58),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_14),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_18),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_34),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_83),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_147),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_192),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_207),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_129),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_157),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_134),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_94),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_60),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_162),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_44),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_10),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_90),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_29),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_220),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_149),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_23),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_86),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_109),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_123),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_82),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_145),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_77),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_173),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_205),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_40),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_202),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_46),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_200),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_222),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_195),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_37),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_121),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_43),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_138),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_0),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_53),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_87),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_189),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_68),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_76),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_35),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_211),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_107),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_155),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_117),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_21),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_64),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_60),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_209),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_39),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_15),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_178),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_40),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_122),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_171),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_9),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_38),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_160),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_78),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_49),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_177),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_165),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_104),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_23),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_181),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_221),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_54),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_16),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_31),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_183),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_19),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_34),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_140),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_39),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_110),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_59),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_112),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_106),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_62),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_7),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_118),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_71),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_79),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_182),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_38),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_139),
.Y(n_436)
);

BUFx5_ASAP7_75t_L g437 ( 
.A(n_30),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_52),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_4),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_9),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_97),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_80),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_62),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_132),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_33),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_229),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_52),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_59),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_29),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_148),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_61),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_447),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_295),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_437),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_247),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_280),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_298),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_299),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_437),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_276),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_437),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_437),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_437),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_285),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_308),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_321),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_434),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_363),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_315),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_303),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_303),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_303),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_325),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_303),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_303),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_310),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_310),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_310),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_284),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_310),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_254),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_274),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_310),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_351),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_236),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_330),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_331),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_363),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_230),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_352),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_235),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_335),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_340),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_277),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_288),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_291),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_342),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_294),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_309),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_312),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_333),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_336),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_337),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_297),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_361),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_344),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_375),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_377),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_400),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_287),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_403),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_410),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_419),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_425),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_429),
.Y(n_524)
);

INVxp33_ASAP7_75t_SL g525 ( 
.A(n_236),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_287),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_430),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_440),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_448),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_241),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_451),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_346),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_284),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_319),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_347),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_319),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_345),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_345),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_367),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_399),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_313),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_248),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_399),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_233),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_241),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_241),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_244),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_313),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_245),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_246),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_255),
.Y(n_551)
);

INVxp33_ASAP7_75t_SL g552 ( 
.A(n_248),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_348),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_256),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_450),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_349),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_241),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_265),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_449),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_266),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_358),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_231),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_231),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_270),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_238),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_238),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_273),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_318),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_381),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_273),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_385),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_318),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_449),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_482),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_456),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_530),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_557),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_474),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_540),
.B(n_318),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_455),
.B(n_250),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_530),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_474),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_475),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_475),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_477),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_530),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_452),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_545),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_456),
.Y(n_591)
);

CKINVDCx6p67_ASAP7_75t_R g592 ( 
.A(n_568),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_564),
.B(n_290),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_557),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_473),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_457),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_477),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_544),
.B(n_547),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_484),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_452),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_473),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_545),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_480),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_549),
.B(n_290),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_550),
.B(n_365),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_R g606 ( 
.A(n_457),
.B(n_232),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_458),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_478),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_472),
.A2(n_252),
.B1(n_406),
.B2(n_360),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_458),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_468),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_470),
.B(n_365),
.Y(n_612)
);

OAI22x1_ASAP7_75t_L g613 ( 
.A1(n_467),
.A2(n_249),
.B1(n_260),
.B2(n_257),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_453),
.A2(n_438),
.B1(n_424),
.B2(n_323),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_545),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_480),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_478),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_468),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_459),
.A2(n_301),
.B(n_281),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_533),
.B(n_293),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_485),
.A2(n_249),
.B1(n_260),
.B2(n_257),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_534),
.B(n_316),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_491),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_551),
.B(n_281),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_545),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_482),
.B(n_301),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_512),
.B(n_387),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_554),
.B(n_427),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_469),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_487),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_469),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_491),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_558),
.B(n_232),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_560),
.B(n_427),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_545),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_546),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_498),
.A2(n_435),
.B1(n_445),
.B2(n_421),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_479),
.B(n_292),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_546),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_546),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_536),
.B(n_234),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_546),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_546),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_461),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_462),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_476),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_476),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_479),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_481),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_523),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_555),
.A2(n_435),
.B1(n_445),
.B2(n_421),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_460),
.B(n_241),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_537),
.B(n_234),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_463),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_481),
.Y(n_655)
);

BUFx8_ASAP7_75t_L g656 ( 
.A(n_538),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_494),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_483),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_464),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_543),
.B(n_237),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_494),
.B(n_267),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_465),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_466),
.A2(n_300),
.B(n_296),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_483),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_486),
.B(n_237),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_486),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_488),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_488),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_606),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_658),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_658),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_627),
.B(n_489),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_652),
.B(n_572),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_595),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_658),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_595),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_593),
.B(n_626),
.C(n_605),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_599),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_595),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_652),
.B(n_495),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_601),
.Y(n_681)
);

CKINVDCx6p67_ASAP7_75t_R g682 ( 
.A(n_592),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_590),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_644),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_644),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_644),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_667),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_601),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_SL g689 ( 
.A(n_613),
.B(n_495),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_601),
.Y(n_690)
);

INVxp33_ASAP7_75t_SL g691 ( 
.A(n_581),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_645),
.Y(n_692)
);

BUFx6f_ASAP7_75t_SL g693 ( 
.A(n_652),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_645),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_580),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_631),
.B(n_500),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_603),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_631),
.B(n_500),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_603),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_574),
.B(n_489),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_574),
.B(n_490),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_603),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_SL g703 ( 
.A1(n_621),
.A2(n_539),
.B1(n_552),
.B2(n_525),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_645),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_620),
.B(n_501),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_616),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_581),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_612),
.B(n_525),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_593),
.A2(n_552),
.B1(n_454),
.B2(n_493),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_616),
.Y(n_710)
);

AO21x2_ASAP7_75t_L g711 ( 
.A1(n_663),
.A2(n_306),
.B(n_305),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_580),
.B(n_490),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_616),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_620),
.B(n_501),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_654),
.Y(n_715)
);

INVx6_ASAP7_75t_L g716 ( 
.A(n_577),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_654),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_623),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_654),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_622),
.B(n_665),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_622),
.B(n_505),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_624),
.A2(n_634),
.B1(n_628),
.B2(n_638),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_659),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_623),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_590),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_623),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_590),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_659),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_632),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_667),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_632),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_632),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_665),
.B(n_492),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_578),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_659),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_638),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_621),
.A2(n_326),
.B1(n_366),
.B2(n_242),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_661),
.B(n_505),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_578),
.Y(n_739)
);

NOR2x1p5_ASAP7_75t_L g740 ( 
.A(n_592),
.B(n_267),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_590),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_578),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_662),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_594),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_641),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

BUFx6f_ASAP7_75t_SL g747 ( 
.A(n_598),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_662),
.B(n_492),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_590),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_662),
.B(n_454),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_590),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_594),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_624),
.A2(n_563),
.B1(n_565),
.B2(n_562),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_625),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_579),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_624),
.A2(n_563),
.B1(n_565),
.B2(n_562),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_624),
.A2(n_567),
.B1(n_570),
.B2(n_566),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_579),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_638),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_641),
.B(n_514),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_583),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_653),
.B(n_542),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_583),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_584),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_584),
.Y(n_765)
);

OAI21xp33_ASAP7_75t_SL g766 ( 
.A1(n_619),
.A2(n_605),
.B(n_604),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_585),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_625),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_638),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_653),
.B(n_514),
.Y(n_770)
);

INVx6_ASAP7_75t_L g771 ( 
.A(n_577),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_585),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_598),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_575),
.B(n_532),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_625),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_586),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_586),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_597),
.Y(n_778)
);

INVx5_ASAP7_75t_L g779 ( 
.A(n_625),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_597),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_660),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_625),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_608),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_660),
.B(n_532),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_598),
.B(n_518),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_608),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_598),
.B(n_535),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_617),
.Y(n_788)
);

CKINVDCx16_ASAP7_75t_R g789 ( 
.A(n_588),
.Y(n_789)
);

BUFx4f_ASAP7_75t_L g790 ( 
.A(n_667),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_617),
.Y(n_791)
);

NOR2x1p5_ASAP7_75t_L g792 ( 
.A(n_591),
.B(n_275),
.Y(n_792)
);

AND3x2_ASAP7_75t_L g793 ( 
.A(n_618),
.B(n_573),
.C(n_559),
.Y(n_793)
);

INVxp33_ASAP7_75t_SL g794 ( 
.A(n_609),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_648),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_649),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_633),
.B(n_535),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_576),
.B(n_553),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_633),
.B(n_553),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_630),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_596),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_649),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_655),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_618),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_L g805 ( 
.A(n_607),
.B(n_571),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_667),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_655),
.Y(n_807)
);

BUFx4f_ASAP7_75t_L g808 ( 
.A(n_667),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_664),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_SL g810 ( 
.A1(n_637),
.A2(n_278),
.B1(n_414),
.B2(n_275),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_611),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_637),
.A2(n_383),
.B1(n_414),
.B2(n_278),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_625),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_635),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_650),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_664),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_635),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_666),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_666),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_668),
.Y(n_820)
);

AND2x6_ASAP7_75t_L g821 ( 
.A(n_628),
.B(n_264),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_635),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_635),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_668),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_613),
.A2(n_389),
.B1(n_391),
.B2(n_386),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_619),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_628),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_629),
.B(n_556),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_745),
.B(n_556),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_695),
.B(n_646),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_674),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_745),
.B(n_561),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_695),
.B(n_657),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_785),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_798),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_781),
.B(n_561),
.Y(n_836)
);

NAND2x1_ASAP7_75t_L g837 ( 
.A(n_716),
.B(n_577),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_720),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_670),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_674),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_773),
.B(n_497),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_781),
.B(n_569),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_677),
.B(n_569),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_797),
.B(n_610),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_677),
.B(n_760),
.Y(n_845)
);

NAND2xp33_ASAP7_75t_L g846 ( 
.A(n_669),
.B(n_647),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_762),
.B(n_799),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_804),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_737),
.A2(n_614),
.B1(n_609),
.B2(n_604),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_669),
.B(n_762),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_770),
.B(n_784),
.Y(n_851)
);

AOI22x1_ASAP7_75t_L g852 ( 
.A1(n_671),
.A2(n_571),
.B1(n_600),
.B2(n_628),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_705),
.B(n_651),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_676),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_676),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_733),
.B(n_634),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_672),
.B(n_827),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_827),
.B(n_634),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_671),
.B(n_634),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_679),
.Y(n_860)
);

BUFx8_ASAP7_75t_L g861 ( 
.A(n_811),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_714),
.B(n_651),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_675),
.B(n_577),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_675),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_L g865 ( 
.A(n_787),
.B(n_279),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_721),
.B(n_409),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_736),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_736),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_804),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_738),
.B(n_656),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_709),
.B(n_614),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_811),
.B(n_471),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_680),
.A2(n_528),
.B(n_522),
.C(n_566),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_736),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_766),
.A2(n_663),
.B(n_324),
.C(n_327),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_759),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_708),
.B(n_656),
.C(n_496),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_773),
.B(n_656),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_712),
.B(n_576),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_759),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_773),
.B(n_499),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_679),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_681),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_759),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_769),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_774),
.B(n_502),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_769),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_673),
.B(n_239),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_696),
.B(n_656),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_681),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_707),
.B(n_503),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_722),
.B(n_576),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_678),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_698),
.B(n_239),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_769),
.B(n_240),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_693),
.A2(n_283),
.B1(n_286),
.B2(n_282),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_693),
.A2(n_370),
.B1(n_369),
.B2(n_368),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_755),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_755),
.B(n_576),
.Y(n_899)
);

INVx8_ASAP7_75t_L g900 ( 
.A(n_693),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_764),
.B(n_582),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_826),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_SL g903 ( 
.A(n_682),
.B(n_240),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_764),
.B(n_582),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_765),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_794),
.B(n_243),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_765),
.B(n_582),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_688),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_801),
.B(n_504),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_R g910 ( 
.A(n_815),
.B(n_289),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_688),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_L g912 ( 
.A(n_821),
.B(n_302),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_772),
.B(n_582),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_772),
.B(n_587),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_800),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_776),
.B(n_587),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_825),
.B(n_243),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_786),
.B(n_251),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_826),
.A2(n_570),
.B1(n_567),
.B2(n_264),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_786),
.B(n_587),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_826),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_801),
.B(n_251),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_740),
.B(n_506),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_795),
.B(n_589),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_795),
.B(n_253),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_790),
.A2(n_643),
.B(n_635),
.Y(n_926)
);

NAND2x1_ASAP7_75t_L g927 ( 
.A(n_716),
.B(n_771),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_796),
.B(n_253),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_690),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_796),
.B(n_802),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_689),
.A2(n_339),
.B1(n_332),
.B2(n_328),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_700),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_716),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_802),
.B(n_589),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_809),
.B(n_589),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_701),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_809),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_805),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_801),
.B(n_507),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_819),
.B(n_602),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_801),
.B(n_258),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_819),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_758),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_703),
.B(n_258),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_747),
.A2(n_388),
.B1(n_317),
.B2(n_311),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_690),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_810),
.A2(n_307),
.B1(n_264),
.B2(n_404),
.Y(n_947)
);

AOI221xp5_ASAP7_75t_L g948 ( 
.A1(n_737),
.A2(n_439),
.B1(n_432),
.B2(n_443),
.C(n_422),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_820),
.B(n_259),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_828),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_758),
.B(n_602),
.Y(n_951)
);

BUFx5_ASAP7_75t_L g952 ( 
.A(n_684),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_L g953 ( 
.A(n_821),
.B(n_304),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_761),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_751),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_761),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_763),
.B(n_602),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_792),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_SL g959 ( 
.A(n_716),
.B(n_264),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_789),
.B(n_259),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_747),
.B(n_824),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_747),
.A2(n_359),
.B1(n_433),
.B2(n_329),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_711),
.A2(n_264),
.B1(n_307),
.B2(n_412),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_763),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_767),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_767),
.B(n_261),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_792),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_777),
.B(n_602),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_789),
.B(n_261),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_824),
.B(n_262),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_793),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_777),
.B(n_778),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_697),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_800),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_790),
.A2(n_643),
.B(n_635),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_SL g976 ( 
.A(n_682),
.B(n_262),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_L g977 ( 
.A(n_766),
.B(n_508),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_740),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_778),
.B(n_667),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_L g980 ( 
.A(n_812),
.B(n_390),
.C(n_314),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_753),
.B(n_263),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_707),
.B(n_509),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_780),
.B(n_393),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_697),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_751),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_683),
.B(n_320),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_756),
.B(n_263),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_780),
.B(n_636),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_783),
.B(n_636),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_783),
.A2(n_436),
.B1(n_431),
.B2(n_405),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_788),
.B(n_636),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_699),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_757),
.B(n_268),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_812),
.B(n_510),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_699),
.Y(n_995)
);

OAI21xp33_ASAP7_75t_L g996 ( 
.A1(n_788),
.A2(n_513),
.B(n_511),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_791),
.B(n_639),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_791),
.B(n_268),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_841),
.B(n_803),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_841),
.B(n_881),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_851),
.B(n_803),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_943),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_881),
.B(n_807),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_834),
.B(n_807),
.Y(n_1004)
);

AO21x1_ASAP7_75t_L g1005 ( 
.A1(n_845),
.A2(n_402),
.B(n_684),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_943),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_921),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_847),
.B(n_816),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_838),
.A2(n_816),
.B(n_818),
.C(n_750),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_954),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_848),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_891),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_956),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_SL g1014 ( 
.A(n_861),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_964),
.Y(n_1015)
);

NAND2x2_ASAP7_75t_L g1016 ( 
.A(n_978),
.B(n_417),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_965),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_982),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_839),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_876),
.B(n_818),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_893),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_847),
.B(n_685),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_838),
.B(n_685),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_872),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_921),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_SL g1026 ( 
.A1(n_871),
.A2(n_691),
.B1(n_443),
.B2(n_418),
.Y(n_1026)
);

NOR2x1p5_ASAP7_75t_L g1027 ( 
.A(n_829),
.B(n_417),
.Y(n_1027)
);

OAI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_853),
.A2(n_862),
.B1(n_857),
.B2(n_849),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_864),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_876),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_831),
.Y(n_1031)
);

OR2x6_ASAP7_75t_L g1032 ( 
.A(n_900),
.B(n_515),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_909),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_835),
.A2(n_771),
.B1(n_821),
.B2(n_692),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_921),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_932),
.B(n_686),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_869),
.Y(n_1037)
);

AND3x2_ASAP7_75t_SL g1038 ( 
.A(n_947),
.B(n_526),
.C(n_518),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_869),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_932),
.B(n_686),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_876),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_900),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_921),
.Y(n_1043)
);

INVx8_ASAP7_75t_L g1044 ( 
.A(n_900),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_936),
.B(n_692),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_840),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_876),
.B(n_694),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_861),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_939),
.B(n_516),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_963),
.A2(n_771),
.B1(n_694),
.B2(n_719),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_933),
.B(n_704),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_915),
.Y(n_1052)
);

OAI22x1_ASAP7_75t_R g1053 ( 
.A1(n_853),
.A2(n_418),
.B1(n_432),
.B2(n_422),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_898),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_854),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_936),
.B(n_704),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_933),
.B(n_715),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_905),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_974),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_930),
.B(n_715),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_930),
.B(n_717),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_937),
.B(n_717),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_906),
.B(n_719),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_927),
.A2(n_808),
.B(n_790),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_967),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_867),
.B(n_517),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_942),
.B(n_723),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_977),
.A2(n_728),
.B(n_723),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_868),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_843),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_955),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_980),
.A2(n_711),
.B1(n_821),
.B2(n_728),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_902),
.B(n_735),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_862),
.A2(n_771),
.B1(n_821),
.B2(n_735),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_910),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_923),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_972),
.Y(n_1077)
);

INVx5_ASAP7_75t_L g1078 ( 
.A(n_902),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_980),
.A2(n_711),
.B1(n_821),
.B2(n_743),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_971),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_832),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_874),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_880),
.B(n_884),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_923),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_856),
.B(n_743),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_L g1086 ( 
.A(n_906),
.B(n_271),
.C(n_269),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_885),
.Y(n_1087)
);

INVx5_ASAP7_75t_L g1088 ( 
.A(n_955),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_855),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_923),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_938),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_837),
.A2(n_879),
.B(n_919),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_SL g1093 ( 
.A(n_948),
.B(n_439),
.C(n_398),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_877),
.B(n_519),
.Y(n_1094)
);

INVx5_ASAP7_75t_L g1095 ( 
.A(n_955),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_955),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_860),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_887),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_919),
.B(n_808),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_961),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_958),
.B(n_886),
.Y(n_1101)
);

INVxp67_ASAP7_75t_SL g1102 ( 
.A(n_985),
.Y(n_1102)
);

AND2x2_ASAP7_75t_SL g1103 ( 
.A(n_963),
.B(n_307),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_899),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_950),
.B(n_938),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_901),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_836),
.B(n_842),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_830),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_950),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_952),
.B(n_808),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_952),
.B(n_751),
.Y(n_1111)
);

O2A1O1Ixp5_ASAP7_75t_L g1112 ( 
.A1(n_875),
.A2(n_748),
.B(n_702),
.C(n_706),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_961),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_918),
.B(n_683),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_882),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_904),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_833),
.Y(n_1117)
);

NAND2x1p5_ASAP7_75t_L g1118 ( 
.A(n_985),
.B(n_687),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_994),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_985),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_883),
.Y(n_1121)
);

INVx4_ASAP7_75t_L g1122 ( 
.A(n_985),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_907),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_918),
.B(n_683),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_852),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_866),
.A2(n_821),
.B1(n_823),
.B2(n_817),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_958),
.B(n_520),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_913),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_925),
.B(n_683),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_890),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_908),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_925),
.B(n_725),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_911),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_866),
.B(n_521),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_844),
.B(n_396),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_929),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_917),
.A2(n_730),
.B(n_687),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_858),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_914),
.Y(n_1139)
);

AND2x2_ASAP7_75t_SL g1140 ( 
.A(n_947),
.B(n_307),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_916),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_920),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_998),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_928),
.B(n_725),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_928),
.B(n_725),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_924),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_934),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_849),
.A2(n_307),
.B1(n_731),
.B2(n_739),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_946),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_973),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_949),
.B(n_725),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_894),
.B(n_524),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_850),
.A2(n_823),
.B1(n_817),
.B2(n_727),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_984),
.Y(n_1154)
);

NOR2x1p5_ASAP7_75t_L g1155 ( 
.A(n_903),
.B(n_976),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_859),
.Y(n_1156)
);

NAND2x1p5_ASAP7_75t_L g1157 ( 
.A(n_959),
.B(n_687),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_892),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_992),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_R g1160 ( 
.A(n_846),
.B(n_269),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_952),
.B(n_751),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_917),
.A2(n_527),
.B(n_529),
.C(n_531),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_935),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_983),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_995),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_983),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_878),
.B(n_526),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_940),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_949),
.B(n_727),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_944),
.A2(n_888),
.B1(n_894),
.B2(n_952),
.Y(n_1170)
);

INVx8_ASAP7_75t_L g1171 ( 
.A(n_895),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_986),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_863),
.Y(n_1173)
);

OR2x4_ASAP7_75t_L g1174 ( 
.A(n_888),
.B(n_401),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_966),
.B(n_727),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_988),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_966),
.B(n_727),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_896),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_931),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_989),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_952),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_952),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_960),
.B(n_407),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_970),
.B(n_741),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_970),
.B(n_741),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_991),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_969),
.B(n_741),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1025),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1182),
.A2(n_953),
.B(n_912),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1054),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1049),
.B(n_1024),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_L g1192 ( 
.A(n_1044),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1012),
.B(n_922),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1172),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1182),
.A2(n_975),
.B(n_926),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1099),
.A2(n_730),
.B(n_687),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_SL g1197 ( 
.A1(n_1063),
.A2(n_873),
.B(n_865),
.C(n_897),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1033),
.B(n_870),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1058),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1081),
.B(n_945),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1025),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1001),
.B(n_941),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_SL g1203 ( 
.A(n_1032),
.Y(n_1203)
);

O2A1O1Ixp5_ASAP7_75t_L g1204 ( 
.A1(n_1137),
.A2(n_889),
.B(n_979),
.C(n_997),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1099),
.A2(n_806),
.B(n_730),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1103),
.A2(n_981),
.B1(n_993),
.B2(n_987),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1001),
.B(n_996),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1059),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1025),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1011),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1081),
.B(n_962),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1107),
.B(n_951),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1021),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1070),
.B(n_957),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1110),
.A2(n_806),
.B(n_730),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1018),
.B(n_968),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1028),
.A2(n_990),
.B1(n_446),
.B2(n_444),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1046),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1063),
.B(n_741),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1037),
.Y(n_1220)
);

CKINVDCx16_ASAP7_75t_R g1221 ( 
.A(n_1021),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1035),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1028),
.B(n_271),
.Y(n_1223)
);

OR2x2_ASAP7_75t_SL g1224 ( 
.A(n_1093),
.B(n_1053),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1008),
.B(n_749),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1070),
.A2(n_729),
.B(n_702),
.C(n_706),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1000),
.B(n_541),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1103),
.A2(n_379),
.B1(n_322),
.B2(n_334),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1086),
.A2(n_731),
.B(n_710),
.C(n_713),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1110),
.A2(n_806),
.B(n_754),
.Y(n_1230)
);

NAND2xp33_ASAP7_75t_SL g1231 ( 
.A(n_1155),
.B(n_1179),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1026),
.A2(n_548),
.B(n_541),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1105),
.B(n_272),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1138),
.B(n_823),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_1037),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1043),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1075),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1138),
.B(n_1134),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1052),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1044),
.B(n_806),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1092),
.A2(n_754),
.B(n_751),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1080),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1105),
.B(n_272),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1068),
.A2(n_775),
.B(n_754),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_R g1245 ( 
.A(n_1178),
.B(n_341),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1091),
.B(n_341),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1039),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1043),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1140),
.A2(n_749),
.B(n_817),
.C(n_768),
.Y(n_1249)
);

AO21x1_ASAP7_75t_L g1250 ( 
.A1(n_1114),
.A2(n_713),
.B(n_710),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1035),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1014),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1119),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1152),
.B(n_823),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1086),
.A2(n_746),
.B(n_752),
.C(n_744),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1039),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1158),
.B(n_749),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1019),
.Y(n_1258)
);

INVx3_ASAP7_75t_SL g1259 ( 
.A(n_1076),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1022),
.B(n_749),
.Y(n_1260)
);

BUFx4f_ASAP7_75t_L g1261 ( 
.A(n_1044),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1000),
.A2(n_1140),
.B1(n_1170),
.B2(n_1117),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1109),
.B(n_408),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1047),
.A2(n_742),
.B(n_739),
.Y(n_1264)
);

NOR3xp33_ASAP7_75t_L g1265 ( 
.A(n_1026),
.B(n_420),
.C(n_416),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1088),
.A2(n_822),
.B(n_814),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1100),
.B(n_408),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1115),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_1014),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1158),
.B(n_768),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1077),
.B(n_768),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1100),
.B(n_411),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1127),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1113),
.B(n_413),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1156),
.B(n_768),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1088),
.A2(n_814),
.B(n_754),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1156),
.B(n_782),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1036),
.B(n_782),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1127),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1101),
.B(n_548),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1040),
.B(n_782),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1043),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1170),
.A2(n_782),
.B(n_817),
.C(n_413),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1113),
.B(n_415),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1023),
.B(n_718),
.Y(n_1285)
);

OAI22x1_ASAP7_75t_L g1286 ( 
.A1(n_1135),
.A2(n_415),
.B1(n_444),
.B2(n_442),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1045),
.B(n_718),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1101),
.B(n_81),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1056),
.B(n_724),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1162),
.A2(n_732),
.B(n_746),
.C(n_744),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1135),
.B(n_416),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1121),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_R g1293 ( 
.A(n_1042),
.B(n_420),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_999),
.B(n_423),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1148),
.A2(n_423),
.B1(n_428),
.B2(n_441),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1183),
.B(n_428),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1035),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1183),
.A2(n_441),
.B(n_442),
.C(n_446),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1088),
.A2(n_814),
.B(n_775),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1108),
.A2(n_392),
.B1(n_343),
.B2(n_350),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1176),
.B(n_726),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1187),
.A2(n_394),
.B(n_353),
.C(n_354),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1029),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1088),
.A2(n_814),
.B(n_775),
.Y(n_1304)
);

INVxp67_ASAP7_75t_L g1305 ( 
.A(n_1065),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1148),
.A2(n_395),
.B1(n_355),
.B2(n_356),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1174),
.B(n_338),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_999),
.B(n_1003),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1162),
.A2(n_729),
.B(n_742),
.C(n_734),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1065),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1035),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1187),
.A2(n_357),
.B(n_362),
.C(n_364),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1066),
.B(n_371),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1095),
.A2(n_814),
.B(n_775),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1066),
.B(n_85),
.Y(n_1315)
);

NOR3xp33_ASAP7_75t_L g1316 ( 
.A(n_1143),
.B(n_372),
.C(n_373),
.Y(n_1316)
);

BUFx8_ASAP7_75t_L g1317 ( 
.A(n_1048),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1003),
.B(n_374),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1043),
.B(n_376),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1095),
.A2(n_822),
.B(n_775),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1098),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1041),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1004),
.B(n_732),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_SL g1324 ( 
.A1(n_1072),
.A2(n_734),
.B(n_752),
.C(n_640),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1130),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1098),
.B(n_378),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1180),
.B(n_380),
.Y(n_1327)
);

NAND3xp33_ASAP7_75t_SL g1328 ( 
.A(n_1160),
.B(n_384),
.C(n_382),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1186),
.B(n_754),
.Y(n_1329)
);

INVx5_ASAP7_75t_L g1330 ( 
.A(n_1071),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1027),
.B(n_0),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1095),
.A2(n_822),
.B(n_813),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1166),
.B(n_1),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1166),
.B(n_1160),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1164),
.B(n_822),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1030),
.Y(n_1336)
);

INVx5_ASAP7_75t_L g1337 ( 
.A(n_1071),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1015),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1072),
.A2(n_822),
.B1(n_642),
.B2(n_640),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1079),
.A2(n_642),
.B1(n_640),
.B2(n_639),
.Y(n_1340)
);

INVx8_ASAP7_75t_L g1341 ( 
.A(n_1095),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1078),
.A2(n_813),
.B(n_779),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1174),
.B(n_1),
.Y(n_1343)
);

INVx4_ASAP7_75t_L g1344 ( 
.A(n_1071),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1104),
.B(n_639),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1164),
.B(n_88),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1218),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_SL g1348 ( 
.A(n_1221),
.B(n_1048),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1238),
.B(n_1171),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1241),
.A2(n_1112),
.B(n_1064),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1250),
.A2(n_1005),
.B(n_1112),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1291),
.B(n_1090),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1202),
.B(n_1296),
.Y(n_1353)
);

OR2x6_ASAP7_75t_L g1354 ( 
.A(n_1341),
.B(n_1288),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1283),
.A2(n_1129),
.B(n_1124),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1195),
.A2(n_1020),
.B(n_1047),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1265),
.A2(n_1079),
.B(n_1167),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1192),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1191),
.B(n_1171),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1264),
.A2(n_1205),
.B(n_1196),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1189),
.A2(n_1230),
.B(n_1215),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1220),
.B(n_1171),
.Y(n_1362)
);

AOI211x1_ASAP7_75t_L g1363 ( 
.A1(n_1223),
.A2(n_1087),
.B(n_1060),
.C(n_1061),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1244),
.A2(n_1020),
.B(n_1073),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1220),
.B(n_1256),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1190),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1274),
.B(n_1200),
.Y(n_1367)
);

BUFx8_ASAP7_75t_SL g1368 ( 
.A(n_1252),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1249),
.A2(n_1050),
.A3(n_1144),
.B(n_1132),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1219),
.A2(n_1151),
.B(n_1145),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1254),
.A2(n_1078),
.B(n_1085),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1288),
.B(n_1082),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1247),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1231),
.A2(n_1167),
.B1(n_1083),
.B2(n_1125),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1213),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1199),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1214),
.B(n_1106),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1192),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1207),
.A2(n_1074),
.B(n_1169),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_L g1380 ( 
.A(n_1330),
.B(n_1030),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1246),
.B(n_1082),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1198),
.A2(n_1185),
.B(n_1177),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1256),
.Y(n_1383)
);

NAND2x1_ASAP7_75t_L g1384 ( 
.A(n_1236),
.B(n_1096),
.Y(n_1384)
);

AOI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1225),
.A2(n_1184),
.B(n_1175),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1346),
.A2(n_1007),
.B(n_1102),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1260),
.A2(n_1078),
.B(n_1007),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1339),
.A2(n_1073),
.B(n_1111),
.Y(n_1388)
);

NAND3x1_ASAP7_75t_L g1389 ( 
.A(n_1343),
.B(n_1084),
.C(n_1016),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1339),
.A2(n_1340),
.B(n_1309),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1233),
.B(n_1116),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1206),
.A2(n_1083),
.B(n_1038),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1212),
.A2(n_1078),
.B(n_1157),
.Y(n_1393)
);

NOR2xp67_ASAP7_75t_SL g1394 ( 
.A(n_1194),
.B(n_1071),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1340),
.A2(n_1142),
.A3(n_1123),
.B(n_1168),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1290),
.A2(n_1111),
.B(n_1161),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1243),
.B(n_1128),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1308),
.B(n_1041),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1210),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1208),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1322),
.B(n_1139),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1258),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1341),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1204),
.A2(n_1161),
.B(n_1051),
.Y(n_1404)
);

O2A1O1Ixp5_ASAP7_75t_SL g1405 ( 
.A1(n_1211),
.A2(n_1017),
.B(n_1069),
.C(n_1057),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1268),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1273),
.B(n_1279),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1239),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1327),
.B(n_1141),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1266),
.A2(n_1299),
.B(n_1276),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1263),
.Y(n_1411)
);

BUFx2_ASAP7_75t_R g1412 ( 
.A(n_1269),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1237),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1259),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1197),
.A2(n_1009),
.B(n_1094),
.C(n_1067),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1236),
.A2(n_1157),
.B(n_1102),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1206),
.A2(n_1146),
.B(n_1147),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1303),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1262),
.A2(n_1163),
.B(n_1034),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1338),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1257),
.A2(n_1062),
.B(n_1126),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1304),
.A2(n_1051),
.B(n_1057),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1216),
.B(n_1173),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1261),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1248),
.A2(n_1118),
.B(n_1282),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1257),
.A2(n_1013),
.B(n_1010),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1270),
.A2(n_1006),
.B(n_1002),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1245),
.B(n_1173),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1334),
.B(n_1173),
.Y(n_1429)
);

NAND2x1p5_ASAP7_75t_L g1430 ( 
.A(n_1261),
.B(n_1096),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1248),
.A2(n_1118),
.B(n_1181),
.Y(n_1431)
);

AOI221x1_ASAP7_75t_L g1432 ( 
.A1(n_1286),
.A2(n_1298),
.B1(n_1295),
.B2(n_1306),
.C(n_1307),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1270),
.A2(n_1136),
.B(n_1165),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1302),
.A2(n_1149),
.A3(n_1130),
.B(n_1154),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1235),
.B(n_1032),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1341),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1228),
.A2(n_1150),
.B1(n_1069),
.B2(n_1173),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1193),
.A2(n_1016),
.B1(n_1032),
.B2(n_1031),
.Y(n_1438)
);

AOI221xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1217),
.A2(n_1159),
.B1(n_1097),
.B2(n_1055),
.C(n_1089),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1282),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1324),
.A2(n_1153),
.B(n_1154),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1321),
.B(n_1280),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1229),
.A2(n_1149),
.B(n_1133),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1314),
.A2(n_1133),
.B(n_1131),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1326),
.B(n_1131),
.Y(n_1445)
);

AO31x2_ASAP7_75t_L g1446 ( 
.A1(n_1312),
.A2(n_1122),
.A3(n_1038),
.B(n_642),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1285),
.A2(n_1122),
.B(n_1120),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1285),
.A2(n_1120),
.B(n_1150),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1329),
.A2(n_1150),
.A3(n_1120),
.B(n_5),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1305),
.A2(n_1150),
.B1(n_1120),
.B2(n_813),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1330),
.A2(n_813),
.B1(n_779),
.B2(n_643),
.Y(n_1451)
);

AOI31xp67_ASAP7_75t_L g1452 ( 
.A1(n_1292),
.A2(n_813),
.A3(n_779),
.B(n_158),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1294),
.B(n_2),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1255),
.A2(n_813),
.B(n_779),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1333),
.B(n_2),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1267),
.B(n_4),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1336),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1280),
.B(n_6),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1325),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1188),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1242),
.Y(n_1461)
);

NOR4xp25_ASAP7_75t_L g1462 ( 
.A(n_1232),
.B(n_6),
.C(n_8),
.D(n_12),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1287),
.A2(n_779),
.B(n_643),
.Y(n_1463)
);

O2A1O1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1272),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1316),
.A2(n_643),
.B(n_16),
.C(n_17),
.Y(n_1465)
);

OR2x6_ASAP7_75t_L g1466 ( 
.A(n_1346),
.B(n_643),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1310),
.B(n_146),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1289),
.A2(n_779),
.B(n_615),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1188),
.Y(n_1469)
);

NAND3x1_ASAP7_75t_L g1470 ( 
.A(n_1331),
.B(n_13),
.C(n_18),
.Y(n_1470)
);

OAI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1232),
.A2(n_1295),
.B(n_1306),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1320),
.A2(n_152),
.B(n_226),
.Y(n_1472)
);

AO31x2_ASAP7_75t_L g1473 ( 
.A1(n_1278),
.A2(n_19),
.A3(n_20),
.B(n_22),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1227),
.B(n_20),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1227),
.B(n_25),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1336),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1281),
.A2(n_615),
.B(n_223),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1313),
.B(n_25),
.Y(n_1478)
);

AO31x2_ASAP7_75t_L g1479 ( 
.A1(n_1345),
.A2(n_26),
.A3(n_27),
.B(n_31),
.Y(n_1479)
);

BUFx10_ASAP7_75t_L g1480 ( 
.A(n_1315),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1226),
.A2(n_137),
.B(n_212),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1277),
.B(n_32),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1277),
.B(n_32),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1301),
.Y(n_1484)
);

AND2x6_ASAP7_75t_L g1485 ( 
.A(n_1315),
.B(n_193),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1301),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1323),
.A2(n_615),
.B(n_185),
.Y(n_1487)
);

AOI221x1_ASAP7_75t_L g1488 ( 
.A1(n_1328),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.C(n_42),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1253),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1188),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1284),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1317),
.Y(n_1492)
);

INVx4_ASAP7_75t_SL g1493 ( 
.A(n_1251),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1332),
.A2(n_130),
.B(n_179),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1330),
.A2(n_615),
.B(n_170),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1271),
.A2(n_103),
.B(n_168),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1271),
.A2(n_144),
.B(n_135),
.Y(n_1497)
);

OAI22x1_ASAP7_75t_L g1498 ( 
.A1(n_1318),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1330),
.A2(n_615),
.B(n_102),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1300),
.B(n_615),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1317),
.Y(n_1501)
);

AO31x2_ASAP7_75t_L g1502 ( 
.A1(n_1234),
.A2(n_45),
.A3(n_46),
.B(n_47),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1275),
.B(n_1319),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1335),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1342),
.A2(n_95),
.B(n_93),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1201),
.B(n_48),
.Y(n_1506)
);

BUFx12f_ASAP7_75t_L g1507 ( 
.A(n_1224),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1251),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1203),
.A2(n_49),
.B(n_50),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1201),
.A2(n_50),
.B(n_58),
.C(n_61),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1209),
.B(n_63),
.Y(n_1511)
);

INVx3_ASAP7_75t_SL g1512 ( 
.A(n_1240),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1222),
.A2(n_91),
.B(n_64),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1293),
.B(n_63),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1240),
.A2(n_65),
.B(n_67),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1222),
.B(n_74),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1297),
.B(n_74),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1251),
.B(n_1311),
.C(n_1297),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1240),
.A2(n_67),
.B(n_69),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1337),
.A2(n_70),
.B(n_73),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1360),
.A2(n_1337),
.B(n_1344),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1375),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1354),
.B(n_1311),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1350),
.A2(n_1337),
.B(n_1311),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1367),
.A2(n_1353),
.B(n_1397),
.C(n_1391),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_R g1526 ( 
.A1(n_1372),
.A2(n_70),
.B(n_1337),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1386),
.B(n_1344),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1361),
.A2(n_1356),
.B(n_1410),
.Y(n_1528)
);

CKINVDCx16_ASAP7_75t_R g1529 ( 
.A(n_1492),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1354),
.B(n_1398),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1439),
.A2(n_1355),
.B(n_1390),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1365),
.B(n_1383),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1455),
.B(n_1407),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1409),
.A2(n_1432),
.B(n_1417),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1376),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1471),
.A2(n_1513),
.B(n_1357),
.C(n_1456),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1411),
.A2(n_1381),
.B1(n_1377),
.B2(n_1352),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1478),
.B(n_1372),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1364),
.A2(n_1422),
.B(n_1404),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1373),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1396),
.A2(n_1388),
.B(n_1481),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1383),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1402),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1444),
.A2(n_1494),
.B(n_1472),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1423),
.B(n_1429),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1505),
.A2(n_1385),
.B(n_1496),
.Y(n_1546)
);

AO31x2_ASAP7_75t_L g1547 ( 
.A1(n_1488),
.A2(n_1371),
.A3(n_1448),
.B(n_1387),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1418),
.Y(n_1548)
);

BUFx2_ASAP7_75t_SL g1549 ( 
.A(n_1358),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1408),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1442),
.B(n_1445),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1420),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1393),
.A2(n_1405),
.B(n_1370),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1382),
.A2(n_1463),
.B(n_1355),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1401),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1395),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1453),
.A2(n_1491),
.B1(n_1428),
.B2(n_1471),
.Y(n_1557)
);

AOI21xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1509),
.A2(n_1413),
.B(n_1498),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1443),
.A2(n_1477),
.B(n_1416),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1504),
.A2(n_1513),
.B1(n_1485),
.B2(n_1379),
.Y(n_1560)
);

AO31x2_ASAP7_75t_L g1561 ( 
.A1(n_1437),
.A2(n_1465),
.A3(n_1447),
.B(n_1486),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1439),
.A2(n_1392),
.B(n_1419),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1354),
.B(n_1398),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1431),
.A2(n_1415),
.B(n_1421),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_SL g1565 ( 
.A1(n_1392),
.A2(n_1482),
.B(n_1483),
.Y(n_1565)
);

AND2x6_ASAP7_75t_L g1566 ( 
.A(n_1484),
.B(n_1374),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1426),
.A2(n_1487),
.B(n_1427),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1399),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1433),
.A2(n_1425),
.B(n_1468),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1514),
.B(n_1349),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1359),
.B(n_1503),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1504),
.A2(n_1485),
.B1(n_1520),
.B2(n_1507),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1362),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1460),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1357),
.A2(n_1500),
.B(n_1374),
.Y(n_1575)
);

XOR2xp5_ASAP7_75t_L g1576 ( 
.A(n_1400),
.B(n_1412),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1358),
.Y(n_1577)
);

NAND2xp33_ASAP7_75t_R g1578 ( 
.A(n_1351),
.B(n_1440),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1459),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1406),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1511),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1506),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1474),
.B(n_1475),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1485),
.A2(n_1458),
.B1(n_1438),
.B2(n_1435),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1438),
.A2(n_1462),
.B1(n_1517),
.B2(n_1516),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1454),
.A2(n_1351),
.B(n_1519),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1434),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1495),
.A2(n_1499),
.B(n_1497),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1466),
.A2(n_1441),
.B(n_1497),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1450),
.A2(n_1384),
.B(n_1451),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1358),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1457),
.A2(n_1476),
.B(n_1440),
.Y(n_1592)
);

INVx8_ASAP7_75t_L g1593 ( 
.A(n_1469),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1378),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1403),
.A2(n_1436),
.B(n_1518),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_SL g1596 ( 
.A1(n_1464),
.A2(n_1509),
.B(n_1501),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1480),
.B(n_1424),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1378),
.Y(n_1598)
);

OAI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1403),
.A2(n_1436),
.B(n_1518),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1449),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1348),
.B(n_1467),
.Y(n_1601)
);

BUFx2_ASAP7_75t_R g1602 ( 
.A(n_1368),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1449),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1466),
.A2(n_1441),
.B(n_1380),
.Y(n_1604)
);

AOI21xp33_ASAP7_75t_L g1605 ( 
.A1(n_1510),
.A2(n_1470),
.B(n_1466),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1489),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1462),
.A2(n_1467),
.B1(n_1512),
.B2(n_1414),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1449),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1434),
.Y(n_1609)
);

BUFx2_ASAP7_75t_R g1610 ( 
.A(n_1490),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1508),
.B(n_1490),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1378),
.Y(n_1612)
);

OA21x2_ASAP7_75t_L g1613 ( 
.A1(n_1452),
.A2(n_1363),
.B(n_1395),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1363),
.B(n_1424),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1389),
.A2(n_1515),
.B(n_1430),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1508),
.B(n_1469),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1369),
.A2(n_1395),
.B(n_1434),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1424),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1369),
.Y(n_1619)
);

OR2x6_ASAP7_75t_L g1620 ( 
.A(n_1469),
.B(n_1493),
.Y(n_1620)
);

AO31x2_ASAP7_75t_L g1621 ( 
.A1(n_1446),
.A2(n_1369),
.A3(n_1473),
.B(n_1479),
.Y(n_1621)
);

OA21x2_ASAP7_75t_L g1622 ( 
.A1(n_1446),
.A2(n_1479),
.B(n_1473),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1446),
.A2(n_1493),
.B(n_1473),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1502),
.B(n_1461),
.Y(n_1624)
);

OAI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1502),
.A2(n_851),
.B1(n_1367),
.B2(n_847),
.C(n_708),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1383),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1629)
);

CKINVDCx6p67_ASAP7_75t_R g1630 ( 
.A(n_1414),
.Y(n_1630)
);

OAI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1367),
.A2(n_851),
.B1(n_847),
.B2(n_708),
.C(n_1296),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1455),
.B(n_1191),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1408),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1350),
.A2(n_1439),
.B(n_1355),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1408),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1386),
.A2(n_1103),
.B(n_1099),
.Y(n_1639)
);

OA21x2_ASAP7_75t_L g1640 ( 
.A1(n_1350),
.A2(n_1439),
.B(n_1355),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1367),
.A2(n_1291),
.B1(n_1296),
.B2(n_851),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_SL g1642 ( 
.A(n_1367),
.B(n_851),
.C(n_1296),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1347),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1358),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1366),
.Y(n_1645)
);

NAND2x1p5_ASAP7_75t_L g1646 ( 
.A(n_1394),
.B(n_1043),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1647)
);

OA21x2_ASAP7_75t_L g1648 ( 
.A1(n_1350),
.A2(n_1439),
.B(n_1355),
.Y(n_1648)
);

OAI21x1_ASAP7_75t_L g1649 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1367),
.A2(n_1103),
.B(n_851),
.C(n_1140),
.Y(n_1650)
);

AO21x1_ASAP7_75t_L g1651 ( 
.A1(n_1367),
.A2(n_851),
.B(n_1296),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1347),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1408),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1367),
.A2(n_1028),
.B1(n_847),
.B2(n_1291),
.Y(n_1654)
);

AOI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1367),
.A2(n_847),
.B1(n_1028),
.B2(n_849),
.C(n_851),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1347),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_SL g1657 ( 
.A1(n_1513),
.A2(n_1392),
.B(n_1417),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1366),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1347),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1661)
);

CKINVDCx6p67_ASAP7_75t_R g1662 ( 
.A(n_1414),
.Y(n_1662)
);

AO31x2_ASAP7_75t_L g1663 ( 
.A1(n_1432),
.A2(n_1137),
.A3(n_1250),
.B(n_1005),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1358),
.Y(n_1664)
);

NOR2x1_ASAP7_75t_SL g1665 ( 
.A(n_1437),
.B(n_1330),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1666)
);

A2O1A1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1367),
.A2(n_1103),
.B(n_851),
.C(n_1140),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1367),
.A2(n_851),
.B(n_1291),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1353),
.B(n_847),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1358),
.Y(n_1670)
);

O2A1O1Ixp33_ASAP7_75t_SL g1671 ( 
.A1(n_1513),
.A2(n_1028),
.B(n_1197),
.C(n_1465),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1367),
.B(n_851),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1386),
.A2(n_1103),
.B(n_1099),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1386),
.A2(n_1103),
.B(n_1099),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1386),
.A2(n_1103),
.B(n_1099),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1347),
.Y(n_1676)
);

AOI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1370),
.A2(n_1385),
.B(n_1382),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1347),
.Y(n_1678)
);

CKINVDCx20_ASAP7_75t_R g1679 ( 
.A(n_1368),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1365),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1347),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1383),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1367),
.A2(n_1291),
.B1(n_1296),
.B2(n_851),
.Y(n_1683)
);

CKINVDCx8_ASAP7_75t_R g1684 ( 
.A(n_1413),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1353),
.B(n_847),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1350),
.A2(n_1439),
.B(n_1355),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1347),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1688)
);

AO31x2_ASAP7_75t_L g1689 ( 
.A1(n_1432),
.A2(n_1137),
.A3(n_1250),
.B(n_1005),
.Y(n_1689)
);

OAI21x1_ASAP7_75t_L g1690 ( 
.A1(n_1360),
.A2(n_1350),
.B(n_1361),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1354),
.B(n_1398),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1358),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1367),
.A2(n_851),
.B(n_1291),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1368),
.Y(n_1694)
);

OA21x2_ASAP7_75t_L g1695 ( 
.A1(n_1350),
.A2(n_1439),
.B(n_1355),
.Y(n_1695)
);

OAI21x1_ASAP7_75t_L g1696 ( 
.A1(n_1350),
.A2(n_1360),
.B(n_1361),
.Y(n_1696)
);

AOI221x1_ASAP7_75t_SL g1697 ( 
.A1(n_1672),
.A2(n_1537),
.B1(n_1685),
.B2(n_1669),
.C(n_1583),
.Y(n_1697)
);

OA21x2_ASAP7_75t_L g1698 ( 
.A1(n_1589),
.A2(n_1617),
.B(n_1553),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1641),
.A2(n_1683),
.B(n_1693),
.C(n_1668),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_1679),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1532),
.B(n_1680),
.Y(n_1701)
);

AOI221x1_ASAP7_75t_SL g1702 ( 
.A1(n_1672),
.A2(n_1583),
.B1(n_1605),
.B2(n_1582),
.C(n_1571),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1591),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1555),
.B(n_1525),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1650),
.A2(n_1667),
.B(n_1536),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1680),
.B(n_1581),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1650),
.A2(n_1667),
.B(n_1639),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1627),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1535),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1627),
.Y(n_1710)
);

AOI21x1_ASAP7_75t_SL g1711 ( 
.A1(n_1526),
.A2(n_1601),
.B(n_1556),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1555),
.B(n_1525),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1631),
.A2(n_1642),
.B(n_1625),
.C(n_1536),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1534),
.B(n_1655),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1654),
.B(n_1566),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1654),
.B(n_1566),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1560),
.A2(n_1607),
.B1(n_1557),
.B2(n_1572),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1560),
.A2(n_1607),
.B1(n_1572),
.B2(n_1675),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1639),
.A2(n_1674),
.B(n_1673),
.Y(n_1719)
);

AOI21x1_ASAP7_75t_SL g1720 ( 
.A1(n_1556),
.A2(n_1570),
.B(n_1523),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1573),
.Y(n_1721)
);

INVx3_ASAP7_75t_SL g1722 ( 
.A(n_1694),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1673),
.A2(n_1675),
.B(n_1674),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1545),
.B(n_1551),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1566),
.B(n_1651),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1533),
.B(n_1632),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1566),
.B(n_1585),
.Y(n_1727)
);

O2A1O1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1642),
.A2(n_1671),
.B(n_1558),
.C(n_1596),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1573),
.B(n_1542),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1671),
.A2(n_1564),
.B(n_1559),
.Y(n_1730)
);

O2A1O1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1565),
.A2(n_1657),
.B(n_1624),
.C(n_1575),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1538),
.B(n_1530),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1530),
.B(n_1563),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1574),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1585),
.A2(n_1584),
.B1(n_1610),
.B2(n_1540),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1584),
.A2(n_1540),
.B1(n_1682),
.B2(n_1645),
.Y(n_1736)
);

INVxp67_ASAP7_75t_L g1737 ( 
.A(n_1568),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1527),
.A2(n_1567),
.B(n_1665),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1566),
.B(n_1543),
.Y(n_1739)
);

OAI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1615),
.A2(n_1548),
.B(n_1658),
.C(n_1552),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_1694),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1550),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1527),
.A2(n_1604),
.B(n_1569),
.Y(n_1743)
);

AOI21x1_ASAP7_75t_SL g1744 ( 
.A1(n_1691),
.A2(n_1578),
.B(n_1623),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1633),
.B(n_1638),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1579),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1653),
.B(n_1550),
.Y(n_1747)
);

BUFx10_ASAP7_75t_L g1748 ( 
.A(n_1597),
.Y(n_1748)
);

O2A1O1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1597),
.A2(n_1522),
.B(n_1618),
.C(n_1664),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1611),
.B(n_1643),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1562),
.A2(n_1580),
.B1(n_1646),
.B2(n_1620),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1562),
.B(n_1652),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1577),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1656),
.B(n_1660),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1620),
.A2(n_1576),
.B(n_1577),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1593),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1562),
.B(n_1656),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1660),
.B(n_1676),
.Y(n_1758)
);

A2O1A1Ixp33_ASAP7_75t_L g1759 ( 
.A1(n_1588),
.A2(n_1604),
.B(n_1586),
.C(n_1554),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1616),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_SL g1761 ( 
.A1(n_1620),
.A2(n_1670),
.B(n_1594),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1684),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1679),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1591),
.A2(n_1594),
.B(n_1670),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1528),
.A2(n_1531),
.B(n_1546),
.Y(n_1765)
);

O2A1O1Ixp5_ASAP7_75t_L g1766 ( 
.A1(n_1619),
.A2(n_1677),
.B(n_1603),
.C(n_1600),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1676),
.B(n_1687),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1678),
.B(n_1687),
.Y(n_1768)
);

OA22x2_ASAP7_75t_L g1769 ( 
.A1(n_1608),
.A2(n_1606),
.B1(n_1692),
.B2(n_1618),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1678),
.B(n_1681),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1598),
.B(n_1644),
.Y(n_1771)
);

OA21x2_ASAP7_75t_L g1772 ( 
.A1(n_1696),
.A2(n_1541),
.B(n_1690),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1529),
.A2(n_1644),
.B1(n_1664),
.B2(n_1598),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1561),
.B(n_1621),
.Y(n_1774)
);

AOI21x1_ASAP7_75t_SL g1775 ( 
.A1(n_1547),
.A2(n_1602),
.B(n_1662),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1561),
.B(n_1621),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1612),
.B(n_1591),
.Y(n_1777)
);

OA21x2_ASAP7_75t_L g1778 ( 
.A1(n_1696),
.A2(n_1628),
.B(n_1688),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1531),
.A2(n_1626),
.B(n_1629),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1634),
.A2(n_1636),
.B(n_1666),
.Y(n_1780)
);

OA21x2_ASAP7_75t_L g1781 ( 
.A1(n_1637),
.A2(n_1649),
.B(n_1661),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1622),
.Y(n_1782)
);

O2A1O1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1612),
.A2(n_1609),
.B(n_1587),
.C(n_1531),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1622),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1594),
.B(n_1670),
.Y(n_1785)
);

NAND2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1595),
.B(n_1599),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1590),
.A2(n_1544),
.B(n_1592),
.C(n_1539),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1594),
.B(n_1670),
.Y(n_1788)
);

NOR2xp67_ASAP7_75t_L g1789 ( 
.A(n_1549),
.B(n_1630),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1521),
.B(n_1621),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1613),
.A2(n_1593),
.B1(n_1686),
.B2(n_1695),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1663),
.B(n_1689),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1663),
.B(n_1689),
.Y(n_1793)
);

OA22x2_ASAP7_75t_L g1794 ( 
.A1(n_1647),
.A2(n_1659),
.B1(n_1613),
.B2(n_1524),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1524),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1635),
.B(n_1640),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1635),
.B(n_1640),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1640),
.B(n_1648),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1648),
.B(n_1686),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1695),
.A2(n_1648),
.B(n_1686),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1695),
.Y(n_1801)
);

AOI21x1_ASAP7_75t_SL g1802 ( 
.A1(n_1614),
.A2(n_851),
.B(n_1353),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1650),
.A2(n_1103),
.B1(n_1667),
.B2(n_1654),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1627),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1650),
.A2(n_1103),
.B1(n_1667),
.B2(n_1654),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1530),
.B(n_1563),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1650),
.A2(n_1103),
.B1(n_1667),
.B2(n_1654),
.Y(n_1807)
);

OA21x2_ASAP7_75t_L g1808 ( 
.A1(n_1589),
.A2(n_1617),
.B(n_1553),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1533),
.B(n_1545),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1533),
.B(n_1545),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1650),
.A2(n_1103),
.B1(n_1667),
.B2(n_1654),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1550),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_SL g1813 ( 
.A(n_1602),
.B(n_1412),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1641),
.B(n_691),
.Y(n_1814)
);

OAI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1650),
.A2(n_1103),
.B1(n_1667),
.B2(n_1654),
.Y(n_1815)
);

AOI21x1_ASAP7_75t_SL g1816 ( 
.A1(n_1614),
.A2(n_851),
.B(n_1353),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1533),
.B(n_1545),
.Y(n_1817)
);

AND2x4_ASAP7_75t_SL g1818 ( 
.A(n_1679),
.B(n_678),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1533),
.B(n_1545),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1532),
.B(n_1680),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1650),
.A2(n_1103),
.B(n_1667),
.Y(n_1821)
);

AOI221x1_ASAP7_75t_SL g1822 ( 
.A1(n_1672),
.A2(n_849),
.B1(n_1028),
.B2(n_853),
.C(n_862),
.Y(n_1822)
);

OA21x2_ASAP7_75t_L g1823 ( 
.A1(n_1589),
.A2(n_1617),
.B(n_1553),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_SL g1824 ( 
.A1(n_1650),
.A2(n_1667),
.B(n_693),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1550),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1555),
.B(n_1525),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_SL g1827 ( 
.A(n_1602),
.B(n_1412),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1627),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1525),
.B(n_1672),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1650),
.A2(n_1103),
.B(n_1667),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1650),
.A2(n_1103),
.B1(n_1667),
.B2(n_1654),
.Y(n_1831)
);

OR2x6_ASAP7_75t_L g1832 ( 
.A(n_1657),
.B(n_1575),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1523),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1650),
.A2(n_1103),
.B1(n_1667),
.B2(n_1654),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1532),
.B(n_1680),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1650),
.A2(n_1103),
.B1(n_1667),
.B2(n_1654),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1555),
.B(n_1525),
.Y(n_1837)
);

AND2x2_ASAP7_75t_SL g1838 ( 
.A(n_1560),
.B(n_1607),
.Y(n_1838)
);

O2A1O1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1631),
.A2(n_851),
.B(n_1693),
.C(n_1668),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1734),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1708),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1700),
.Y(n_1842)
);

AO21x2_ASAP7_75t_L g1843 ( 
.A1(n_1800),
.A2(n_1765),
.B(n_1779),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1792),
.B(n_1709),
.Y(n_1844)
);

INVxp33_ASAP7_75t_L g1845 ( 
.A(n_1809),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_SL g1846 ( 
.A(n_1813),
.B(n_1827),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1752),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1829),
.B(n_1701),
.Y(n_1848)
);

AND2x4_ASAP7_75t_SL g1849 ( 
.A(n_1748),
.B(n_1806),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1786),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1774),
.B(n_1776),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1752),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1739),
.B(n_1832),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1757),
.Y(n_1854)
);

AO21x2_ASAP7_75t_L g1855 ( 
.A1(n_1719),
.A2(n_1730),
.B(n_1759),
.Y(n_1855)
);

AO21x2_ASAP7_75t_L g1856 ( 
.A1(n_1743),
.A2(n_1707),
.B(n_1798),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1757),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1804),
.Y(n_1858)
);

AO21x2_ASAP7_75t_L g1859 ( 
.A1(n_1799),
.A2(n_1830),
.B(n_1821),
.Y(n_1859)
);

INVx5_ASAP7_75t_L g1860 ( 
.A(n_1832),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1739),
.B(n_1832),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1828),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1723),
.A2(n_1705),
.B(n_1839),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1786),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1746),
.Y(n_1865)
);

INVxp33_ASAP7_75t_L g1866 ( 
.A(n_1810),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1782),
.Y(n_1867)
);

AO21x2_ASAP7_75t_L g1868 ( 
.A1(n_1787),
.A2(n_1791),
.B(n_1801),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1784),
.Y(n_1869)
);

AND2x4_ASAP7_75t_SL g1870 ( 
.A(n_1748),
.B(n_1806),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1769),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1721),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1725),
.B(n_1715),
.Y(n_1873)
);

AO21x1_ASAP7_75t_SL g1874 ( 
.A1(n_1727),
.A2(n_1725),
.B(n_1712),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1715),
.B(n_1716),
.Y(n_1875)
);

NAND2x1_ASAP7_75t_L g1876 ( 
.A(n_1824),
.B(n_1738),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1790),
.Y(n_1877)
);

INVxp67_ASAP7_75t_SL g1878 ( 
.A(n_1704),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1710),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1766),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1769),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1716),
.B(n_1727),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1795),
.Y(n_1883)
);

BUFx2_ASAP7_75t_L g1884 ( 
.A(n_1712),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1820),
.Y(n_1885)
);

INVx4_ASAP7_75t_L g1886 ( 
.A(n_1825),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1750),
.B(n_1817),
.Y(n_1887)
);

AOI21x1_ASAP7_75t_L g1888 ( 
.A1(n_1826),
.A2(n_1837),
.B(n_1751),
.Y(n_1888)
);

NAND3xp33_ASAP7_75t_L g1889 ( 
.A(n_1699),
.B(n_1713),
.C(n_1728),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1835),
.B(n_1724),
.Y(n_1890)
);

BUFx5_ASAP7_75t_L g1891 ( 
.A(n_1797),
.Y(n_1891)
);

AO21x2_ASAP7_75t_L g1892 ( 
.A1(n_1793),
.A2(n_1826),
.B(n_1837),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1838),
.A2(n_1717),
.B1(n_1718),
.B2(n_1735),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1760),
.B(n_1697),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1783),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1747),
.Y(n_1896)
);

AOI21x1_ASAP7_75t_L g1897 ( 
.A1(n_1751),
.A2(n_1714),
.B(n_1718),
.Y(n_1897)
);

AO21x2_ASAP7_75t_L g1898 ( 
.A1(n_1803),
.A2(n_1836),
.B(n_1805),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1819),
.B(n_1733),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1706),
.B(n_1729),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1796),
.B(n_1714),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1753),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1702),
.B(n_1822),
.Y(n_1903)
);

OA21x2_ASAP7_75t_L g1904 ( 
.A1(n_1803),
.A2(n_1836),
.B(n_1834),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1754),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1758),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1767),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1768),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1698),
.B(n_1808),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1770),
.Y(n_1910)
);

AO21x2_ASAP7_75t_L g1911 ( 
.A1(n_1805),
.A2(n_1834),
.B(n_1831),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1794),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1745),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1794),
.Y(n_1914)
);

OA21x2_ASAP7_75t_L g1915 ( 
.A1(n_1807),
.A2(n_1831),
.B(n_1815),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1736),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1833),
.B(n_1726),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1736),
.B(n_1731),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1717),
.A2(n_1735),
.B1(n_1807),
.B2(n_1815),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1823),
.Y(n_1920)
);

OAI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1889),
.A2(n_1814),
.B1(n_1811),
.B2(n_1740),
.C(n_1737),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1867),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1867),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1869),
.Y(n_1924)
);

OAI33xp33_ASAP7_75t_L g1925 ( 
.A1(n_1903),
.A2(n_1811),
.A3(n_1773),
.B1(n_1749),
.B2(n_1763),
.B3(n_1741),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1919),
.A2(n_1732),
.B1(n_1833),
.B2(n_1773),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1883),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1878),
.B(n_1742),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1884),
.B(n_1812),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1884),
.B(n_1901),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1912),
.B(n_1914),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1912),
.B(n_1914),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1891),
.B(n_1772),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1898),
.A2(n_1911),
.B1(n_1893),
.B2(n_1863),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1891),
.B(n_1778),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1847),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1873),
.B(n_1781),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1873),
.B(n_1859),
.Y(n_1938)
);

OR2x2_ASAP7_75t_L g1939 ( 
.A(n_1901),
.B(n_1780),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1859),
.B(n_1781),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1892),
.B(n_1788),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1892),
.B(n_1785),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1859),
.B(n_1777),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1844),
.B(n_1771),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1877),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1844),
.B(n_1703),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1856),
.B(n_1744),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1856),
.B(n_1764),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1847),
.B(n_1761),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1856),
.B(n_1755),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1852),
.B(n_1756),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1852),
.B(n_1722),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1849),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1854),
.B(n_1762),
.Y(n_1954)
);

NOR2xp67_ASAP7_75t_L g1955 ( 
.A(n_1854),
.B(n_1789),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_SL g1956 ( 
.A1(n_1898),
.A2(n_1818),
.B1(n_1711),
.B2(n_1775),
.Y(n_1956)
);

INVx2_ASAP7_75t_SL g1957 ( 
.A(n_1877),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1857),
.B(n_1816),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1857),
.B(n_1802),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1880),
.B(n_1720),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1880),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1876),
.Y(n_1962)
);

AOI221xp5_ASAP7_75t_L g1963 ( 
.A1(n_1921),
.A2(n_1918),
.B1(n_1894),
.B2(n_1848),
.C(n_1916),
.Y(n_1963)
);

AOI222xp33_ASAP7_75t_L g1964 ( 
.A1(n_1921),
.A2(n_1934),
.B1(n_1925),
.B2(n_1926),
.C1(n_1875),
.C2(n_1882),
.Y(n_1964)
);

OAI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1956),
.A2(n_1876),
.B1(n_1846),
.B2(n_1904),
.C(n_1915),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1952),
.B(n_1845),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1922),
.Y(n_1967)
);

AOI211xp5_ASAP7_75t_L g1968 ( 
.A1(n_1950),
.A2(n_1875),
.B(n_1882),
.C(n_1881),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1944),
.B(n_1853),
.Y(n_1969)
);

AOI221xp5_ASAP7_75t_L g1970 ( 
.A1(n_1925),
.A2(n_1938),
.B1(n_1959),
.B2(n_1958),
.C(n_1961),
.Y(n_1970)
);

OR2x6_ASAP7_75t_L g1971 ( 
.A(n_1962),
.B(n_1881),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1922),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1930),
.B(n_1900),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1952),
.Y(n_1974)
);

AOI31xp33_ASAP7_75t_L g1975 ( 
.A1(n_1956),
.A2(n_1842),
.A3(n_1866),
.B(n_1871),
.Y(n_1975)
);

INVx1_ASAP7_75t_SL g1976 ( 
.A(n_1952),
.Y(n_1976)
);

AOI211xp5_ASAP7_75t_L g1977 ( 
.A1(n_1950),
.A2(n_1861),
.B(n_1853),
.C(n_1896),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1950),
.A2(n_1904),
.B1(n_1915),
.B2(n_1871),
.C(n_1890),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1954),
.A2(n_1898),
.B1(n_1911),
.B2(n_1915),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1923),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1962),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1944),
.B(n_1946),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1930),
.B(n_1900),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1941),
.B(n_1885),
.Y(n_1984)
);

NAND4xp25_ASAP7_75t_SL g1985 ( 
.A(n_1938),
.B(n_1861),
.C(n_1895),
.D(n_1899),
.Y(n_1985)
);

OA21x2_ASAP7_75t_L g1986 ( 
.A1(n_1940),
.A2(n_1920),
.B(n_1909),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1954),
.A2(n_1911),
.B1(n_1913),
.B2(n_1860),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1942),
.B(n_1840),
.Y(n_1988)
);

AOI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1954),
.A2(n_1860),
.B1(n_1874),
.B2(n_1872),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1953),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1923),
.Y(n_1991)
);

OAI221xp5_ASAP7_75t_SL g1992 ( 
.A1(n_1938),
.A2(n_1895),
.B1(n_1879),
.B2(n_1851),
.C(n_1850),
.Y(n_1992)
);

AOI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1931),
.A2(n_1860),
.B1(n_1874),
.B2(n_1932),
.Y(n_1993)
);

AOI211xp5_ASAP7_75t_SL g1994 ( 
.A1(n_1948),
.A2(n_1864),
.B(n_1851),
.C(n_1862),
.Y(n_1994)
);

AOI222xp33_ASAP7_75t_L g1995 ( 
.A1(n_1947),
.A2(n_1860),
.B1(n_1887),
.B2(n_1841),
.C1(n_1842),
.C2(n_1910),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1924),
.Y(n_1996)
);

AOI222xp33_ASAP7_75t_L g1997 ( 
.A1(n_1947),
.A2(n_1887),
.B1(n_1907),
.B2(n_1905),
.C1(n_1906),
.C2(n_1899),
.Y(n_1997)
);

AND2x6_ASAP7_75t_SL g1998 ( 
.A(n_1928),
.B(n_1917),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1928),
.B(n_1908),
.Y(n_1999)
);

OAI211xp5_ASAP7_75t_L g2000 ( 
.A1(n_1960),
.A2(n_1897),
.B(n_1888),
.C(n_1850),
.Y(n_2000)
);

AO21x2_ASAP7_75t_L g2001 ( 
.A1(n_1940),
.A2(n_1843),
.B(n_1868),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1936),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1944),
.B(n_1917),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_SL g2004 ( 
.A1(n_1948),
.A2(n_1855),
.B1(n_1886),
.B2(n_1870),
.Y(n_2004)
);

OAI211xp5_ASAP7_75t_L g2005 ( 
.A1(n_1960),
.A2(n_1888),
.B(n_1858),
.C(n_1886),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1927),
.Y(n_2006)
);

OAI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1955),
.A2(n_1902),
.B1(n_1858),
.B2(n_1865),
.Y(n_2007)
);

A2O1A1Ixp33_ASAP7_75t_L g2008 ( 
.A1(n_1947),
.A2(n_1962),
.B(n_1960),
.C(n_1949),
.Y(n_2008)
);

CKINVDCx20_ASAP7_75t_R g2009 ( 
.A(n_1953),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1931),
.A2(n_1932),
.B1(n_1855),
.B2(n_1929),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1971),
.B(n_1937),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1971),
.B(n_2008),
.Y(n_2012)
);

AND2x4_ASAP7_75t_SL g2013 ( 
.A(n_2009),
.B(n_1962),
.Y(n_2013)
);

OAI21xp5_ASAP7_75t_SL g2014 ( 
.A1(n_1975),
.A2(n_1962),
.B(n_1870),
.Y(n_2014)
);

INVx4_ASAP7_75t_SL g2015 ( 
.A(n_1981),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1970),
.B(n_1937),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1986),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1976),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_2006),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1971),
.B(n_1937),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1967),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1972),
.Y(n_2022)
);

INVx4_ASAP7_75t_SL g2023 ( 
.A(n_1981),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1980),
.Y(n_2024)
);

NOR2x1p5_ASAP7_75t_L g2025 ( 
.A(n_1974),
.B(n_1962),
.Y(n_2025)
);

OA21x2_ASAP7_75t_L g2026 ( 
.A1(n_2008),
.A2(n_1933),
.B(n_1935),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1965),
.A2(n_1949),
.B(n_1929),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1991),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1977),
.B(n_2007),
.Y(n_2029)
);

NAND3xp33_ASAP7_75t_SL g2030 ( 
.A(n_1963),
.B(n_1943),
.C(n_1945),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1996),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_2001),
.Y(n_2032)
);

INVxp67_ASAP7_75t_SL g2033 ( 
.A(n_2002),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1990),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_2001),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2002),
.Y(n_2036)
);

NOR2x1_ASAP7_75t_SL g2037 ( 
.A(n_2005),
.B(n_1957),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1984),
.Y(n_2038)
);

BUFx2_ASAP7_75t_L g2039 ( 
.A(n_1998),
.Y(n_2039)
);

NAND3xp33_ASAP7_75t_L g2040 ( 
.A(n_1964),
.B(n_1962),
.C(n_1951),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1982),
.B(n_1943),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_1988),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1973),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1983),
.Y(n_2044)
);

OAI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_2000),
.A2(n_1943),
.B(n_1931),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_2010),
.B(n_1939),
.Y(n_2046)
);

INVxp67_ASAP7_75t_SL g2047 ( 
.A(n_2037),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2021),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2021),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2012),
.B(n_1969),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_2040),
.B(n_1966),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2022),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2012),
.B(n_2039),
.Y(n_2053)
);

INVx5_ASAP7_75t_L g2054 ( 
.A(n_2012),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2039),
.B(n_1994),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2039),
.B(n_2004),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_2034),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_2040),
.B(n_1966),
.Y(n_2058)
);

NAND4xp25_ASAP7_75t_SL g2059 ( 
.A(n_2016),
.B(n_2045),
.C(n_1968),
.D(n_1979),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2022),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2027),
.B(n_2003),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_2017),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2024),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2024),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2028),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2025),
.B(n_2010),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2027),
.B(n_1997),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2018),
.B(n_1999),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2011),
.B(n_1987),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2011),
.B(n_1987),
.Y(n_2070)
);

NAND4xp25_ASAP7_75t_L g2071 ( 
.A(n_2030),
.B(n_1979),
.C(n_1978),
.D(n_1992),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2020),
.B(n_1993),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2020),
.B(n_1993),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2020),
.B(n_1989),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_2034),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2026),
.B(n_1989),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_2043),
.B(n_1985),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2042),
.B(n_1995),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2042),
.B(n_2007),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2017),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2026),
.B(n_1957),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_2043),
.B(n_1936),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2031),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2044),
.B(n_1951),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_2034),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2041),
.B(n_2037),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_2013),
.B(n_1902),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2017),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2051),
.B(n_2016),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2082),
.B(n_2044),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2048),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2086),
.B(n_2015),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_2059),
.B(n_2030),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2086),
.B(n_2015),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2058),
.B(n_2044),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2048),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2049),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2049),
.Y(n_2098)
);

INVxp67_ASAP7_75t_L g2099 ( 
.A(n_2053),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2052),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2053),
.B(n_2038),
.Y(n_2101)
);

INVxp67_ASAP7_75t_SL g2102 ( 
.A(n_2047),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2052),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2054),
.B(n_2015),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2054),
.B(n_2015),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2060),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2057),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2057),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2055),
.B(n_2038),
.Y(n_2109)
);

INVx2_ASAP7_75t_SL g2110 ( 
.A(n_2054),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2055),
.B(n_2045),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2060),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2067),
.B(n_2029),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2075),
.B(n_2029),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2063),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2075),
.B(n_2041),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2085),
.B(n_2041),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_2071),
.A2(n_2056),
.B(n_2078),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2082),
.B(n_2046),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2063),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_2056),
.B(n_2014),
.Y(n_2121)
);

OR2x2_ASAP7_75t_L g2122 ( 
.A(n_2084),
.B(n_2046),
.Y(n_2122)
);

OR2x2_ASAP7_75t_L g2123 ( 
.A(n_2085),
.B(n_2046),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2064),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2054),
.B(n_2015),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2064),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2061),
.B(n_2036),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_2054),
.B(n_2023),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2065),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2123),
.B(n_2077),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2099),
.B(n_2118),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2092),
.B(n_2054),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2107),
.Y(n_2133)
);

INVxp67_ASAP7_75t_L g2134 ( 
.A(n_2121),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2091),
.Y(n_2135)
);

INVx1_ASAP7_75t_SL g2136 ( 
.A(n_2104),
.Y(n_2136)
);

INVx1_ASAP7_75t_SL g2137 ( 
.A(n_2092),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2096),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2097),
.Y(n_2139)
);

NAND2x1_ASAP7_75t_L g2140 ( 
.A(n_2128),
.B(n_2081),
.Y(n_2140)
);

NAND2x1_ASAP7_75t_SL g2141 ( 
.A(n_2104),
.B(n_2066),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_SL g2142 ( 
.A(n_2093),
.B(n_2071),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2113),
.B(n_2050),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2094),
.B(n_2050),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2094),
.B(n_2074),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2105),
.B(n_2074),
.Y(n_2146)
);

CKINVDCx20_ASAP7_75t_R g2147 ( 
.A(n_2121),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2093),
.B(n_2069),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2089),
.B(n_2107),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2108),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_2128),
.Y(n_2151)
);

INVx1_ASAP7_75t_SL g2152 ( 
.A(n_2123),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2108),
.B(n_2069),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2098),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2095),
.B(n_2077),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2100),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2105),
.B(n_2066),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_2110),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2125),
.B(n_2072),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2134),
.B(n_2102),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2133),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2133),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2145),
.B(n_2114),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2151),
.Y(n_2164)
);

AND2x4_ASAP7_75t_SL g2165 ( 
.A(n_2132),
.B(n_2128),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2142),
.B(n_2111),
.Y(n_2166)
);

INVxp67_ASAP7_75t_L g2167 ( 
.A(n_2145),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2133),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_2146),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2150),
.Y(n_2170)
);

INVxp67_ASAP7_75t_SL g2171 ( 
.A(n_2141),
.Y(n_2171)
);

A2O1A1Ixp33_ASAP7_75t_L g2172 ( 
.A1(n_2142),
.A2(n_2014),
.B(n_2076),
.C(n_2125),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2144),
.B(n_2109),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2150),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_2151),
.B(n_2110),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2159),
.B(n_2101),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_2147),
.B(n_2127),
.Y(n_2177)
);

AOI21xp33_ASAP7_75t_SL g2178 ( 
.A1(n_2148),
.A2(n_2079),
.B(n_2119),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2150),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2151),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_R g2181 ( 
.A(n_2131),
.B(n_2152),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2135),
.Y(n_2182)
);

INVx2_ASAP7_75t_SL g2183 ( 
.A(n_2165),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2165),
.B(n_2144),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_SL g2185 ( 
.A1(n_2166),
.A2(n_2137),
.B(n_2149),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2171),
.B(n_2159),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2180),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2173),
.B(n_2146),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_2163),
.B(n_2143),
.Y(n_2189)
);

OAI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_2166),
.A2(n_2141),
.B(n_2132),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2169),
.B(n_2157),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2167),
.B(n_2136),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2180),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2177),
.B(n_2136),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2175),
.B(n_2157),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_2177),
.B(n_2155),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2175),
.B(n_2151),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_2164),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2178),
.B(n_2153),
.Y(n_2199)
);

NOR3xp33_ASAP7_75t_L g2200 ( 
.A(n_2194),
.B(n_2160),
.C(n_2176),
.Y(n_2200)
);

OAI221xp5_ASAP7_75t_SL g2201 ( 
.A1(n_2185),
.A2(n_2172),
.B1(n_2155),
.B2(n_2130),
.C(n_2181),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2195),
.B(n_2188),
.Y(n_2202)
);

AOI211xp5_ASAP7_75t_SL g2203 ( 
.A1(n_2196),
.A2(n_2158),
.B(n_2172),
.C(n_2179),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2195),
.B(n_2181),
.Y(n_2204)
);

XNOR2x2_ASAP7_75t_L g2205 ( 
.A(n_2190),
.B(n_2161),
.Y(n_2205)
);

AOI211xp5_ASAP7_75t_L g2206 ( 
.A1(n_2196),
.A2(n_2130),
.B(n_2182),
.C(n_2170),
.Y(n_2206)
);

NAND3xp33_ASAP7_75t_L g2207 ( 
.A(n_2183),
.B(n_2168),
.C(n_2162),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2188),
.B(n_2174),
.Y(n_2208)
);

O2A1O1Ixp5_ASAP7_75t_L g2209 ( 
.A1(n_2199),
.A2(n_2140),
.B(n_2154),
.C(n_2156),
.Y(n_2209)
);

O2A1O1Ixp33_ASAP7_75t_L g2210 ( 
.A1(n_2183),
.A2(n_2156),
.B(n_2154),
.C(n_2139),
.Y(n_2210)
);

OAI21xp33_ASAP7_75t_L g2211 ( 
.A1(n_2184),
.A2(n_2117),
.B(n_2116),
.Y(n_2211)
);

AOI222xp33_ASAP7_75t_L g2212 ( 
.A1(n_2186),
.A2(n_2139),
.B1(n_2138),
.B2(n_2135),
.C1(n_2076),
.C2(n_2070),
.Y(n_2212)
);

O2A1O1Ixp5_ASAP7_75t_L g2213 ( 
.A1(n_2203),
.A2(n_2140),
.B(n_2184),
.C(n_2192),
.Y(n_2213)
);

NAND5xp2_ASAP7_75t_L g2214 ( 
.A(n_2201),
.B(n_2191),
.C(n_2197),
.D(n_2193),
.E(n_2187),
.Y(n_2214)
);

AOI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2204),
.A2(n_2191),
.B1(n_2198),
.B2(n_2189),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_2206),
.B(n_2119),
.Y(n_2216)
);

OAI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2209),
.A2(n_2138),
.B(n_2122),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2202),
.A2(n_2106),
.B(n_2103),
.Y(n_2218)
);

AOI221xp5_ASAP7_75t_L g2219 ( 
.A1(n_2200),
.A2(n_2129),
.B1(n_2126),
.B2(n_2124),
.C(n_2112),
.Y(n_2219)
);

NAND3xp33_ASAP7_75t_L g2220 ( 
.A(n_2213),
.B(n_2207),
.C(n_2212),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2215),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2216),
.B(n_2208),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2217),
.B(n_2211),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2218),
.B(n_2210),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2219),
.B(n_2115),
.Y(n_2225)
);

NOR2x1_ASAP7_75t_SL g2226 ( 
.A(n_2214),
.B(n_2120),
.Y(n_2226)
);

O2A1O1Ixp33_ASAP7_75t_SL g2227 ( 
.A1(n_2224),
.A2(n_2205),
.B(n_2019),
.C(n_2033),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2222),
.B(n_2072),
.Y(n_2228)
);

NOR3xp33_ASAP7_75t_SL g2229 ( 
.A(n_2220),
.B(n_2221),
.C(n_2225),
.Y(n_2229)
);

AOI21xp5_ASAP7_75t_L g2230 ( 
.A1(n_2226),
.A2(n_2122),
.B(n_2090),
.Y(n_2230)
);

HB1xp67_ASAP7_75t_L g2231 ( 
.A(n_2223),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2225),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2228),
.B(n_2090),
.Y(n_2233)
);

OR2x2_ASAP7_75t_L g2234 ( 
.A(n_2231),
.B(n_2068),
.Y(n_2234)
);

NOR3xp33_ASAP7_75t_L g2235 ( 
.A(n_2232),
.B(n_2087),
.C(n_2070),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2233),
.Y(n_2236)
);

OAI22xp5_ASAP7_75t_SL g2237 ( 
.A1(n_2236),
.A2(n_2234),
.B1(n_2229),
.B2(n_2227),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_2237),
.Y(n_2238)
);

AOI21xp5_ASAP7_75t_L g2239 ( 
.A1(n_2237),
.A2(n_2230),
.B(n_2235),
.Y(n_2239)
);

OAI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2239),
.A2(n_2238),
.B(n_2080),
.Y(n_2240)
);

OAI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_2238),
.A2(n_2088),
.B1(n_2062),
.B2(n_2080),
.Y(n_2241)
);

OAI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_2240),
.A2(n_2088),
.B1(n_2062),
.B2(n_2080),
.Y(n_2242)
);

HB1xp67_ASAP7_75t_L g2243 ( 
.A(n_2241),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2243),
.Y(n_2244)
);

INVxp33_ASAP7_75t_L g2245 ( 
.A(n_2244),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_2245),
.B(n_2242),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_2246),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2247),
.A2(n_2088),
.B1(n_2062),
.B2(n_2073),
.Y(n_2248)
);

AOI211xp5_ASAP7_75t_L g2249 ( 
.A1(n_2248),
.A2(n_2035),
.B(n_2032),
.C(n_2083),
.Y(n_2249)
);


endmodule