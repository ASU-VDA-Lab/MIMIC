module real_aes_7176_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_0), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_1), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_2), .A2(n_185), .B1(n_368), .B2(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g318 ( .A(n_3), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_4), .A2(n_89), .B1(n_406), .B2(n_407), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_5), .A2(n_17), .B1(n_410), .B2(n_411), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g296 ( .A(n_6), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_7), .A2(n_19), .B1(n_463), .B2(n_464), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_8), .B(n_508), .Y(n_507) );
AOI222xp33_ASAP7_75t_L g510 ( .A1(n_9), .A2(n_66), .B1(n_207), .B2(n_280), .C1(n_348), .C2(n_397), .Y(n_510) );
INVx1_ASAP7_75t_L g312 ( .A(n_10), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_11), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_12), .A2(n_105), .B1(n_418), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_13), .A2(n_52), .B1(n_678), .B2(n_680), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_14), .A2(n_141), .B1(n_349), .B2(n_483), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_15), .A2(n_98), .B1(n_369), .B2(n_475), .Y(n_648) );
AOI222xp33_ASAP7_75t_L g609 ( .A1(n_16), .A2(n_100), .B1(n_175), .B2(n_398), .C1(n_406), .C2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_18), .A2(n_116), .B1(n_386), .B2(n_389), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_20), .Y(n_288) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_21), .A2(n_136), .B1(n_450), .B2(n_451), .Y(n_449) );
AOI222xp33_ASAP7_75t_L g484 ( .A1(n_22), .A2(n_65), .B1(n_117), .B2(n_410), .C1(n_485), .C2(n_486), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_23), .B(n_389), .Y(n_558) );
INVx1_ASAP7_75t_L g667 ( .A(n_24), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_24), .A2(n_667), .B1(n_671), .B2(n_704), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_25), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_26), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_27), .Y(n_354) );
AO22x2_ASAP7_75t_L g243 ( .A1(n_28), .A2(n_67), .B1(n_244), .B2(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g626 ( .A(n_28), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_29), .B(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_30), .A2(n_158), .B1(n_418), .B2(n_424), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g334 ( .A1(n_31), .A2(n_220), .B1(n_290), .B2(n_335), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_32), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_33), .A2(n_221), .B1(n_333), .B2(n_420), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_34), .A2(n_57), .B1(n_503), .B2(n_685), .Y(n_684) );
AOI222xp33_ASAP7_75t_L g396 ( .A1(n_35), .A2(n_157), .B1(n_202), .B2(n_348), .C1(n_397), .C2(n_398), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_36), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_37), .A2(n_199), .B1(n_335), .B2(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_38), .B(n_386), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_39), .A2(n_143), .B1(n_394), .B2(n_446), .Y(n_445) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_40), .A2(n_71), .B1(n_244), .B2(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g627 ( .A(n_40), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_41), .A2(n_111), .B1(n_255), .B2(n_259), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_42), .A2(n_213), .B1(n_413), .B2(n_414), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_43), .A2(n_64), .B1(n_471), .B2(n_473), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_44), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_45), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_46), .A2(n_102), .B1(n_468), .B2(n_522), .Y(n_521) );
AOI222xp33_ASAP7_75t_L g592 ( .A1(n_47), .A2(n_153), .B1(n_208), .B2(n_280), .C1(n_397), .C2(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_48), .A2(n_56), .B1(n_335), .B2(n_572), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_49), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_50), .A2(n_178), .B1(n_375), .B2(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_51), .A2(n_125), .B1(n_349), .B2(n_411), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_53), .A2(n_148), .B1(n_420), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_54), .A2(n_160), .B1(n_368), .B2(n_420), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_55), .Y(n_340) );
XNOR2x2_ASAP7_75t_L g491 ( .A(n_58), .B(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_59), .A2(n_132), .B1(n_540), .B2(n_541), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_60), .A2(n_194), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_61), .A2(n_181), .B1(n_480), .B2(n_481), .Y(n_479) );
AOI22xp5_ASAP7_75t_SL g321 ( .A1(n_62), .A2(n_123), .B1(n_322), .B2(n_324), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_63), .A2(n_124), .B1(n_333), .B2(n_418), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_68), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_69), .A2(n_115), .B1(n_410), .B2(n_541), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_70), .A2(n_216), .B1(n_372), .B2(n_373), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_72), .A2(n_167), .B1(n_286), .B2(n_381), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_73), .Y(n_595) );
AND2x2_ASAP7_75t_L g229 ( .A(n_74), .B(n_230), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_75), .A2(n_210), .B1(n_377), .B2(n_380), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_76), .A2(n_106), .B1(n_472), .B2(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g573 ( .A(n_77), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_78), .A2(n_164), .B1(n_420), .B2(n_421), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_79), .A2(n_113), .B1(n_475), .B2(n_477), .Y(n_474) );
AOI22xp5_ASAP7_75t_SL g330 ( .A1(n_80), .A2(n_191), .B1(n_331), .B2(n_333), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_81), .A2(n_150), .B1(n_348), .B2(n_349), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_82), .Y(n_524) );
INVx1_ASAP7_75t_L g226 ( .A(n_83), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_84), .A2(n_135), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_85), .A2(n_121), .B1(n_255), .B2(n_280), .Y(n_440) );
XOR2x2_ASAP7_75t_L g359 ( .A(n_86), .B(n_360), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_87), .A2(n_151), .B1(n_450), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g264 ( .A(n_88), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_90), .A2(n_128), .B1(n_446), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_91), .A2(n_197), .B1(n_580), .B2(n_604), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_92), .A2(n_630), .B1(n_658), .B2(n_659), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_92), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_93), .A2(n_177), .B1(n_280), .B2(n_411), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_94), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_95), .A2(n_139), .B1(n_298), .B2(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_96), .B(n_386), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_97), .A2(n_145), .B1(n_418), .B2(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_99), .B(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_101), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_103), .B(n_414), .Y(n_543) );
INVx1_ASAP7_75t_L g562 ( .A(n_104), .Y(n_562) );
INVx1_ASAP7_75t_L g316 ( .A(n_107), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_108), .A2(n_189), .B1(n_381), .B2(n_425), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_109), .A2(n_192), .B1(n_349), .B2(n_392), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_110), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_112), .A2(n_223), .B(n_231), .C(n_628), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_114), .A2(n_217), .B1(n_377), .B2(n_468), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_118), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_119), .Y(n_611) );
INVx2_ASAP7_75t_L g230 ( .A(n_120), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_122), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_126), .A2(n_187), .B1(n_259), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_127), .A2(n_170), .B1(n_392), .B2(n_407), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_129), .Y(n_634) );
AND2x6_ASAP7_75t_L g225 ( .A(n_130), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_130), .Y(n_620) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_131), .A2(n_186), .B1(n_244), .B2(n_248), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_133), .A2(n_205), .B1(n_328), .B2(n_421), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_134), .A2(n_165), .B1(n_455), .B2(n_582), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g273 ( .A(n_137), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_138), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_140), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_142), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_144), .Y(n_352) );
AOI22xp33_ASAP7_75t_SL g570 ( .A1(n_146), .A2(n_159), .B1(n_425), .B2(n_528), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_147), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g453 ( .A1(n_149), .A2(n_203), .B1(n_333), .B2(n_418), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_152), .Y(n_457) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_154), .A2(n_200), .B1(n_244), .B2(n_245), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_155), .A2(n_215), .B1(n_406), .B2(n_446), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_156), .Y(n_654) );
INVx1_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_162), .A2(n_172), .B1(n_467), .B2(n_468), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_163), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_166), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_168), .Y(n_703) );
INVx1_ASAP7_75t_L g309 ( .A(n_169), .Y(n_309) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_171), .A2(n_204), .B1(n_455), .B2(n_456), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_173), .B(n_290), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_174), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_176), .A2(n_201), .B1(n_381), .B2(n_591), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_179), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_180), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_182), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_183), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_184), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_186), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_188), .B(n_414), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_190), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_193), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_195), .A2(n_206), .B1(n_414), .B2(n_508), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_196), .A2(n_513), .B1(n_514), .B2(n_547), .Y(n_512) );
INVx1_ASAP7_75t_L g547 ( .A(n_196), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_198), .Y(n_692) );
INVx1_ASAP7_75t_L g623 ( .A(n_200), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_209), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_211), .A2(n_214), .B1(n_363), .B2(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g244 ( .A(n_212), .Y(n_244) );
INVx1_ASAP7_75t_L g246 ( .A(n_212), .Y(n_246) );
OA22x2_ASAP7_75t_L g458 ( .A1(n_218), .A2(n_459), .B1(n_460), .B2(n_487), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_218), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_219), .Y(n_403) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_226), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_227), .A2(n_618), .B(n_666), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_550), .B1(n_551), .B2(n_614), .C(n_615), .Y(n_231) );
INVxp67_ASAP7_75t_L g614 ( .A(n_232), .Y(n_614) );
XNOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_431), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_355), .B1(n_356), .B2(n_430), .Y(n_233) );
INVx2_ASAP7_75t_L g430 ( .A(n_234), .Y(n_430) );
XOR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_317), .Y(n_234) );
XNOR2x1_ASAP7_75t_L g235 ( .A(n_236), .B(n_316), .Y(n_235) );
AND3x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_283), .C(n_300), .Y(n_236) );
NOR3xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_263), .C(n_272), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_254), .Y(n_238) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_240), .Y(n_345) );
OAI22xp5_ASAP7_75t_SL g633 ( .A1(n_240), .A2(n_265), .B1(n_634), .B2(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g691 ( .A(n_240), .Y(n_691) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_249), .Y(n_240) );
INVx2_ASAP7_75t_L g315 ( .A(n_241), .Y(n_315) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_247), .Y(n_241) );
AND2x2_ASAP7_75t_L g267 ( .A(n_242), .B(n_247), .Y(n_267) );
AND2x2_ASAP7_75t_L g287 ( .A(n_242), .B(n_271), .Y(n_287) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g258 ( .A(n_243), .B(n_253), .Y(n_258) );
AND2x2_ASAP7_75t_L g262 ( .A(n_243), .B(n_247), .Y(n_262) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g248 ( .A(n_246), .Y(n_248) );
INVx2_ASAP7_75t_L g271 ( .A(n_247), .Y(n_271) );
INVx1_ASAP7_75t_L g383 ( .A(n_247), .Y(n_383) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_250), .B(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g286 ( .A(n_250), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g388 ( .A(n_250), .B(n_315), .Y(n_388) );
AND2x6_ASAP7_75t_L g390 ( .A(n_250), .B(n_267), .Y(n_390) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g257 ( .A(n_251), .Y(n_257) );
INVx1_ASAP7_75t_L g261 ( .A(n_251), .Y(n_261) );
INVx1_ASAP7_75t_L g277 ( .A(n_251), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_251), .B(n_253), .Y(n_292) );
AND2x2_ASAP7_75t_L g276 ( .A(n_252), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g307 ( .A(n_253), .B(n_261), .Y(n_307) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_255), .Y(n_348) );
BUFx12f_ASAP7_75t_L g406 ( .A(n_255), .Y(n_406) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g282 ( .A(n_257), .B(n_271), .Y(n_282) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_258), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g281 ( .A(n_258), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g394 ( .A(n_258), .B(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_259), .Y(n_349) );
BUFx2_ASAP7_75t_SL g407 ( .A(n_259), .Y(n_407) );
BUFx3_ASAP7_75t_L g446 ( .A(n_259), .Y(n_446) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx1_ASAP7_75t_L g644 ( .A(n_260), .Y(n_644) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x6_ASAP7_75t_L g275 ( .A(n_262), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g643 ( .A(n_262), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B1(n_268), .B2(n_269), .Y(n_263) );
OA211x2_ASAP7_75t_L g605 ( .A1(n_265), .A2(n_606), .B(n_607), .C(n_608), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_265), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_688) );
BUFx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g339 ( .A(n_266), .Y(n_339) );
AND2x4_ASAP7_75t_L g298 ( .A(n_267), .B(n_276), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_267), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g326 ( .A(n_267), .B(n_307), .Y(n_326) );
INVx4_ASAP7_75t_L g342 ( .A(n_269), .Y(n_342) );
AND2x2_ASAP7_75t_L g290 ( .A(n_270), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_278), .B2(n_279), .Y(n_272) );
INVx2_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
INVx4_ASAP7_75t_L g351 ( .A(n_275), .Y(n_351) );
INVx2_ASAP7_75t_L g404 ( .A(n_275), .Y(n_404) );
BUFx3_ASAP7_75t_L g485 ( .A(n_275), .Y(n_485) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_275), .Y(n_610) );
INVx2_ASAP7_75t_L g696 ( .A(n_275), .Y(n_696) );
AND2x2_ASAP7_75t_L g295 ( .A(n_276), .B(n_287), .Y(n_295) );
AND2x6_ASAP7_75t_L g314 ( .A(n_276), .B(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g540 ( .A(n_279), .Y(n_540) );
INVx4_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g353 ( .A(n_280), .Y(n_353) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_281), .Y(n_398) );
BUFx4f_ASAP7_75t_SL g410 ( .A(n_281), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_284), .B(n_293), .Y(n_283) );
OAI21xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_288), .B(n_289), .Y(n_284) );
OAI221xp5_ASAP7_75t_SL g681 ( .A1(n_285), .A2(n_303), .B1(n_682), .B2(n_683), .C(n_684), .Y(n_681) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_286), .Y(n_335) );
BUFx3_ASAP7_75t_L g368 ( .A(n_286), .Y(n_368) );
BUFx3_ASAP7_75t_L g589 ( .A(n_286), .Y(n_589) );
BUFx3_ASAP7_75t_L g604 ( .A(n_286), .Y(n_604) );
AND2x4_ASAP7_75t_L g304 ( .A(n_287), .B(n_291), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_287), .B(n_307), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_287), .B(n_307), .Y(n_323) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x6_ASAP7_75t_L g382 ( .A(n_292), .B(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .B1(n_297), .B2(n_299), .Y(n_293) );
INVx3_ASAP7_75t_L g328 ( .A(n_294), .Y(n_328) );
INVx3_ASAP7_75t_L g420 ( .A(n_294), .Y(n_420) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_SL g372 ( .A(n_295), .Y(n_372) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_295), .Y(n_472) );
BUFx2_ASAP7_75t_SL g532 ( .A(n_295), .Y(n_532) );
INVx3_ASAP7_75t_L g424 ( .A(n_297), .Y(n_424) );
INVx2_ASAP7_75t_L g463 ( .A(n_297), .Y(n_463) );
INVx2_ASAP7_75t_L g582 ( .A(n_297), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_297), .A2(n_651), .B1(n_652), .B2(n_654), .Y(n_650) );
INVx6_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx3_ASAP7_75t_L g375 ( .A(n_298), .Y(n_375) );
BUFx3_ASAP7_75t_L g456 ( .A(n_298), .Y(n_456) );
BUFx3_ASAP7_75t_L g528 ( .A(n_298), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_308), .C(n_311), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_305), .B2(n_306), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
BUFx3_ASAP7_75t_L g369 ( .A(n_304), .Y(n_369) );
BUFx2_ASAP7_75t_L g477 ( .A(n_304), .Y(n_477) );
BUFx2_ASAP7_75t_SL g497 ( .A(n_304), .Y(n_497) );
BUFx3_ASAP7_75t_L g580 ( .A(n_304), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g535 ( .A(n_310), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx5_ASAP7_75t_SL g421 ( .A(n_313), .Y(n_421) );
INVx1_ASAP7_75t_L g495 ( .A(n_313), .Y(n_495) );
INVx2_ASAP7_75t_SL g567 ( .A(n_313), .Y(n_567) );
INVx4_ASAP7_75t_L g653 ( .A(n_313), .Y(n_653) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_313), .Y(n_674) );
INVx11_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx11_ASAP7_75t_L g332 ( .A(n_314), .Y(n_332) );
XNOR2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NAND3x1_ASAP7_75t_SL g319 ( .A(n_320), .B(n_329), .C(n_336), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_327), .Y(n_320) );
INVx1_ASAP7_75t_L g465 ( .A(n_322), .Y(n_465) );
BUFx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx3_ASAP7_75t_L g366 ( .A(n_323), .Y(n_366) );
BUFx3_ASAP7_75t_L g418 ( .A(n_323), .Y(n_418) );
BUFx3_ASAP7_75t_L g501 ( .A(n_323), .Y(n_501) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx4_ASAP7_75t_L g379 ( .A(n_325), .Y(n_379) );
INVx5_ASAP7_75t_L g425 ( .A(n_325), .Y(n_425) );
INVx1_ASAP7_75t_L g450 ( .A(n_325), .Y(n_450) );
INVx2_ASAP7_75t_L g591 ( .A(n_325), .Y(n_591) );
BUFx3_ASAP7_75t_L g686 ( .A(n_325), .Y(n_686) );
INVx8_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_334), .Y(n_329) );
INVx4_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx4_ASAP7_75t_L g363 ( .A(n_332), .Y(n_363) );
INVx3_ASAP7_75t_L g455 ( .A(n_332), .Y(n_455) );
INVx2_ASAP7_75t_SL g473 ( .A(n_332), .Y(n_473) );
INVx4_ASAP7_75t_L g476 ( .A(n_335), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_344), .C(n_350), .Y(n_336) );
OAI22xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_340), .B1(n_341), .B2(n_343), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g506 ( .A(n_339), .Y(n_506) );
OAI22xp5_ASAP7_75t_SL g639 ( .A1(n_341), .A2(n_640), .B1(n_641), .B2(n_645), .Y(n_639) );
INVx3_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g698 ( .A(n_342), .Y(n_698) );
OAI21xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_346), .B(n_347), .Y(n_344) );
BUFx4f_ASAP7_75t_L g541 ( .A(n_348), .Y(n_541) );
OAI22xp5_ASAP7_75t_SL g350 ( .A1(n_351), .A2(n_352), .B1(n_353), .B2(n_354), .Y(n_350) );
INVx4_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
OAI21xp5_ASAP7_75t_SL g537 ( .A1(n_351), .A2(n_538), .B(n_539), .Y(n_537) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_351), .A2(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AO22x1_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_399), .B1(n_428), .B2(n_429), .Y(n_358) );
INVx1_ASAP7_75t_L g428 ( .A(n_359), .Y(n_428) );
NAND4xp75_ASAP7_75t_L g360 ( .A(n_361), .B(n_370), .C(n_384), .D(n_396), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_367), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g520 ( .A(n_369), .Y(n_520) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_376), .Y(n_370) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI221xp5_ASAP7_75t_SL g673 ( .A1(n_374), .A2(n_674), .B1(n_675), .B2(n_676), .C(n_677), .Y(n_673) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx2_ASAP7_75t_L g467 ( .A(n_379), .Y(n_467) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_379), .Y(n_522) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g451 ( .A(n_381), .Y(n_451) );
BUFx2_ASAP7_75t_L g468 ( .A(n_381), .Y(n_468) );
INVx6_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g503 ( .A(n_382), .Y(n_503) );
INVx1_ASAP7_75t_SL g572 ( .A(n_382), .Y(n_572) );
INVx1_ASAP7_75t_L g395 ( .A(n_383), .Y(n_395) );
AND2x2_ASAP7_75t_SL g384 ( .A(n_385), .B(n_391), .Y(n_384) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx5_ASAP7_75t_L g413 ( .A(n_387), .Y(n_413) );
INVx2_ASAP7_75t_L g444 ( .A(n_387), .Y(n_444) );
INVx2_ASAP7_75t_L g508 ( .A(n_387), .Y(n_508) );
INVx4_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx4f_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
BUFx2_ASAP7_75t_L g481 ( .A(n_390), .Y(n_481) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx3_ASAP7_75t_L g411 ( .A(n_394), .Y(n_411) );
BUFx2_ASAP7_75t_L g483 ( .A(n_394), .Y(n_483) );
BUFx2_ASAP7_75t_L g586 ( .A(n_394), .Y(n_586) );
INVx3_ASAP7_75t_SL g429 ( .A(n_399), .Y(n_429) );
XOR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_427), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_415), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_408), .Y(n_401) );
OAI21xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B(n_405), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_404), .A2(n_439), .B(n_440), .Y(n_438) );
OAI21xp5_ASAP7_75t_SL g561 ( .A1(n_404), .A2(n_562), .B(n_563), .Y(n_561) );
BUFx4f_ASAP7_75t_SL g486 ( .A(n_406), .Y(n_486) );
INVx2_ASAP7_75t_L g594 ( .A(n_406), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g694 ( .A(n_410), .Y(n_694) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_413), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_422), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
BUFx3_ASAP7_75t_L g680 ( .A(n_418), .Y(n_680) );
INVx1_ASAP7_75t_L g525 ( .A(n_421), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_426), .Y(n_422) );
AOI22xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_433), .B1(n_489), .B2(n_490), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B1(n_458), .B2(n_488), .Y(n_433) );
INVx4_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
XOR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_457), .Y(n_435) );
NAND3x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_447), .C(n_452), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .C(n_445), .Y(n_441) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g488 ( .A(n_458), .Y(n_488) );
INVx1_ASAP7_75t_SL g487 ( .A(n_460), .Y(n_487) );
NAND4xp75_ASAP7_75t_L g460 ( .A(n_461), .B(n_469), .C(n_478), .D(n_484), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g679 ( .A(n_472), .Y(n_679) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx4_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_479), .B(n_482), .Y(n_478) );
INVx1_ASAP7_75t_L g702 ( .A(n_486), .Y(n_702) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_511), .B1(n_548), .B2(n_549), .Y(n_490) );
INVx1_ASAP7_75t_L g549 ( .A(n_491), .Y(n_549) );
NAND4xp75_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .C(n_504), .D(n_510), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_502), .Y(n_498) );
BUFx4f_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OA211x2_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_507), .C(n_509), .Y(n_504) );
INVx1_ASAP7_75t_L g548 ( .A(n_511), .Y(n_548) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_515), .B(n_536), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_523), .C(n_529), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_526), .B2(n_527), .Y(n_523) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_533), .B2(n_534), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_531), .A2(n_534), .B1(n_656), .B2(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_542), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .C(n_546), .Y(n_542) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B1(n_574), .B2(n_575), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
XOR2x2_ASAP7_75t_SL g554 ( .A(n_555), .B(n_573), .Y(n_554) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_556), .B(n_564), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .C(n_560), .Y(n_557) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AO22x1_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_596), .B1(n_612), .B2(n_613), .Y(n_575) );
INVx2_ASAP7_75t_SL g612 ( .A(n_576), .Y(n_612) );
XOR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_595), .Y(n_576) );
NAND4xp75_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .C(n_587), .D(n_592), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_SL g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_SL g613 ( .A(n_596), .Y(n_613) );
XOR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_611), .Y(n_596) );
NAND4xp75_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .C(n_605), .D(n_609), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NOR2x1_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .Y(n_616) );
OR2x2_ASAP7_75t_SL g707 ( .A(n_617), .B(n_622), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_619), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_619), .B(n_663), .Y(n_666) );
CKINVDCx16_ASAP7_75t_R g663 ( .A(n_620), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
OAI322xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_660), .A3(n_661), .B1(n_664), .B2(n_667), .C1(n_668), .C2(n_705), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_630), .Y(n_659) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_646), .Y(n_631) );
NOR3xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_636), .C(n_639), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_641), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x6_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_650), .C(n_655), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g704 ( .A(n_671), .Y(n_704) );
AND2x2_ASAP7_75t_SL g671 ( .A(n_672), .B(n_687), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_681), .Y(n_672) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_693), .C(n_700), .Y(n_687) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
OAI222xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_699), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_707), .Y(n_706) );
endmodule