module fake_jpeg_337_n_659 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_659);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_659;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g180 ( 
.A(n_59),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_60),
.B(n_63),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g224 ( 
.A(n_61),
.Y(n_224)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_71),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_75),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_25),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_76),
.Y(n_134)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_77),
.Y(n_189)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_79),
.Y(n_225)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_80),
.Y(n_181)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_83),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_32),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_87),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_17),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_90),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_17),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_100),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_20),
.B(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_94),
.B(n_108),
.Y(n_148)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx12f_ASAP7_75t_SL g96 ( 
.A(n_26),
.Y(n_96)
);

BUFx12f_ASAP7_75t_SL g194 ( 
.A(n_96),
.Y(n_194)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_39),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_101),
.Y(n_208)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_102),
.Y(n_210)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_104),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_105),
.B(n_106),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_20),
.B(n_19),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_110),
.Y(n_227)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_29),
.B(n_14),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_112),
.B(n_118),
.Y(n_204)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_24),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_117),
.B(n_119),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_36),
.B(n_41),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_41),
.B(n_15),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_40),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_24),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_127),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_124),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_33),
.B(n_31),
.C(n_35),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_24),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_57),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_128),
.B(n_52),
.Y(n_201)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_26),
.Y(n_129)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_30),
.Y(n_130)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_133),
.B(n_161),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_81),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_162),
.B(n_195),
.Y(n_243)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_164),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_77),
.Y(n_168)
);

INVx11_ASAP7_75t_L g247 ( 
.A(n_168),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_59),
.Y(n_169)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_68),
.B(n_52),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_171),
.Y(n_262)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_172),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_174),
.B(n_57),
.Y(n_238)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_76),
.Y(n_183)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_185),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_126),
.B(n_50),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_188),
.B(n_206),
.Y(n_260)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_70),
.Y(n_192)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_93),
.Y(n_195)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_83),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_65),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_199),
.Y(n_291)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_205),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_44),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_121),
.B(n_44),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_211),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_64),
.B(n_43),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_111),
.Y(n_212)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_66),
.Y(n_213)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_73),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_96),
.B(n_54),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_43),
.C(n_56),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_79),
.B(n_31),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_52),
.Y(n_230)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_95),
.Y(n_218)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_82),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_222),
.Y(n_250)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_84),
.Y(n_221)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_83),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_103),
.Y(n_223)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_223),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g352 ( 
.A1(n_230),
.A2(n_238),
.B(n_241),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_180),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_232),
.B(n_237),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_234),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_131),
.A2(n_124),
.B1(n_120),
.B2(n_88),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_235),
.A2(n_254),
.B1(n_255),
.B2(n_259),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_54),
.B1(n_109),
.B2(n_74),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_236),
.A2(n_301),
.B1(n_159),
.B2(n_165),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_37),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_188),
.A2(n_37),
.B1(n_56),
.B2(n_55),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_239),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_246),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_249),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_148),
.A2(n_143),
.B1(n_142),
.B2(n_226),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_142),
.A2(n_92),
.B1(n_116),
.B2(n_101),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_145),
.Y(n_256)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_256),
.Y(n_340)
);

BUFx12_ASAP7_75t_L g257 ( 
.A(n_151),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_257),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_143),
.A2(n_99),
.B1(n_69),
.B2(n_54),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_264),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_23),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_270),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_145),
.Y(n_266)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_146),
.Y(n_267)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_146),
.Y(n_269)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_204),
.B(n_23),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_160),
.B(n_55),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_288),
.Y(n_330)
);

CKINVDCx12_ASAP7_75t_R g274 ( 
.A(n_169),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_274),
.Y(n_350)
);

BUFx12f_ASAP7_75t_L g276 ( 
.A(n_151),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_276),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_163),
.Y(n_277)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_277),
.Y(n_346)
);

CKINVDCx12_ASAP7_75t_R g278 ( 
.A(n_134),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_189),
.Y(n_279)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_178),
.B(n_147),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_280),
.A2(n_297),
.B(n_298),
.Y(n_311)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_281),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_135),
.A2(n_125),
.B1(n_123),
.B2(n_57),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_282),
.A2(n_283),
.B1(n_306),
.B2(n_139),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_135),
.A2(n_47),
.B1(n_35),
.B2(n_33),
.Y(n_283)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_182),
.Y(n_285)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_225),
.Y(n_286)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_154),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_190),
.Y(n_289)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_155),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_290),
.B(n_294),
.Y(n_343)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_191),
.Y(n_292)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_149),
.Y(n_293)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_141),
.B(n_47),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_141),
.B(n_53),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_302),
.Y(n_344)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_163),
.Y(n_296)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_296),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_187),
.B(n_1),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_187),
.B(n_1),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_167),
.Y(n_299)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_166),
.Y(n_300)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_155),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_301)
);

CKINVDCx9p33_ASAP7_75t_R g302 ( 
.A(n_134),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_181),
.Y(n_303)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_137),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_305),
.A2(n_170),
.B1(n_3),
.B2(n_5),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_140),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_175),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_308),
.Y(n_322)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_150),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_156),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_309),
.B(n_310),
.Y(n_370)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_166),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_238),
.A2(n_176),
.B1(n_171),
.B2(n_227),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_313),
.A2(n_354),
.B1(n_307),
.B2(n_231),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_223),
.B1(n_220),
.B2(n_197),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_314),
.A2(n_336),
.B(n_347),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_316),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_245),
.A2(n_159),
.B1(n_217),
.B2(n_210),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_260),
.B(n_152),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_321),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_320),
.A2(n_334),
.B1(n_357),
.B2(n_256),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_261),
.B(n_158),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_229),
.B(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_328),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_262),
.A2(n_177),
.B1(n_208),
.B2(n_170),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_230),
.A2(n_190),
.B(n_138),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_244),
.B(n_168),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_341),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_301),
.A2(n_132),
.B1(n_144),
.B2(n_153),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_299),
.A2(n_227),
.B1(n_184),
.B2(n_186),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_348),
.A2(n_246),
.B(n_240),
.Y(n_389)
);

A2O1A1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_237),
.A2(n_198),
.B(n_136),
.C(n_184),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_349),
.B(n_234),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_243),
.B(n_209),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_356),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_263),
.B(n_157),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g408 ( 
.A(n_353),
.B(n_355),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_235),
.A2(n_208),
.B1(n_186),
.B2(n_177),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_271),
.B(n_173),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_265),
.B(n_173),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_268),
.B(n_2),
.C(n_6),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_359),
.B(n_360),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_252),
.B(n_258),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_275),
.B(n_2),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_364),
.B(n_369),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_250),
.B(n_2),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_364),
.Y(n_379)
);

AOI32xp33_ASAP7_75t_L g367 ( 
.A1(n_248),
.A2(n_7),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_306),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_272),
.B(n_12),
.Y(n_369)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_236),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_372),
.B(n_401),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_319),
.B(n_228),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_382),
.Y(n_427)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_322),
.Y(n_376)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_379),
.B(n_383),
.Y(n_428)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_342),
.Y(n_380)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_322),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_328),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_384),
.A2(n_394),
.B(n_341),
.Y(n_447)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_322),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_386),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_330),
.B(n_231),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_387),
.B(n_390),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_318),
.A2(n_310),
.B1(n_269),
.B2(n_296),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_388),
.A2(n_395),
.B1(n_399),
.B2(n_402),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_389),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_328),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_343),
.B(n_287),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_391),
.B(n_396),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_321),
.B(n_272),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_409),
.Y(n_420)
);

OR2x2_ASAP7_75t_SL g394 ( 
.A(n_336),
.B(n_284),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_314),
.A2(n_300),
.B1(n_266),
.B2(n_267),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_335),
.B(n_291),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_356),
.B(n_366),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_357),
.A2(n_277),
.B1(n_286),
.B2(n_248),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_403),
.B(n_404),
.Y(n_438)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_355),
.Y(n_404)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_331),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_405),
.Y(n_445)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_242),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_410),
.B(n_413),
.Y(n_439)
);

OA22x2_ASAP7_75t_SL g411 ( 
.A1(n_312),
.A2(n_291),
.B1(n_240),
.B2(n_264),
.Y(n_411)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_411),
.A2(n_389),
.B(n_415),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_351),
.B(n_249),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_412),
.B(n_417),
.Y(n_455)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_344),
.B(n_289),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_416),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_347),
.A2(n_264),
.B1(n_251),
.B2(n_233),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_415),
.A2(n_419),
.B1(n_361),
.B2(n_338),
.Y(n_431)
);

BUFx12_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_311),
.B(n_233),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_324),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_337),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_368),
.A2(n_251),
.B1(n_276),
.B2(n_247),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_375),
.A2(n_348),
.B1(n_354),
.B2(n_313),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_422),
.B(n_426),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_375),
.A2(n_369),
.B1(n_329),
.B2(n_353),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_397),
.A2(n_350),
.B(n_361),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_437),
.B(n_450),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_431),
.B(n_458),
.Y(n_484)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_432),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_406),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_378),
.A2(n_369),
.B1(n_364),
.B2(n_333),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_435),
.A2(n_451),
.B1(n_457),
.B2(n_413),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_338),
.B(n_371),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_378),
.A2(n_353),
.B1(n_370),
.B2(n_332),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_444),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_392),
.B(n_400),
.C(n_398),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_453),
.C(n_456),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_359),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_447),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_383),
.B(n_327),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_449),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_411),
.A2(n_346),
.B1(n_333),
.B2(n_324),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_377),
.A2(n_326),
.B(n_341),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_407),
.B(n_377),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_411),
.A2(n_346),
.B1(n_340),
.B2(n_315),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_379),
.B(n_358),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_459),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_392),
.B(n_325),
.C(n_365),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_406),
.B(n_326),
.C(n_365),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_374),
.A2(n_395),
.B1(n_402),
.B2(n_388),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_408),
.A2(n_340),
.B1(n_362),
.B2(n_363),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_496),
.Y(n_528)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_454),
.Y(n_461)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_461),
.Y(n_498)
);

INVx8_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_462),
.B(n_473),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_420),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_463),
.B(n_471),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_414),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_485),
.C(n_456),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_427),
.B(n_416),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_466),
.B(n_469),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_468),
.A2(n_472),
.B(n_447),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_420),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_442),
.B(n_419),
.Y(n_473)
);

INVx13_ASAP7_75t_L g474 ( 
.A(n_445),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_474),
.Y(n_506)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_432),
.Y(n_475)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_475),
.Y(n_507)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_448),
.Y(n_476)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_476),
.Y(n_510)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_454),
.Y(n_477)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_477),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_405),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_479),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_446),
.B(n_403),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_425),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_483),
.B(n_492),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_394),
.C(n_401),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_451),
.A2(n_385),
.B1(n_376),
.B2(n_382),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_487),
.A2(n_493),
.B1(n_436),
.B2(n_458),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_441),
.B(n_408),
.Y(n_488)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_488),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_425),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_489),
.B(n_494),
.Y(n_532)
);

NOR2x1_ASAP7_75t_SL g490 ( 
.A(n_433),
.B(n_372),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_455),
.Y(n_521)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_441),
.Y(n_491)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_491),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_437),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_446),
.B(n_323),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_434),
.A2(n_385),
.B1(n_410),
.B2(n_408),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_495),
.A2(n_436),
.B1(n_421),
.B2(n_458),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_386),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_499),
.B(n_508),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_505),
.C(n_531),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_504),
.A2(n_526),
.B1(n_422),
.B2(n_404),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_467),
.B(n_465),
.C(n_496),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_480),
.Y(n_509)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_509),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_460),
.B(n_428),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_511),
.B(n_524),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_471),
.A2(n_421),
.B(n_439),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_512),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_482),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_516),
.B(n_520),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_518),
.A2(n_470),
.B1(n_515),
.B2(n_516),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_472),
.A2(n_458),
.B(n_431),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_519),
.B(n_523),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_482),
.Y(n_520)
);

XNOR2x1_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_481),
.Y(n_551)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_491),
.Y(n_522)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_522),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_488),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_467),
.B(n_480),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_484),
.A2(n_468),
.B(n_492),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_525),
.B(n_529),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_484),
.A2(n_470),
.B1(n_483),
.B2(n_463),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_476),
.B(n_430),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_527),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_486),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_484),
.A2(n_423),
.B1(n_434),
.B2(n_457),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_530),
.A2(n_486),
.B1(n_475),
.B2(n_464),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_485),
.B(n_438),
.C(n_444),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g534 ( 
.A(n_497),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_534),
.B(n_532),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_536),
.A2(n_538),
.B1(n_517),
.B2(n_514),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_505),
.B(n_438),
.C(n_495),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_539),
.B(n_545),
.C(n_546),
.Y(n_570)
);

XOR2x2_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_490),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_540),
.A2(n_551),
.B(n_562),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_521),
.A2(n_424),
.B1(n_462),
.B2(n_427),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_541),
.B(n_549),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_455),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_542),
.B(n_554),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_502),
.B(n_464),
.C(n_452),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_524),
.B(n_435),
.C(n_440),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_528),
.B(n_445),
.C(n_426),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_548),
.B(n_559),
.C(n_506),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_531),
.B(n_428),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_503),
.A2(n_423),
.B1(n_481),
.B2(n_449),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_552),
.B(n_506),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_527),
.B(n_459),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_555),
.A2(n_520),
.B1(n_510),
.B2(n_507),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_518),
.B(n_409),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_557),
.B(n_558),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_508),
.B(n_363),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_515),
.B(n_339),
.C(n_380),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_362),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_522),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_512),
.B(n_416),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_562),
.B(n_525),
.Y(n_567)
);

A2O1A1Ixp33_ASAP7_75t_SL g565 ( 
.A1(n_551),
.A2(n_513),
.B(n_501),
.C(n_519),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_565),
.A2(n_577),
.B(n_556),
.Y(n_598)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_535),
.Y(n_566)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_566),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_572),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_569),
.Y(n_601)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_543),
.Y(n_571)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_571),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_573),
.B(n_580),
.Y(n_595)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_561),
.Y(n_574)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_574),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_533),
.B(n_510),
.C(n_507),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_575),
.B(n_578),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_554),
.Y(n_576)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_576),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_553),
.A2(n_500),
.B1(n_501),
.B2(n_513),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_544),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_579),
.Y(n_588)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_559),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_547),
.B(n_530),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_581),
.B(n_582),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_547),
.B(n_542),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_583),
.A2(n_585),
.B1(n_537),
.B2(n_550),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_584),
.B(n_564),
.Y(n_593)
);

AO221x1_ASAP7_75t_L g586 ( 
.A1(n_585),
.A2(n_575),
.B1(n_568),
.B2(n_474),
.C(n_545),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_586),
.B(n_589),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_587),
.B(n_593),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_570),
.B(n_533),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_565),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_597),
.B(n_598),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_570),
.B(n_539),
.C(n_548),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_599),
.B(n_582),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_565),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_600),
.B(n_514),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_584),
.B(n_517),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_602),
.B(n_560),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_596),
.B(n_572),
.C(n_581),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_605),
.B(n_607),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_599),
.B(n_594),
.C(n_596),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_608),
.B(n_609),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_597),
.A2(n_576),
.B(n_565),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_604),
.B(n_564),
.C(n_563),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_610),
.B(n_611),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_604),
.B(n_563),
.C(n_546),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_587),
.B(n_567),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_614),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_613),
.B(n_619),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_588),
.B(n_540),
.C(n_557),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_595),
.B(n_588),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_617),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_601),
.B(n_558),
.C(n_499),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_618),
.Y(n_631)
);

OA21x2_ASAP7_75t_L g619 ( 
.A1(n_598),
.A2(n_498),
.B(n_477),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_593),
.B(n_498),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_621),
.B(n_602),
.C(n_603),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_622),
.B(n_625),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_605),
.B(n_601),
.C(n_603),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_616),
.A2(n_600),
.B1(n_595),
.B2(n_592),
.Y(n_627)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_627),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_606),
.A2(n_592),
.B1(n_612),
.B2(n_619),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_631),
.Y(n_639)
);

FAx1_ASAP7_75t_SL g629 ( 
.A(n_620),
.B(n_590),
.CI(n_591),
.CON(n_629),
.SN(n_629)
);

AOI31xp67_ASAP7_75t_L g640 ( 
.A1(n_629),
.A2(n_611),
.A3(n_331),
.B(n_339),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_619),
.A2(n_590),
.B1(n_591),
.B2(n_418),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_633),
.B(n_620),
.C(n_621),
.Y(n_637)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_637),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_632),
.B(n_610),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_638),
.B(n_639),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_640),
.A2(n_629),
.B(n_627),
.C(n_633),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_624),
.B(n_630),
.C(n_625),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_641),
.B(n_634),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_626),
.A2(n_345),
.B1(n_242),
.B2(n_247),
.Y(n_642)
);

OAI21xp33_ASAP7_75t_L g646 ( 
.A1(n_642),
.A2(n_643),
.B(n_253),
.Y(n_646)
);

AOI321xp33_ASAP7_75t_L g643 ( 
.A1(n_623),
.A2(n_257),
.A3(n_276),
.B1(n_345),
.B2(n_253),
.C(n_11),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_644),
.B(n_645),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_639),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_646),
.A2(n_647),
.B(n_634),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_SL g650 ( 
.A(n_648),
.B(n_636),
.C(n_635),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_650),
.A2(n_7),
.B(n_9),
.Y(n_654)
);

AOI31xp33_ASAP7_75t_L g653 ( 
.A1(n_651),
.A2(n_649),
.A3(n_622),
.B(n_257),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_653),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_655),
.B(n_652),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_656),
.B(n_654),
.Y(n_657)
);

AOI211xp5_ASAP7_75t_L g658 ( 
.A1(n_657),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_658)
);

XNOR2xp5_ASAP7_75t_L g659 ( 
.A(n_658),
.B(n_11),
.Y(n_659)
);


endmodule