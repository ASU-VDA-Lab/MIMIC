module fake_jpeg_4703_n_297 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_38),
.B(n_23),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_40),
.Y(n_73)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_20),
.B(n_0),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_55),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_60),
.B1(n_30),
.B2(n_19),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_21),
.B1(n_26),
.B2(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_53),
.A2(n_54),
.B1(n_81),
.B2(n_17),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_21),
.B1(n_25),
.B2(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_56),
.B(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_62),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_26),
.B1(n_33),
.B2(n_22),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_26),
.Y(n_71)
);

NOR2x1_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_97),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_82),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_39),
.A2(n_17),
.B(n_12),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_92),
.B(n_95),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_43),
.B(n_29),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_38),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_34),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_43),
.B(n_23),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_98),
.B1(n_18),
.B2(n_30),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_38),
.A2(n_24),
.B(n_33),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_46),
.A2(n_34),
.B1(n_30),
.B2(n_19),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_111),
.B1(n_115),
.B2(n_78),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_120),
.B1(n_85),
.B2(n_73),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_18),
.B1(n_22),
.B2(n_14),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g112 ( 
.A(n_60),
.B(n_71),
.Y(n_112)
);

XNOR2x1_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_33),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_22),
.B1(n_8),
.B2(n_9),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_9),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_52),
.A2(n_33),
.B1(n_16),
.B2(n_17),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_72),
.A2(n_16),
.B1(n_33),
.B2(n_24),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_72),
.B1(n_78),
.B2(n_67),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_71),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_129),
.A2(n_161),
.B(n_107),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_100),
.B(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_130),
.B(n_153),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_77),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_142),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_133),
.A2(n_141),
.B1(n_145),
.B2(n_147),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_134),
.B(n_143),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_128),
.B(n_16),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_90),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_59),
.C(n_77),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_155),
.C(n_159),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_138),
.A2(n_148),
.B1(n_118),
.B2(n_123),
.Y(n_179)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_67),
.B1(n_69),
.B2(n_64),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_79),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_105),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_75),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_152),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_69),
.B1(n_57),
.B2(n_86),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_150),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_83),
.B1(n_57),
.B2(n_51),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_66),
.A3(n_73),
.B1(n_84),
.B2(n_33),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_151),
.Y(n_184)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_50),
.B1(n_94),
.B2(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_75),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_88),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_123),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_63),
.B1(n_73),
.B2(n_33),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_125),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_157),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_61),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_104),
.B(n_8),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_104),
.A2(n_117),
.B1(n_101),
.B2(n_108),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_8),
.C(n_1),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_88),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_16),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

AOI32xp33_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_122),
.A3(n_121),
.B1(n_107),
.B2(n_128),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_166),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_168),
.C1(n_183),
.C2(n_174),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_167),
.A2(n_0),
.B(n_1),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_116),
.B1(n_96),
.B2(n_126),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_141),
.B1(n_140),
.B2(n_138),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_170),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_131),
.A2(n_126),
.B1(n_108),
.B2(n_118),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_96),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_198),
.C(n_145),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_178),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_179),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_180),
.B(n_181),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_142),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_192),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_63),
.B1(n_24),
.B2(n_2),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_133),
.B1(n_153),
.B2(n_146),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_195),
.Y(n_200)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_197),
.B(n_2),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_132),
.B(n_24),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_203),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_SL g239 ( 
.A1(n_202),
.A2(n_187),
.B(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_208),
.C(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_130),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_205),
.B(n_219),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_149),
.C(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_218),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_140),
.B(n_156),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_211),
.A2(n_214),
.B(n_205),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_157),
.C(n_24),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_24),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_217),
.C(n_191),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_214),
.A2(n_225),
.B(n_165),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_1),
.C(n_2),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_3),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_178),
.B(n_3),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_221),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_193),
.B1(n_181),
.B2(n_184),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_202),
.B1(n_218),
.B2(n_199),
.Y(n_247)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_184),
.B(n_183),
.C(n_204),
.D(n_200),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_240),
.B(n_243),
.Y(n_261)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_200),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_231),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_213),
.C(n_212),
.Y(n_249)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_238),
.Y(n_248)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_239),
.A2(n_210),
.B1(n_187),
.B2(n_220),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_245),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_183),
.B(n_180),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

OAI211xp5_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_243),
.B(n_239),
.C(n_235),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_250),
.C(n_251),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_233),
.C(n_227),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_203),
.C(n_217),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_253),
.A2(n_235),
.B1(n_246),
.B2(n_234),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_186),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_259),
.C(n_232),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_236),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_224),
.B1(n_187),
.B2(n_215),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_238),
.B1(n_242),
.B2(n_236),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

NAND4xp25_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.C(n_258),
.D(n_253),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_249),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_245),
.B1(n_246),
.B2(n_232),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_271),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_169),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_273),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_242),
.C(n_226),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_251),
.C(n_247),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_175),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_263),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_281),
.B(n_266),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_262),
.B(n_252),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_237),
.B(n_248),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_260),
.B(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_255),
.C(n_259),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_SL g286 ( 
.A1(n_282),
.A2(n_265),
.B(n_269),
.C(n_229),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_278),
.Y(n_283)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_186),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_276),
.B(n_280),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_260),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_294),
.B(n_290),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_292),
.B(n_281),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_274),
.C(n_185),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_241),
.Y(n_297)
);


endmodule