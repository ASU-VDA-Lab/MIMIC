module fake_jpeg_8191_n_33 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_1),
.Y(n_18)
);

AND2x6_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_9),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_19),
.A2(n_21),
.B(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_2),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_4),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_4),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_10),
.B1(n_14),
.B2(n_7),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.C(n_25),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_21),
.A2(n_11),
.B1(n_13),
.B2(n_8),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_5),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_25),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_23),
.B1(n_27),
.B2(n_29),
.Y(n_33)
);


endmodule