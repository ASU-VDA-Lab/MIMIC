module fake_jpeg_17663_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_8),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OR2x2_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_0),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_11),
.B1(n_16),
.B2(n_13),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_13),
.B1(n_15),
.B2(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_15),
.B1(n_13),
.B2(n_18),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_46),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_15),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_14),
.B(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

OAI32xp33_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_22),
.A3(n_12),
.B1(n_14),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_18),
.B1(n_19),
.B2(n_14),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_1),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_55),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_57),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_45),
.C(n_41),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_44),
.C(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_28),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_55),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_39),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_69),
.C(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_44),
.B(n_37),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_57),
.B(n_49),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_28),
.B1(n_35),
.B2(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_35),
.B1(n_24),
.B2(n_42),
.Y(n_71)
);

OA21x2_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_33),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_53),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_2),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_82),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_78),
.B1(n_80),
.B2(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_48),
.B1(n_52),
.B2(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_84),
.B(n_52),
.Y(n_86)
);

XNOR2x2_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_50),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_69),
.C(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_90),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.C(n_92),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_65),
.C(n_62),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_85),
.B(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_72),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_75),
.C(n_5),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_95),
.B(n_82),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_83),
.B(n_76),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_80),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_96),
.C(n_82),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_84),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_99),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_4),
.B(n_5),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_100),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_101),
.Y(n_103)
);

NOR2xp67_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_4),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_102),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_107),
.B(n_108),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_8),
.C(n_105),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_109),
.Y(n_110)
);


endmodule