module fake_jpeg_1739_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_66),
.Y(n_69)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_45),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_46),
.B1(n_49),
.B2(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_55),
.B1(n_53),
.B2(n_51),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_60),
.B1(n_46),
.B2(n_49),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_59),
.B1(n_1),
.B2(n_3),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_45),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_96),
.B1(n_4),
.B2(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_90),
.Y(n_112)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_57),
.B1(n_59),
.B2(n_48),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_95),
.B(n_9),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_9),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_19),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_57),
.B1(n_59),
.B2(n_3),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_69),
.B1(n_76),
.B2(n_23),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_76),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_43),
.B1(n_29),
.B2(n_32),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_7),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_11),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_10),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_30),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_11),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_95),
.B(n_12),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_34),
.B(n_36),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_129),
.B1(n_120),
.B2(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_17),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_18),
.B1(n_22),
.B2(n_26),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_27),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_106),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_28),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_136),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_97),
.C(n_35),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_37),
.Y(n_154)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_147),
.B1(n_115),
.B2(n_116),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_123),
.B1(n_127),
.B2(n_138),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_154),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_123),
.B1(n_127),
.B2(n_40),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_139),
.B(n_140),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_146),
.B(n_147),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_136),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_150),
.B(n_148),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_162),
.C(n_157),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_155),
.B(n_142),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.C(n_154),
.Y(n_165)
);

AO21x2_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_135),
.B(n_41),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_157),
.B(n_134),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_38),
.Y(n_169)
);


endmodule