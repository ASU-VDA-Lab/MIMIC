module fake_jpeg_14675_n_214 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx9p33_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_1),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_17),
.C(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_1),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_15),
.B1(n_19),
.B2(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_53),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_19),
.B1(n_21),
.B2(n_18),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_37),
.B1(n_19),
.B2(n_21),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_79),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_67),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_78),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_39),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_82),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_20),
.B(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_104),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_57),
.B1(n_43),
.B2(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_51),
.B1(n_62),
.B2(n_72),
.Y(n_115)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_21),
.B(n_34),
.C(n_56),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_62),
.B(n_46),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_56),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_67),
.B(n_38),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_99),
.C(n_50),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_76),
.CI(n_63),
.CON(n_98),
.SN(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_65),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_17),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_27),
.B1(n_51),
.B2(n_18),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_101),
.B1(n_102),
.B2(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_116),
.B1(n_89),
.B2(n_66),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_122),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_80),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_98),
.C(n_103),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_25),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_138),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_127),
.B1(n_125),
.B2(n_118),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_92),
.C(n_88),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_131),
.C(n_135),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_92),
.C(n_102),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_133),
.B1(n_115),
.B2(n_117),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_97),
.B1(n_72),
.B2(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_25),
.Y(n_158)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_106),
.C(n_107),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_109),
.B(n_106),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_157),
.B(n_134),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_109),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_151),
.C(n_131),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_154),
.B1(n_158),
.B2(n_140),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_152),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_105),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_155),
.B(n_159),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_118),
.B1(n_111),
.B2(n_112),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_113),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_110),
.B(n_114),
.C(n_49),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_66),
.B1(n_69),
.B2(n_35),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_143),
.B1(n_134),
.B2(n_31),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_69),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_160),
.A2(n_149),
.B(n_148),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_130),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_164),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_167),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_133),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_164),
.B1(n_169),
.B2(n_166),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_166),
.A2(n_31),
.B(n_3),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_126),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_169),
.B(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_47),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_172),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_157),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_47),
.C(n_31),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_28),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_181),
.B(n_171),
.C(n_173),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_177),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_10),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_178),
.B(n_12),
.Y(n_193)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

AND2x4_ASAP7_75t_SL g181 ( 
.A(n_172),
.B(n_2),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_167),
.B1(n_163),
.B2(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_30),
.B(n_5),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_180),
.C(n_185),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_181),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_14),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_193),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_177),
.B(n_12),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_188),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_189),
.A2(n_175),
.B(n_185),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_198),
.B(n_192),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_190),
.A2(n_3),
.B(n_4),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_186),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_201),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_195),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_30),
.C(n_8),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_209),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_202),
.A2(n_192),
.B(n_200),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_208),
.A2(n_210),
.B(n_7),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_30),
.B(n_8),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_212),
.A2(n_7),
.B(n_35),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_211),
.Y(n_214)
);


endmodule