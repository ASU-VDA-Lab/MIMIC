module fake_jpeg_15827_n_121 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_31),
.B1(n_15),
.B2(n_26),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_49),
.B1(n_30),
.B2(n_14),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_31),
.B1(n_26),
.B2(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_29),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_18),
.B1(n_31),
.B2(n_23),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_60),
.B1(n_22),
.B2(n_20),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_23),
.B1(n_22),
.B2(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_69),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_32),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_30),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_33),
.C(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_73),
.Y(n_76)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_72),
.B(n_56),
.C(n_53),
.D(n_62),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_78),
.C(n_69),
.Y(n_96)
);

NOR4xp25_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_56),
.C(n_49),
.D(n_52),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_51),
.B1(n_50),
.B2(n_74),
.Y(n_79)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_75),
.B(n_61),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_64),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_85),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_30),
.B(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_87),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_57),
.C(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_24),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_96),
.B(n_92),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_63),
.B(n_64),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_77),
.C(n_76),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_99),
.C(n_21),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_83),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_85),
.C(n_1),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_101),
.B(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_7),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

OAI321xp33_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_95),
.A3(n_94),
.B1(n_93),
.B2(n_88),
.C(n_21),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_107),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_14),
.C(n_13),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_103),
.B(n_8),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_109),
.B(n_112),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_6),
.B(n_11),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_109),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_115),
.Y(n_119)
);

AOI221xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_120),
.Y(n_121)
);


endmodule