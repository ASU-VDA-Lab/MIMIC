module fake_jpeg_8148_n_279 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_21),
.B1(n_30),
.B2(n_34),
.Y(n_50)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_21),
.B1(n_27),
.B2(n_30),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_41),
.B1(n_37),
.B2(n_35),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_52),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_51),
.B(n_18),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_27),
.B1(n_34),
.B2(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_SL g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_57),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_29),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_35),
.B1(n_62),
.B2(n_42),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_74),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_81),
.B(n_88),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_26),
.B(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_76),
.B(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_80),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_85),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_17),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_27),
.B1(n_18),
.B2(n_37),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_41),
.B(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_0),
.B(n_1),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_75),
.Y(n_104)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_42),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_103),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_111),
.B1(n_71),
.B2(n_93),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_57),
.B1(n_35),
.B2(n_37),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_118),
.B1(n_69),
.B2(n_72),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_58),
.B(n_63),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_105),
.B(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_70),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_42),
.B(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_38),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_28),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_31),
.B(n_28),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_64),
.B1(n_55),
.B2(n_54),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_49),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_131),
.B(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_124),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_32),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_126),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_98),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_82),
.B1(n_73),
.B2(n_90),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_147),
.B1(n_108),
.B2(n_80),
.Y(n_152)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_110),
.B1(n_117),
.B2(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_137),
.B(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_66),
.B(n_78),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_76),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_95),
.C(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_84),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_73),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_91),
.B(n_83),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_87),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_109),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_148),
.A2(n_152),
.B1(n_145),
.B2(n_129),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_123),
.B(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_150),
.B(n_171),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_104),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_159),
.B(n_162),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_158),
.C(n_164),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_95),
.B1(n_112),
.B2(n_102),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_168),
.B1(n_147),
.B2(n_133),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_109),
.C(n_71),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_115),
.B(n_32),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_122),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_137),
.B(n_131),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_107),
.C(n_102),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_102),
.B(n_107),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_173),
.B(n_174),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_112),
.B1(n_97),
.B2(n_49),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_107),
.C(n_97),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_130),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_22),
.B(n_20),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_97),
.B(n_22),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_179),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_180),
.B(n_189),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_188),
.B1(n_171),
.B2(n_38),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

AO21x2_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_126),
.B(n_120),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_185),
.A2(n_193),
.B1(n_195),
.B2(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_158),
.C(n_153),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_138),
.C(n_144),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_121),
.B1(n_20),
.B2(n_23),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_196),
.B1(n_198),
.B2(n_148),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_16),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_38),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_49),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_204),
.C(n_212),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_161),
.C(n_153),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_168),
.B1(n_167),
.B2(n_159),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_166),
.B1(n_173),
.B2(n_149),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_149),
.C(n_156),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_155),
.C(n_38),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_216),
.C(n_218),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_155),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_221),
.B1(n_3),
.B2(n_4),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_23),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_23),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_209),
.B(n_182),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_5),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_185),
.B(n_199),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_225),
.A2(n_226),
.B(n_227),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_211),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_213),
.A2(n_191),
.B(n_184),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_184),
.B(n_193),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_203),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_183),
.B1(n_200),
.B2(n_3),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_201),
.B1(n_220),
.B2(n_207),
.Y(n_239)
);

HAxp5_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_1),
.CON(n_235),
.SN(n_235)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_7),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_3),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_207),
.B1(n_5),
.B2(n_6),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_242),
.B1(n_248),
.B2(n_236),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_215),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_246),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_212),
.C(n_5),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_247),
.C(n_224),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_231),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_234),
.B(n_237),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_229),
.B(n_231),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_253),
.B(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_252),
.B(n_254),
.Y(n_266)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_225),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_241),
.A2(n_230),
.B1(n_228),
.B2(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_232),
.B1(n_227),
.B2(n_233),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_247),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_10),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_265),
.B(n_258),
.C(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_263),
.C(n_257),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_222),
.B(n_233),
.Y(n_263)
);

NOR3xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_8),
.C(n_9),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_10),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_271),
.B1(n_11),
.B2(n_12),
.Y(n_274)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_271),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_275),
.C(n_272),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_11),
.Y(n_279)
);


endmodule