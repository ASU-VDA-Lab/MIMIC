module fake_jpeg_31315_n_526 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_58),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_53),
.B(n_86),
.Y(n_140)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_87),
.Y(n_120)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_16),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_28),
.Y(n_89)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_50),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_100),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_36),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_19),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_148),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_47),
.B1(n_50),
.B2(n_49),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_123),
.A2(n_135),
.B1(n_39),
.B2(n_41),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_141),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_99),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_153),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_68),
.A2(n_51),
.B(n_24),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_139),
.A2(n_25),
.B(n_43),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_19),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_36),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_143),
.B(n_144),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_55),
.B(n_27),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_54),
.B(n_20),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_63),
.B(n_20),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_13),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_59),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_56),
.A2(n_51),
.B1(n_43),
.B2(n_35),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_39),
.B1(n_25),
.B2(n_35),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_88),
.B(n_49),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_32),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_64),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_76),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_27),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_168),
.B(n_196),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_169),
.B(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_171),
.Y(n_267)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_174),
.A2(n_178),
.B1(n_165),
.B2(n_65),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_105),
.A2(n_82),
.B1(n_97),
.B2(n_91),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_175),
.A2(n_182),
.B1(n_184),
.B2(n_188),
.Y(n_243)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_214),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_118),
.A2(n_97),
.B1(n_83),
.B2(n_88),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_85),
.B1(n_79),
.B2(n_77),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_164),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_186),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_137),
.A2(n_73),
.B1(n_72),
.B2(n_71),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_190),
.Y(n_254)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_139),
.A2(n_60),
.B1(n_10),
.B2(n_16),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_194),
.B(n_213),
.Y(n_252)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_120),
.B(n_9),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_128),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_197),
.B(n_198),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_10),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_199),
.Y(n_266)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_200),
.Y(n_268)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_204),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_141),
.B(n_10),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_202),
.B(n_205),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_119),
.B(n_15),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_207),
.Y(n_258)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_208),
.B(n_211),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_125),
.B(n_15),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_209),
.B(n_210),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_110),
.B(n_15),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

BUFx8_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_122),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_215),
.B(n_217),
.Y(n_259)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_132),
.B(n_14),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_126),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_223),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_13),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_221),
.B(n_222),
.Y(n_270)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_152),
.C(n_130),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_226),
.B(n_220),
.C(n_219),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_109),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_230),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_167),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_167),
.A2(n_160),
.B1(n_157),
.B2(n_109),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_237),
.B(n_250),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_142),
.B(n_130),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_242),
.A2(n_152),
.B(n_175),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_115),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_184),
.A2(n_135),
.B1(n_134),
.B2(n_147),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_165),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_253),
.A2(n_242),
.B1(n_262),
.B2(n_191),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_179),
.B(n_145),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_262),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_188),
.A2(n_66),
.B1(n_61),
.B2(n_147),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_265),
.B1(n_203),
.B2(n_212),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_214),
.B(n_116),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_182),
.A2(n_116),
.B1(n_134),
.B2(n_145),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_256),
.B(n_230),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_271),
.B(n_273),
.Y(n_335)
);

AO22x1_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_252),
.B1(n_253),
.B2(n_261),
.Y(n_272)
);

AO21x2_ASAP7_75t_SL g321 ( 
.A1(n_272),
.A2(n_277),
.B(n_244),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_255),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_60),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_264),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_195),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_282),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_234),
.B(n_232),
.C(n_227),
.Y(n_277)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_280),
.A2(n_239),
.B(n_235),
.Y(n_333)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_281),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_259),
.B(n_241),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_291),
.B1(n_296),
.B2(n_244),
.Y(n_320)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_285),
.Y(n_345)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_286),
.B(n_287),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_206),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_226),
.B(n_216),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_292),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_290),
.B(n_298),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_246),
.B(n_270),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_228),
.B(n_211),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_293),
.B(n_295),
.Y(n_323)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_207),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_265),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_186),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_231),
.B(n_185),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_299),
.B(n_300),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_159),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_303),
.Y(n_326)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_305),
.Y(n_336)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_224),
.Y(n_305)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_309),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_243),
.B(n_161),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_236),
.Y(n_309)
);

INVx5_ASAP7_75t_SL g310 ( 
.A(n_224),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_310),
.A2(n_232),
.B1(n_247),
.B2(n_263),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_248),
.B(n_13),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_11),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_264),
.B(n_142),
.C(n_161),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_233),
.C(n_239),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_277),
.A2(n_264),
.B(n_244),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_313),
.A2(n_330),
.B(n_278),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_SL g316 ( 
.A(n_272),
.B(n_280),
.C(n_271),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_316),
.A2(n_312),
.B(n_292),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_333),
.B(n_296),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_337),
.C(n_289),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_320),
.A2(n_329),
.B1(n_331),
.B2(n_349),
.Y(n_376)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_272),
.A2(n_225),
.B1(n_229),
.B2(n_269),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_322),
.A2(n_328),
.B1(n_332),
.B2(n_340),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_346),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_276),
.A2(n_245),
.B1(n_171),
.B2(n_189),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_291),
.A2(n_225),
.B1(n_247),
.B2(n_229),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_283),
.A2(n_224),
.B(n_263),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_284),
.A2(n_308),
.B1(n_296),
.B2(n_276),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_283),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_288),
.A2(n_213),
.B1(n_192),
.B2(n_235),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_343),
.B(n_311),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_138),
.C(n_146),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_308),
.A2(n_267),
.B1(n_133),
.B2(n_146),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_278),
.Y(n_350)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_351),
.A2(n_359),
.B(n_365),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_346),
.C(n_337),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_371),
.Y(n_388)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_356),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_342),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_357),
.B(n_360),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_273),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_364),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_318),
.B(n_304),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_318),
.B(n_290),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_343),
.Y(n_406)
);

AOI322xp5_ASAP7_75t_L g362 ( 
.A1(n_316),
.A2(n_282),
.A3(n_274),
.B1(n_279),
.B2(n_306),
.C1(n_301),
.C2(n_294),
.Y(n_362)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_362),
.B(n_373),
.C(n_8),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_326),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_363),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_305),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_348),
.A2(n_309),
.B(n_307),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_285),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_370),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_314),
.Y(n_367)
);

INVx11_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_320),
.A2(n_281),
.B1(n_303),
.B2(n_302),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_368),
.A2(n_322),
.B1(n_348),
.B2(n_321),
.Y(n_394)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_286),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_313),
.A2(n_310),
.B(n_133),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_339),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_334),
.Y(n_401)
);

A2O1A1O1Ixp25_ASAP7_75t_L g373 ( 
.A1(n_330),
.A2(n_321),
.B(n_325),
.C(n_319),
.D(n_339),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_310),
.Y(n_375)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_345),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_379),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_340),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_380),
.Y(n_404)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_381),
.Y(n_411)
);

NAND2x1_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_321),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_386),
.B(n_375),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_351),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_397),
.C(n_398),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_324),
.C(n_333),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_331),
.C(n_329),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_376),
.A2(n_334),
.B1(n_315),
.B2(n_349),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_381),
.Y(n_403)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_403),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_406),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_342),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_407),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_378),
.A2(n_138),
.B1(n_1),
.B2(n_2),
.Y(n_408)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_408),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_376),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_409),
.A2(n_371),
.B(n_361),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_356),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_400),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_416),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_415),
.A2(n_426),
.B1(n_433),
.B2(n_394),
.Y(n_441)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_382),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_422),
.Y(n_457)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_421),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_359),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_354),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_423),
.B(n_432),
.Y(n_442)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_393),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_427),
.Y(n_456)
);

XNOR2x2_ASAP7_75t_SL g458 ( 
.A(n_425),
.B(n_386),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_388),
.A2(n_377),
.B1(n_352),
.B2(n_372),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_363),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_435),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_360),
.C(n_355),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_365),
.C(n_410),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_388),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_395),
.A2(n_352),
.B1(n_380),
.B2(n_373),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_383),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_384),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_436),
.B(n_405),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_390),
.Y(n_439)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_439),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_445),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_428),
.A2(n_395),
.B1(n_384),
.B2(n_404),
.Y(n_444)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_444),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_388),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_446),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_428),
.A2(n_404),
.B1(n_399),
.B2(n_378),
.Y(n_449)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_450),
.B(n_459),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_415),
.A2(n_389),
.B1(n_391),
.B2(n_386),
.Y(n_451)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_451),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_391),
.C(n_350),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_454),
.C(n_418),
.Y(n_471)
);

FAx1_ASAP7_75t_SL g453 ( 
.A(n_432),
.B(n_406),
.CI(n_389),
.CON(n_453),
.SN(n_453)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_410),
.C(n_402),
.Y(n_454)
);

AO22x1_ASAP7_75t_L g467 ( 
.A1(n_458),
.A2(n_425),
.B1(n_426),
.B2(n_431),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_430),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_454),
.B(n_437),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_464),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_440),
.B(n_390),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_467),
.B(n_441),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_468),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_453),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_470),
.B(n_445),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_450),
.C(n_457),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_456),
.A2(n_433),
.B(n_427),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_472),
.A2(n_474),
.B(n_444),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_456),
.A2(n_438),
.B1(n_414),
.B2(n_417),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_451),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_458),
.A2(n_414),
.B(n_424),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_477),
.B(n_489),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_471),
.B(n_452),
.C(n_457),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_478),
.B(n_479),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_409),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_482),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_484),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_442),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_422),
.C(n_442),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_485),
.B(n_488),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_474),
.A2(n_443),
.B(n_455),
.Y(n_486)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_486),
.Y(n_494)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_487),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_449),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_448),
.C(n_421),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_467),
.A2(n_419),
.B(n_385),
.Y(n_491)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_491),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_482),
.A2(n_476),
.B(n_466),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_495),
.B(n_499),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_460),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_473),
.B(n_469),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_489),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_479),
.C(n_487),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_508),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_493),
.B(n_465),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_507),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_502),
.B(n_484),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_480),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_510),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_490),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_501),
.B(n_369),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_511),
.A2(n_393),
.B(n_494),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_512),
.A2(n_513),
.B(n_500),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_504),
.A2(n_496),
.B(n_499),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_517),
.A2(n_514),
.B1(n_374),
.B2(n_434),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_505),
.C(n_379),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_SL g521 ( 
.A(n_518),
.B(n_519),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_516),
.A2(n_508),
.B(n_509),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_520),
.A2(n_411),
.B(n_434),
.Y(n_522)
);

AOI322xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_521),
.A3(n_357),
.B1(n_403),
.B2(n_411),
.C1(n_6),
.C2(n_0),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_1),
.C(n_4),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_4),
.C(n_5),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_7),
.Y(n_526)
);


endmodule