module fake_jpeg_17297_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_71),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_65),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_62),
.B1(n_56),
.B2(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_84),
.B1(n_89),
.B2(n_1),
.Y(n_111)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_91),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_57),
.B1(n_58),
.B2(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_47),
.B1(n_49),
.B2(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_56),
.C(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_58),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_96),
.B(n_103),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_66),
.B(n_55),
.C(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_59),
.B1(n_51),
.B2(n_3),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_121)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_20),
.B1(n_45),
.B2(n_43),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_122),
.B1(n_123),
.B2(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_1),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_4),
.Y(n_131)
);

NAND2x1_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_2),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_95),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_102),
.B1(n_107),
.B2(n_108),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_129),
.B(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_118),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_122),
.C(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_122),
.B1(n_121),
.B2(n_131),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_141),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_115),
.C(n_124),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_32),
.B(n_46),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_120),
.B1(n_116),
.B2(n_26),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_130),
.C(n_31),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_134),
.B1(n_116),
.B2(n_120),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_144),
.B1(n_5),
.B2(n_6),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_34),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_21),
.B1(n_41),
.B2(n_40),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_18),
.C(n_22),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_147),
.B(n_149),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_145),
.C(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_150),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_13),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_12),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_35),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_11),
.B(n_39),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_38),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_98),
.C(n_93),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_36),
.B(n_118),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_6),
.B(n_8),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_8),
.B(n_9),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_9),
.C(n_10),
.Y(n_164)
);


endmodule