module real_jpeg_22304_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_249;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_211;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_0),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_0),
.A2(n_32),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_0),
.A2(n_32),
.B1(n_68),
.B2(n_69),
.Y(n_110)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_3),
.B(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_3),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_3),
.B(n_31),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_68),
.B1(n_69),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_5),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_80),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_80),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_80),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_6),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_42),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_26),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_8),
.A2(n_68),
.B(n_70),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_8),
.B(n_71),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_8),
.A2(n_10),
.B(n_25),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_8),
.B(n_141),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_8),
.A2(n_52),
.B(n_55),
.C(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_73),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_9),
.A2(n_68),
.B(n_72),
.C(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_35),
.B(n_38),
.C(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_10),
.B(n_38),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_123),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_122),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_104),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_16),
.B(n_104),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_81),
.C(n_90),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_17),
.A2(n_18),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.C(n_63),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_19),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_20),
.B(n_33),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_21),
.B(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_22),
.B(n_28),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_23),
.A2(n_29),
.B(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_24),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_26),
.A2(n_36),
.B(n_39),
.C(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_26),
.B(n_34),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_26),
.B(n_94),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_26),
.A2(n_38),
.B(n_57),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_27),
.A2(n_30),
.B(n_131),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_27),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_28),
.B(n_183),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_29),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B(n_43),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_34),
.A2(n_96),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_35),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_35),
.B(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_35),
.B(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_37),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_39),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_43),
.B(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_45),
.B(n_84),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_45),
.B(n_191),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_47),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_58),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_50),
.A2(n_60),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_50),
.B(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_51),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_54),
.B(n_55),
.C(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_52),
.B(n_73),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_53),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_54),
.A2(n_61),
.B(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_58),
.B(n_140),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_59),
.B(n_141),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_61),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_72),
.B(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_76),
.Y(n_112)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_72),
.B(n_79),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_108),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_76),
.B(n_110),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_81),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B(n_89),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_83),
.B(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_140),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_105),
.CI(n_121),
.CON(n_104),
.SN(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_93),
.A2(n_99),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_93),
.B(n_218),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_93),
.A2(n_95),
.B1(n_99),
.B2(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_95),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_97),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_101),
.B(n_103),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_104),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_113),
.B2(n_114),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_136),
.C(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_116),
.B1(n_138),
.B2(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_280),
.B(n_286),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_268),
.B(n_279),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_174),
.B(n_250),
.C(n_267),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_163),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_127),
.B(n_163),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_143),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_129),
.B(n_135),
.C(n_143),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_130),
.B(n_133),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_132),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_137),
.B(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_153),
.B1(n_154),
.B2(n_162),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_152),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_145),
.B(n_152),
.C(n_153),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_164),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_166),
.Y(n_247)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_169),
.B(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_170),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_182),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_249),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_243),
.B(n_248),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_229),
.B(n_242),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_214),
.B(n_228),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_203),
.B(n_213),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_192),
.B(n_202),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_184),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_188),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_197),
.B(n_201),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_210),
.C(n_212),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_216),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_221),
.B1(n_222),
.B2(n_227),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_217),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_226),
.C(n_227),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_231),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_238),
.C(n_241),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_238),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_239),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_252),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_265),
.B2(n_266),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_256),
.C(n_266),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_270),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_278),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_276),
.C(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);


endmodule