module fake_jpeg_25235_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_22),
.B1(n_31),
.B2(n_24),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_42),
.C(n_40),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_22),
.B1(n_28),
.B2(n_30),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_51),
.B1(n_20),
.B2(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_53),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_19),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_31),
.B1(n_33),
.B2(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_31),
.B1(n_21),
.B2(n_27),
.Y(n_70)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_39),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_40),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_76),
.B1(n_85),
.B2(n_38),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_73),
.B(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_1),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_1),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_19),
.B1(n_33),
.B2(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_26),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_42),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_25),
.B1(n_33),
.B2(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_113),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_100),
.B1(n_20),
.B2(n_21),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_106),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_49),
.B1(n_56),
.B2(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_82),
.B1(n_69),
.B2(n_49),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_88),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_80),
.B1(n_84),
.B2(n_88),
.Y(n_130)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_94),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_29),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_66),
.B(n_74),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_124),
.B1(n_129),
.B2(n_134),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_123),
.B(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_97),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_100),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_127),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_75),
.B(n_66),
.C(n_67),
.D(n_81),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_75),
.B1(n_64),
.B2(n_84),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_67),
.C(n_16),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_132),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_84),
.B1(n_58),
.B2(n_60),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_83),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_106),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_108),
.C(n_95),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_148),
.C(n_153),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_154),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_93),
.B1(n_86),
.B2(n_88),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_157),
.B1(n_162),
.B2(n_24),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_90),
.C(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_151),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_90),
.B1(n_101),
.B2(n_105),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_126),
.B1(n_137),
.B2(n_78),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_102),
.C(n_59),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_55),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_102),
.C(n_59),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_101),
.B1(n_105),
.B2(n_80),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_55),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_133),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_78),
.B1(n_72),
.B2(n_27),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_165),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_131),
.B1(n_129),
.B2(n_120),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_178),
.B1(n_141),
.B2(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_170),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_18),
.C(n_34),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_168),
.B(n_175),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_125),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_171),
.B(n_152),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_176),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_136),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_125),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_159),
.B1(n_158),
.B2(n_155),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_24),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_181),
.C(n_153),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_24),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_186),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_198),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_157),
.B1(n_162),
.B2(n_159),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_182),
.B(n_173),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_197),
.B(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_141),
.B1(n_140),
.B2(n_158),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_154),
.B1(n_145),
.B2(n_34),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_175),
.A2(n_18),
.B(n_34),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_204),
.B(n_210),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_174),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_205),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_182),
.C(n_173),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_191),
.C(n_186),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_192),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_181),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_194),
.C(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_185),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_3),
.B(n_4),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_16),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_220),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_193),
.C(n_187),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_190),
.B1(n_195),
.B2(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_221),
.B(n_222),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_198),
.C(n_7),
.Y(n_222)
);

OA21x2_ASAP7_75t_SL g224 ( 
.A1(n_218),
.A2(n_209),
.B(n_200),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_230),
.B(n_217),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_200),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_228),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_205),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_206),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_6),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_235),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_227),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_8),
.Y(n_236)
);

NAND4xp25_ASAP7_75t_SL g238 ( 
.A(n_236),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_238)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_10),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_236),
.A3(n_232),
.B1(n_11),
.B2(n_13),
.C1(n_9),
.C2(n_15),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_243),
.C(n_11),
.Y(n_244)
);

OAI211xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_14),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_245),
.Y(n_248)
);


endmodule