module fake_jpeg_857_n_187 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_66),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_63),
.B1(n_46),
.B2(n_60),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_93),
.B1(n_77),
.B2(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_92),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_48),
.C(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_60),
.B1(n_58),
.B2(n_52),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_52),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_58),
.B1(n_48),
.B2(n_56),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_53),
.B(n_55),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_3),
.B(n_4),
.Y(n_128)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_109),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

AOI31xp33_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_61),
.A3(n_54),
.B(n_51),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_51),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_55),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_104),
.C(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_114),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_93),
.B1(n_95),
.B2(n_57),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_133),
.B1(n_128),
.B2(n_119),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_132),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_44),
.B1(n_61),
.B2(n_20),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_130),
.B1(n_25),
.B2(n_24),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_125),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_0),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_43),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_134),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_114),
.B(n_112),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_42),
.B1(n_41),
.B2(n_39),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

BUFx4f_ASAP7_75t_SL g156 ( 
.A(n_142),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_105),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_10),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_100),
.B(n_32),
.C(n_31),
.D(n_28),
.Y(n_144)
);

OA21x2_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_152),
.B(n_9),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_6),
.C(n_8),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_150),
.B1(n_18),
.B2(n_11),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_133),
.B1(n_118),
.B2(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_5),
.Y(n_152)
);

AO32x1_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_12),
.C(n_13),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_157),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_23),
.C(n_21),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_159),
.C(n_160),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_150),
.B1(n_147),
.B2(n_144),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_10),
.C(n_12),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_148),
.C(n_143),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_151),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_169),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_161),
.C(n_162),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_178),
.B1(n_153),
.B2(n_14),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_167),
.B(n_163),
.CI(n_156),
.CON(n_178),
.SN(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_171),
.C(n_163),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_180),
.B(n_181),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_173),
.C(n_166),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_177),
.B(n_178),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_13),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_15),
.C(n_16),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_15),
.C(n_16),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_17),
.Y(n_187)
);


endmodule