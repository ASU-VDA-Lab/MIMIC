module fake_jpeg_2447_n_97 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_30),
.B1(n_32),
.B2(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_49),
.B1(n_36),
.B2(n_39),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_27),
.B1(n_31),
.B2(n_29),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_27),
.B1(n_29),
.B2(n_34),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_41),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_14),
.C(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_58),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_13),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_15),
.Y(n_58)
);

NOR3xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_44),
.C(n_46),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_64),
.C(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_46),
.B1(n_45),
.B2(n_38),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_66),
.B1(n_3),
.B2(n_5),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_68),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_72),
.B1(n_6),
.B2(n_7),
.Y(n_81)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_75),
.Y(n_82)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_5),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_10),
.Y(n_86)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_9),
.Y(n_85)
);

NOR4xp25_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_18),
.C(n_25),
.D(n_24),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_17),
.B(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_6),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_81),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_8),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_88),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_90),
.A2(n_80),
.B1(n_72),
.B2(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_89),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_86),
.B1(n_87),
.B2(n_22),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_12),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_26),
.Y(n_97)
);


endmodule