module fake_jpeg_29662_n_522 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_522);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_522;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_12),
.B(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_48),
.Y(n_146)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_49),
.Y(n_149)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_59),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_72),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_75),
.Y(n_121)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_0),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_0),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_29),
.Y(n_119)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_41),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_46),
.B(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_102),
.B(n_110),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_44),
.B1(n_19),
.B2(n_30),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_104),
.A2(n_124),
.B1(n_154),
.B2(n_158),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_62),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_54),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_96),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_119),
.B(n_29),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_51),
.A2(n_20),
.B1(n_41),
.B2(n_39),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_43),
.C(n_30),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_19),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_67),
.B(n_45),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_151),
.Y(n_186)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_52),
.B(n_17),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_28),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_64),
.A2(n_17),
.B1(n_39),
.B2(n_38),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_66),
.A2(n_16),
.B1(n_38),
.B2(n_37),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_163),
.Y(n_233)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_164),
.Y(n_241)
);

BUFx16f_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_166),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_196),
.C(n_45),
.Y(n_223)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_113),
.B(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_169),
.B(n_177),
.Y(n_227)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_175),
.B(n_199),
.Y(n_246)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_118),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_96),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_180),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_115),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_197),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_138),
.A2(n_65),
.B1(n_75),
.B2(n_48),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_182),
.A2(n_190),
.B1(n_206),
.B2(n_104),
.Y(n_214)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_63),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_184),
.B(n_207),
.Y(n_240)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_189),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_123),
.A2(n_65),
.B1(n_75),
.B2(n_48),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

BUFx24_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_128),
.B(n_44),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_120),
.B(n_19),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_203),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_205),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_162),
.A2(n_95),
.B1(n_89),
.B2(n_84),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_101),
.B(n_28),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_144),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_214),
.B(n_215),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_181),
.B(n_125),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_192),
.A2(n_157),
.B1(n_155),
.B2(n_126),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g269 ( 
.A1(n_219),
.A2(n_200),
.B1(n_183),
.B2(n_173),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_166),
.Y(n_265)
);

AOI32xp33_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_149),
.A3(n_155),
.B1(n_157),
.B2(n_126),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_147),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_197),
.A2(n_127),
.B1(n_142),
.B2(n_141),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_244),
.B1(n_178),
.B2(n_142),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_206),
.A2(n_111),
.B1(n_133),
.B2(n_81),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_63),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_190),
.B(n_182),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_203),
.Y(n_256)
);

AO22x1_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_196),
.B1(n_167),
.B2(n_186),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_248),
.A2(n_263),
.B(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_37),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_253),
.B(n_36),
.Y(n_296)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_215),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_256),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_258),
.A2(n_261),
.B1(n_269),
.B2(n_241),
.Y(n_302)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_20),
.C(n_34),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_201),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_260),
.B(n_267),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_130),
.B1(n_141),
.B2(n_163),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_147),
.B(n_170),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_237),
.B(n_218),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_218),
.Y(n_298)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_271),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_214),
.A2(n_130),
.B1(n_78),
.B2(n_79),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_215),
.B(n_168),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_185),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_164),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_273),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_221),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_188),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_275),
.B(n_276),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_212),
.B(n_76),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_229),
.A2(n_194),
.B1(n_211),
.B2(n_241),
.Y(n_277)
);

OR2x2_ASAP7_75t_SL g279 ( 
.A(n_221),
.B(n_166),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_237),
.C(n_217),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_250),
.A2(n_244),
.B1(n_228),
.B2(n_211),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_284),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_252),
.A2(n_243),
.B1(n_239),
.B2(n_236),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_249),
.A2(n_243),
.B1(n_239),
.B2(n_236),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_297),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_248),
.B(n_229),
.C(n_224),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_298),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_295),
.A2(n_304),
.B(n_270),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_311),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_172),
.B1(n_174),
.B2(n_205),
.Y(n_297)
);

AO21x2_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_216),
.B(n_233),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g321 ( 
.A1(n_299),
.A2(n_268),
.B(n_269),
.Y(n_321)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_274),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_303),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_231),
.B(n_213),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_273),
.B(n_34),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_279),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_260),
.A2(n_234),
.B1(n_230),
.B2(n_213),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_222),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_278),
.A2(n_231),
.B1(n_234),
.B2(n_230),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_272),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_275),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_321),
.Y(n_348)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_315),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_316),
.B(n_320),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_265),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_337),
.C(n_340),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_SL g354 ( 
.A(n_318),
.B(n_307),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_280),
.A2(n_278),
.B(n_248),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_322),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_253),
.Y(n_323)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_334),
.Y(n_347)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_326),
.Y(n_368)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_327),
.Y(n_345)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_276),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_335),
.Y(n_349)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_242),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_264),
.B(n_258),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_336),
.A2(n_338),
.B(n_341),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_256),
.C(n_271),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_262),
.B(n_254),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_266),
.C(n_267),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_299),
.A2(n_251),
.B1(n_269),
.B2(n_242),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_269),
.C(n_222),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_340),
.C(n_337),
.Y(n_356)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_289),
.B(n_269),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_289),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_301),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_313),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_346),
.B(n_359),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_288),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_356),
.C(n_367),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_SL g405 ( 
.A(n_354),
.B(n_283),
.C(n_297),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_336),
.A2(n_295),
.B(n_299),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_358),
.A2(n_312),
.B(n_332),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_303),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_322),
.B(n_308),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_360),
.B(n_361),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_328),
.Y(n_361)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_319),
.B(n_306),
.C(n_293),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_327),
.Y(n_369)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_369),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_328),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_372),
.Y(n_380)
);

AO21x2_ASAP7_75t_L g371 ( 
.A1(n_321),
.A2(n_299),
.B(n_310),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_371),
.A2(n_321),
.B1(n_299),
.B2(n_332),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_324),
.B(n_281),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g374 ( 
.A(n_325),
.B(n_306),
.CI(n_281),
.CON(n_374),
.SN(n_374)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_312),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_287),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_284),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_329),
.B(n_294),
.Y(n_376)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_376),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_294),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_350),
.C(n_356),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_369),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_387),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_399),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_347),
.A2(n_314),
.B1(n_364),
.B2(n_349),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_388),
.A2(n_393),
.B1(n_395),
.B2(n_401),
.Y(n_429)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_348),
.Y(n_409)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_355),
.A2(n_314),
.B1(n_333),
.B2(n_343),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_347),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_396),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_351),
.A2(n_301),
.B1(n_333),
.B2(n_344),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_376),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_363),
.Y(n_397)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_397),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_367),
.C(n_319),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_404),
.C(n_374),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_368),
.B(n_362),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_371),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_355),
.A2(n_338),
.B1(n_334),
.B2(n_331),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_SL g402 ( 
.A(n_354),
.B(n_318),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_402),
.A2(n_405),
.B1(n_371),
.B2(n_373),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_352),
.B(n_320),
.C(n_285),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_406),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_377),
.C(n_365),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_407),
.B(n_428),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_392),
.A2(n_366),
.B1(n_365),
.B2(n_358),
.Y(n_408)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_421),
.C(n_426),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_404),
.B(n_381),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_411),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_348),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_417),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_398),
.B(n_348),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_401),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_420),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_374),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_371),
.Y(n_421)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_424),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_425),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_371),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_384),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_380),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_451),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_386),
.C(n_383),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_417),
.C(n_415),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_429),
.A2(n_386),
.B1(n_396),
.B2(n_405),
.Y(n_440)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_440),
.Y(n_452)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_419),
.Y(n_441)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_444),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_430),
.A2(n_383),
.B(n_378),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_SL g460 ( 
.A(n_443),
.B(n_287),
.C(n_216),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_416),
.Y(n_444)
);

NOR2x1p5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_378),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_418),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_422),
.A2(n_406),
.B1(n_391),
.B2(n_389),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_446),
.A2(n_450),
.B1(n_421),
.B2(n_309),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_382),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_448),
.B(n_449),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_414),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_422),
.A2(n_353),
.B1(n_373),
.B2(n_403),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_434),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_436),
.A2(n_409),
.B(n_411),
.Y(n_455)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_458),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_457),
.B(n_462),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_431),
.A2(n_420),
.B1(n_282),
.B2(n_251),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_466),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_287),
.C(n_165),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_165),
.C(n_176),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_463),
.B(n_464),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_432),
.A2(n_36),
.B1(n_187),
.B2(n_139),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_216),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_468),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_439),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_171),
.C(n_156),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_116),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_447),
.Y(n_468)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_445),
.B(n_147),
.CI(n_193),
.CON(n_469),
.SN(n_469)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_469),
.B(n_459),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_452),
.A2(n_443),
.B(n_445),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_471),
.A2(n_476),
.B(n_461),
.Y(n_488)
);

OA21x2_ASAP7_75t_SL g472 ( 
.A1(n_468),
.A2(n_433),
.B(n_446),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_472),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_454),
.A2(n_433),
.B(n_450),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_463),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_465),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_456),
.A2(n_2),
.B(n_4),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_44),
.B1(n_131),
.B2(n_6),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_481),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_453),
.A2(n_193),
.B1(n_143),
.B2(n_7),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_482),
.B(n_485),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_457),
.A2(n_143),
.B1(n_5),
.B2(n_7),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_4),
.Y(n_498)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_488),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_473),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_492),
.B(n_495),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_490),
.B(n_493),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_480),
.A2(n_469),
.B(n_462),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_467),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_486),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_497),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_143),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_498),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_4),
.Y(n_499)
);

NAND3xp33_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_4),
.C(n_5),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_483),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_504),
.Y(n_510)
);

NAND3xp33_ASAP7_75t_SL g504 ( 
.A(n_489),
.B(n_476),
.C(n_482),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_505),
.A2(n_508),
.B(n_491),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_492),
.A2(n_479),
.B(n_7),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_509),
.B(n_511),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_506),
.A2(n_502),
.B(n_503),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_501),
.A2(n_494),
.B(n_487),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_512),
.B(n_513),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_504),
.A2(n_5),
.B(n_9),
.Y(n_513)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_510),
.B(n_507),
.CI(n_11),
.CON(n_514),
.SN(n_514)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_10),
.C(n_12),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_517),
.B(n_518),
.C(n_516),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_515),
.A2(n_10),
.B(n_12),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_519),
.B(n_12),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_14),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_521),
.B(n_14),
.Y(n_522)
);


endmodule