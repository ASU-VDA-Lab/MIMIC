module fake_jpeg_18109_n_67 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_55;
wire n_64;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_43;
wire n_37;
wire n_50;
wire n_29;
wire n_32;
wire n_66;

INVx3_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_9),
.B(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_1),
.B1(n_5),
.B2(n_8),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_45),
.B(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_5),
.B1(n_34),
.B2(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_36),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_22),
.A2(n_41),
.B1(n_20),
.B2(n_32),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_49),
.B(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_52),
.B(n_44),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_58),
.B1(n_50),
.B2(n_51),
.Y(n_60)
);

OAI21x1_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_50),
.B(n_53),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_53),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_33),
.C(n_35),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_29),
.C(n_24),
.Y(n_64)
);

AOI322xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.A3(n_29),
.B1(n_42),
.B2(n_23),
.C1(n_54),
.C2(n_27),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_47),
.B(n_42),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_48),
.B1(n_24),
.B2(n_39),
.Y(n_67)
);


endmodule