module real_jpeg_23803_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_31),
.B1(n_38),
.B2(n_40),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_4),
.A2(n_7),
.B1(n_31),
.B2(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_50),
.C(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_4),
.B(n_49),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_4),
.B(n_38),
.C(n_69),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_4),
.B(n_24),
.C(n_35),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_4),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_4),
.B(n_83),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_4),
.B(n_100),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_39),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_39),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_6),
.A2(n_39),
.B1(n_51),
.B2(n_52),
.Y(n_99)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_80),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_8),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_9),
.A2(n_25),
.B1(n_38),
.B2(n_40),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_11),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_120),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_119),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_101),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_16),
.B(n_101),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_75),
.C(n_84),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_17),
.A2(n_18),
.B1(n_75),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_45),
.B2(n_46),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_19),
.B(n_47),
.C(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_21),
.A2(n_32),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_21),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_27),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_22),
.A2(n_29),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_24),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_26),
.B(n_29),
.Y(n_114)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_26),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_28),
.A2(n_94),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_32),
.A2(n_126),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_32),
.B(n_176),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_32),
.A2(n_107),
.B1(n_109),
.B2(n_126),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_32),
.B(n_107),
.C(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B(n_41),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_33),
.A2(n_41),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_33),
.B(n_131),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_37),
.A2(n_42),
.B1(n_43),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_38),
.Y(n_40)
);

OA22x2_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_40),
.B1(n_69),
.B2(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_38),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_42),
.B(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_43),
.Y(n_131)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_64),
.B1(n_65),
.B2(n_74),
.Y(n_46)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_47),
.A2(n_74),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_55),
.B(n_58),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_59),
.B1(n_62),
.B2(n_86),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_54),
.B1(n_56),
.B2(n_61),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_52),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_52),
.B(n_162),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B(n_72),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_73),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_73),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_99),
.B(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_109),
.C(n_129),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_75),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_81),
.Y(n_105)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_81),
.A2(n_82),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_81),
.A2(n_82),
.B1(n_159),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_153),
.C(n_159),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_82),
.B(n_92),
.C(n_192),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_84),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.C(n_97),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_85),
.A2(n_97),
.B1(n_110),
.B2(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_91),
.A2(n_92),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_92),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_92),
.B(n_184),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_96),
.B(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_146),
.C(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_97),
.A2(n_136),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_109),
.B1(n_129),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_112),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_149),
.B(n_210),
.C(n_215),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_138),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_122),
.B(n_138),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_134),
.B2(n_137),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_133),
.C(n_137),
.Y(n_211)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.C(n_145),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_140),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_148),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_146),
.B(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_209),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_168),
.B(n_208),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_165),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_152),
.B(n_165),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_154),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_173),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_201),
.B(n_207),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_195),
.B(n_200),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_187),
.B(n_194),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_186),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_174),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_185),
.Y(n_177)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_188),
.B(n_189),
.Y(n_194)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_196),
.B(n_197),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_202),
.B(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_212),
.Y(n_215)
);


endmodule