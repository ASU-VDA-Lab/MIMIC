module fake_jpeg_3505_n_466 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_466);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_466;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_48),
.Y(n_56)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_7),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_60),
.B(n_83),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_14),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_100),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_25),
.B(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_84),
.B(n_36),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_37),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_97),
.A2(n_30),
.B1(n_39),
.B2(n_32),
.Y(n_143)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_30),
.B(n_31),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_27),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_60),
.A2(n_34),
.B(n_27),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_116),
.C(n_125),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_23),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_68),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_88),
.A2(n_34),
.B1(n_20),
.B2(n_32),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_138),
.A2(n_81),
.B1(n_41),
.B2(n_47),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_36),
.B1(n_45),
.B2(n_28),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_69),
.A2(n_34),
.B1(n_21),
.B2(n_43),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_93),
.B1(n_78),
.B2(n_70),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_98),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_156),
.Y(n_161)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_160),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_103),
.A2(n_72),
.B1(n_69),
.B2(n_61),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_189),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_57),
.B(n_72),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_163),
.A2(n_119),
.B(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_164),
.Y(n_233)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_103),
.A2(n_99),
.B1(n_96),
.B2(n_95),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_167),
.A2(n_175),
.B1(n_202),
.B2(n_53),
.Y(n_228)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_31),
.B1(n_39),
.B2(n_86),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_171),
.B1(n_179),
.B2(n_181),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_105),
.B(n_64),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_63),
.B1(n_90),
.B2(n_85),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_177),
.A2(n_192),
.B1(n_200),
.B2(n_119),
.Y(n_219)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_52),
.B1(n_67),
.B2(n_66),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_62),
.B1(n_58),
.B2(n_40),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_28),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_184),
.B(n_191),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_45),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_195),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_110),
.B(n_17),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_17),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_201),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_135),
.A2(n_43),
.B1(n_21),
.B2(n_41),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_120),
.A2(n_41),
.B1(n_17),
.B2(n_43),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_203),
.A2(n_130),
.B1(n_147),
.B2(n_128),
.Y(n_211)
);

AOI32xp33_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_136),
.A3(n_133),
.B1(n_131),
.B2(n_122),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_137),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_211),
.A2(n_174),
.B1(n_178),
.B2(n_160),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_112),
.B1(n_154),
.B2(n_115),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_214),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_161),
.B(n_155),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_226),
.C(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_219),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_171),
.A2(n_128),
.B1(n_147),
.B2(n_126),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_228),
.B1(n_162),
.B2(n_167),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_187),
.C(n_195),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_163),
.A2(n_134),
.B(n_124),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_162),
.B(n_123),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_123),
.C(n_124),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_244),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_241),
.A2(n_251),
.B1(n_258),
.B2(n_259),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_233),
.B1(n_216),
.B2(n_213),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_243),
.A2(n_218),
.B(n_234),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_212),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_205),
.B(n_161),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_187),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_231),
.A2(n_192),
.B(n_188),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_249),
.A2(n_0),
.B(n_1),
.Y(n_296)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_228),
.A2(n_175),
.B1(n_157),
.B2(n_126),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_252),
.B(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_169),
.B1(n_157),
.B2(n_113),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_254),
.A2(n_261),
.B1(n_263),
.B2(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_204),
.A2(n_198),
.B1(n_194),
.B2(n_186),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_210),
.A2(n_189),
.B1(n_191),
.B2(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_168),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_265),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_121),
.B1(n_141),
.B2(n_185),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_215),
.B(n_159),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_121),
.B1(n_141),
.B2(n_172),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_206),
.A2(n_221),
.B1(n_227),
.B2(n_224),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_232),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_201),
.B1(n_199),
.B2(n_43),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_21),
.C(n_47),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_216),
.C(n_225),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_269),
.B(n_259),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_271),
.A2(n_272),
.B(n_249),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_240),
.A2(n_225),
.B1(n_229),
.B2(n_233),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_260),
.Y(n_274)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_268),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_209),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_278),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_241),
.A2(n_209),
.B1(n_213),
.B2(n_232),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_282),
.A2(n_289),
.B1(n_264),
.B2(n_254),
.Y(n_302)
);

OAI32xp33_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_217),
.A3(n_238),
.B1(n_223),
.B2(n_229),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_285),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g285 ( 
.A1(n_242),
.A2(n_217),
.B1(n_238),
.B2(n_223),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_235),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_291),
.C(n_293),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_243),
.B1(n_257),
.B2(n_258),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_296),
.B(n_243),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_222),
.C(n_220),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_222),
.C(n_220),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_245),
.B(n_235),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_268),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_289),
.B1(n_281),
.B2(n_274),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_300),
.B1(n_254),
.B2(n_277),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_290),
.B1(n_282),
.B2(n_284),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_269),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_304),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_265),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_303),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_240),
.B(n_249),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_305),
.A2(n_322),
.B(n_240),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_252),
.A3(n_248),
.B1(n_253),
.B2(n_262),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_308),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_244),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_286),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_295),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_310),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_284),
.B(n_239),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_311),
.B(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_291),
.B(n_255),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_294),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_318),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_320),
.C(n_276),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_295),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_296),
.Y(n_319)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_319),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_267),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_311),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_351),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_329),
.C(n_335),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_290),
.C(n_271),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_336),
.A2(n_349),
.B1(n_350),
.B2(n_331),
.Y(n_366)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_314),
.Y(n_337)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_342),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_292),
.C(n_270),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_345),
.C(n_316),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_270),
.C(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_347),
.A2(n_322),
.B(n_305),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_285),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_348),
.B(n_306),
.Y(n_360)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_327),
.B(n_320),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_353),
.B(n_360),
.Y(n_395)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_261),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_344),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_362),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_302),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_358),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_328),
.A2(n_304),
.B(n_308),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_330),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_326),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_368),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_309),
.B1(n_319),
.B2(n_323),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_366),
.B1(n_367),
.B2(n_369),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_309),
.B1(n_318),
.B2(n_310),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_328),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_337),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_347),
.A2(n_323),
.B(n_275),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_342),
.A2(n_277),
.B1(n_323),
.B2(n_273),
.Y(n_372)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_329),
.B(n_283),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_338),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_368),
.A2(n_331),
.B1(n_334),
.B2(n_338),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_377),
.A2(n_381),
.B1(n_387),
.B2(n_394),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_325),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_379),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_371),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_345),
.C(n_335),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_388),
.C(n_353),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_363),
.A2(n_338),
.B1(n_340),
.B2(n_348),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_382),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_385),
.Y(n_402)
);

XOR2x2_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_365),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_333),
.B1(n_285),
.B2(n_263),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_333),
.C(n_250),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_355),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_359),
.A2(n_248),
.B1(n_266),
.B2(n_8),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_388),
.A2(n_358),
.B(n_360),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_381),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_400),
.B(n_401),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_376),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_403),
.Y(n_424)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_391),
.Y(n_404)
);

BUFx24_ASAP7_75t_SL g427 ( 
.A(n_404),
.Y(n_427)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_405),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_413),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_396),
.A2(n_375),
.B1(n_369),
.B2(n_356),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_408),
.A2(n_412),
.B1(n_384),
.B2(n_389),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_373),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_390),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_373),
.C(n_375),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_410),
.B(n_411),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_370),
.C(n_361),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_393),
.A2(n_370),
.B1(n_361),
.B2(n_374),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_374),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_400),
.B(n_395),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_409),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_418),
.A2(n_426),
.B(n_410),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_420),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_384),
.C(n_389),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_377),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_421),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_422),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_411),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_406),
.A2(n_387),
.B1(n_382),
.B2(n_8),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_425),
.A2(n_3),
.B1(n_4),
.B2(n_10),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_399),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_426)
);

NOR2x1_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_433),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_431),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_416),
.B(n_403),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_407),
.C(n_1),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_435),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_4),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_0),
.C(n_1),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_438),
.Y(n_448)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_439),
.B(n_440),
.Y(n_449)
);

INVx6_ASAP7_75t_L g440 ( 
.A(n_427),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_441),
.B(n_424),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_444),
.B(n_445),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_421),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_424),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_447),
.A2(n_450),
.B(n_426),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_430),
.A2(n_434),
.B(n_435),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_446),
.Y(n_451)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_451),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_436),
.Y(n_452)
);

NOR3xp33_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_456),
.C(n_13),
.Y(n_459)
);

AO21x2_ASAP7_75t_L g458 ( 
.A1(n_454),
.A2(n_443),
.B(n_12),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_433),
.C(n_440),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_455),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_3),
.Y(n_456)
);

OAI21xp33_ASAP7_75t_SL g462 ( 
.A1(n_458),
.A2(n_459),
.B(n_2),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_460),
.B(n_452),
.C(n_453),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_461),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_463),
.B(n_457),
.C(n_462),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_464),
.A2(n_2),
.B(n_460),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_465),
.B(n_2),
.Y(n_466)
);


endmodule