module real_jpeg_7334_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_0),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_0),
.Y(n_238)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g362 ( 
.A(n_1),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_1),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_1),
.Y(n_432)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_1),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_2),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_2),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_2),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_2),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_2),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_2),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_3),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_3),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_3),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_3),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_3),
.B(n_172),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_4),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_4),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_4),
.Y(n_345)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_5),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_6),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_7),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_7),
.Y(n_194)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_7),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_8),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_8),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_8),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_8),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_8),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_8),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_8),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_9),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_9),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_9),
.B(n_142),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_9),
.B(n_347),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_9),
.B(n_149),
.Y(n_408)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_13),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_13),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_13),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_13),
.B(n_313),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_13),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_13),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_13),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_13),
.B(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_14),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_14),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_14),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_14),
.B(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_14),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_14),
.B(n_45),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_15),
.B(n_216),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_15),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_15),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_15),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_15),
.B(n_159),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_15),
.B(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_16),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_16),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_16),
.B(n_99),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_16),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_17),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_17),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_17),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_17),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_17),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_17),
.B(n_333),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_17),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_17),
.B(n_430),
.Y(n_429)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_45),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_19),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_19),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_19),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_19),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_19),
.B(n_387),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_19),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_19),
.B(n_485),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_539),
.B(n_541),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_46),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_26),
.A2(n_27),
.B1(n_36),
.B2(n_62),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_36),
.C(n_42),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_28),
.B(n_379),
.Y(n_378)
);

INVx6_ASAP7_75t_L g485 ( 
.A(n_29),
.Y(n_485)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_30),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_50),
.C(n_57),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_40),
.Y(n_315)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_41),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_41),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_72),
.C(n_74),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_47),
.B(n_529),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_63),
.C(n_65),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_48),
.A2(n_49),
.B1(n_525),
.B2(n_526),
.Y(n_524)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_66),
.C(n_68),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_56),
.A2(n_57),
.B1(n_68),
.B2(n_486),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_60),
.Y(n_389)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_61),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_63),
.B(n_65),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_66),
.A2(n_67),
.B1(n_488),
.B2(n_489),
.Y(n_487)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_68),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_68),
.A2(n_441),
.B1(n_442),
.B2(n_486),
.Y(n_503)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_530),
.Y(n_529)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_74),
.Y(n_530)
);

AO21x1_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_459),
.B(n_532),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_415),
.B(n_458),
.Y(n_78)
);

AOI21x1_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_366),
.B(n_414),
.Y(n_79)
);

OAI21x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_319),
.B(n_365),
.Y(n_80)
);

AOI21x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_281),
.B(n_318),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_204),
.B(n_280),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_187),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_84),
.B(n_187),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_130),
.B2(n_186),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_85),
.B(n_131),
.C(n_169),
.Y(n_317)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_107),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_87),
.B(n_108),
.C(n_129),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_101),
.C(n_105),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_88),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_192)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_101),
.B(n_105),
.Y(n_203)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_116),
.B1(n_128),
.B2(n_129),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B(n_115),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_111),
.Y(n_115)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_115),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_115),
.B(n_286),
.C(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g547 ( 
.A(n_116),
.Y(n_547)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.CI(n_124),
.CON(n_116),
.SN(n_116)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_117),
.B(n_120),
.C(n_124),
.Y(n_316)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_169),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_145),
.C(n_161),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_137),
.C(n_141),
.Y(n_185)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_140),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_140),
.Y(n_444)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_145),
.A2(n_146),
.B1(n_161),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_157),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_147),
.A2(n_148),
.B1(n_157),
.B2(n_158),
.Y(n_273)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_149),
.Y(n_439)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_150),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_151),
.B(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_155),
.Y(n_250)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_156),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_156),
.Y(n_343)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_156),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_156),
.Y(n_455)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_163),
.B(n_449),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_163),
.B(n_468),
.Y(n_467)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_183),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_170),
.B(n_184),
.C(n_185),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_171),
.B(n_179),
.C(n_181),
.Y(n_296)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_174),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_179),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.C(n_202),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_188),
.B(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_191),
.B(n_202),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.C(n_195),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_192),
.B(n_193),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_195),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_198),
.Y(n_244)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_200),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21x1_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_275),
.B(n_279),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_260),
.B(n_274),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_241),
.B(n_259),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_229),
.B(n_240),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_217),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_217),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_213),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_212),
.Y(n_356)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_212),
.Y(n_381)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_224),
.B2(n_225),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_221),
.C(n_224),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_227),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_235),
.B(n_239),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_232),
.Y(n_239)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_233),
.Y(n_397)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_258),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_258),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_245),
.C(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_253),
.C(n_257),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_257),
.Y(n_251)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_263),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_270),
.C(n_271),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_317),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_282),
.B(n_317),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_298),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_285),
.C(n_298),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_295),
.B2(n_297),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_291),
.C(n_292),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_301),
.C(n_310),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_310),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_302),
.B(n_304),
.C(n_306),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g449 ( 
.A(n_309),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_316),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_314),
.C(n_316),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_321),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_322),
.B(n_338),
.C(n_363),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_338),
.B1(n_363),
.B2(n_364),
.Y(n_323)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_324),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_337),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_328),
.C(n_329),
.Y(n_368)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_336),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_331),
.B(n_332),
.C(n_336),
.Y(n_403)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_349),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_350),
.C(n_351),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_339),
.Y(n_545)
);

FAx1_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_344),
.CI(n_346),
.CON(n_339),
.SN(n_339)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_340),
.B(n_344),
.C(n_346),
.Y(n_411)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_360),
.B2(n_361),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_353)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_354),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_359),
.C(n_360),
.Y(n_383)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_357),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_357),
.A2(n_359),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_359),
.B(n_373),
.C(n_378),
.Y(n_427)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_413),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_413),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_368),
.B(n_370),
.C(n_399),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_399),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_382),
.B2(n_398),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_383),
.C(n_384),
.Y(n_421)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_376),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_375),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_377),
.A2(n_378),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_377),
.B(n_436),
.C(n_441),
.Y(n_504)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_382),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_395),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_390),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_386),
.B(n_390),
.C(n_395),
.Y(n_446)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_402),
.B2(n_412),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_403),
.C(n_404),
.Y(n_417)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_402),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_411),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_408),
.B1(n_409),
.B2(n_410),
.Y(n_405)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_406),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_408),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_409),
.C(n_425),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_408),
.A2(n_410),
.B1(n_429),
.B2(n_433),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_410),
.B(n_427),
.C(n_433),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_411),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_457),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_457),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_417),
.B(n_419),
.C(n_434),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_434),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_420),
.B(n_424),
.C(n_426),
.Y(n_512)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_429),
.Y(n_433)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_445),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_446),
.C(n_447),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_440),
.Y(n_435)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_484),
.C(n_486),
.Y(n_483)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_450),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_448),
.B(n_453),
.C(n_456),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_453),
.B1(n_454),
.B2(n_456),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_451),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_454),
.Y(n_453)
);

NOR3xp33_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_517),
.C(n_527),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_513),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_462),
.A2(n_536),
.B(n_537),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_506),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_463),
.B(n_506),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_480),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_464),
.B(n_481),
.C(n_501),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.C(n_478),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_465),
.B(n_508),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_466),
.A2(n_478),
.B1(n_479),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_466),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_471),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_467),
.B(n_472),
.C(n_473),
.Y(n_493)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_477),
.Y(n_499)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_501),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_492),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_487),
.B1(n_490),
.B2(n_491),
.Y(n_482)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_483),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_491),
.C(n_492),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_487),
.Y(n_491)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_493),
.B(n_497),
.C(n_500),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_497),
.B1(n_498),
.B2(n_500),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_495),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_498),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_504),
.C(n_505),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_511),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_505),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_510),
.C(n_512),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_510),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_512),
.B(n_515),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_516),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_516),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_535),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_520),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_522),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_523),
.C(n_524),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_524),
.Y(n_522)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_533),
.B(n_534),
.C(n_538),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_531),
.Y(n_538)
);

INVx8_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_540),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_544),
.Y(n_541)
);

BUFx12f_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);


endmodule