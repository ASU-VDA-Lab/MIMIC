module fake_jpeg_29853_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_8),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_75),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_66),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_87),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_76),
.Y(n_86)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_65),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_90),
.A2(n_70),
.B1(n_46),
.B2(n_61),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_106),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_47),
.B(n_56),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_109),
.B(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_1),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_104),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_98),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_63),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_6),
.C(n_7),
.Y(n_129)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_50),
.B1(n_58),
.B2(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_59),
.C(n_57),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_55),
.C(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_23),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_125),
.B(n_20),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_116),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_118),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_123),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_5),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_25),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_130),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_24),
.B(n_39),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_5),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_6),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_7),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_27),
.C(n_10),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_26),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_141),
.B1(n_118),
.B2(n_129),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_143),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_21),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_146),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_140),
.B1(n_133),
.B2(n_138),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_120),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_154),
.C(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_153),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_157),
.A3(n_158),
.B1(n_152),
.B2(n_148),
.C1(n_155),
.C2(n_151),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_144),
.B1(n_147),
.B2(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

OAI321xp33_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_148),
.A3(n_158),
.B1(n_135),
.B2(n_34),
.C(n_35),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_29),
.B(n_31),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_32),
.B(n_37),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_164),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_166),
.Y(n_167)
);


endmodule