module fake_jpeg_11743_n_488 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_488);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_488;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_50),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_51),
.B(n_53),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_17),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_56),
.B(n_79),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_58),
.B(n_74),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_61),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_27),
.B(n_0),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_33),
.C(n_49),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_0),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_47),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_37),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_89),
.Y(n_151)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_32),
.Y(n_92)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_69),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_19),
.B1(n_40),
.B2(n_30),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_111),
.A2(n_19),
.B1(n_94),
.B2(n_91),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_49),
.Y(n_163)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_158),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_159),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_53),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_160),
.B(n_165),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_163),
.A2(n_171),
.B(n_192),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_93),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_171),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_55),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_33),
.B1(n_49),
.B2(n_22),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_166),
.A2(n_173),
.B1(n_181),
.B2(n_188),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_114),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_179),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_78),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_129),
.A2(n_22),
.B1(n_30),
.B2(n_88),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_128),
.B(n_130),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_77),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_190),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_142),
.A2(n_22),
.B1(n_30),
.B2(n_88),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_154),
.C(n_153),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_182),
.B(n_97),
.Y(n_231)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

BUFx16f_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_185),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_116),
.B(n_46),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_196),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_101),
.A2(n_87),
.B1(n_69),
.B2(n_40),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_111),
.A2(n_96),
.B1(n_81),
.B2(n_95),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_28),
.B1(n_99),
.B2(n_21),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_104),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_194),
.B1(n_52),
.B2(n_72),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_41),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_201),
.Y(n_234)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_193),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_106),
.A2(n_86),
.B1(n_85),
.B2(n_64),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

AO22x1_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_112),
.B1(n_75),
.B2(n_34),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_127),
.A2(n_87),
.B1(n_28),
.B2(n_41),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_199),
.A2(n_124),
.B1(n_21),
.B2(n_47),
.Y(n_250)
);

CKINVDCx9p33_ASAP7_75t_R g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_200),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_110),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_100),
.B(n_36),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_206),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_113),
.B(n_50),
.Y(n_208)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_120),
.B1(n_132),
.B2(n_121),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_209),
.A2(n_210),
.B1(n_237),
.B2(n_252),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_144),
.B1(n_132),
.B2(n_121),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_213),
.A2(n_232),
.B1(n_175),
.B2(n_168),
.Y(n_279)
);

AO21x2_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_117),
.B(n_98),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_221),
.B1(n_222),
.B2(n_170),
.Y(n_265)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_164),
.A2(n_80),
.A3(n_105),
.B1(n_134),
.B2(n_107),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_231),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_SL g278 ( 
.A1(n_219),
.A2(n_250),
.B(n_36),
.Y(n_278)
);

AO22x2_ASAP7_75t_L g221 ( 
.A1(n_163),
.A2(n_57),
.B1(n_63),
.B2(n_67),
.Y(n_221)
);

AO21x2_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_144),
.B(n_100),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_200),
.C(n_205),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_19),
.B1(n_43),
.B2(n_48),
.Y(n_232)
);

OA22x2_ASAP7_75t_SL g238 ( 
.A1(n_163),
.A2(n_71),
.B1(n_68),
.B2(n_139),
.Y(n_238)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_182),
.B(n_46),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_27),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_195),
.A2(n_45),
.B(n_34),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_43),
.C(n_35),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_193),
.A2(n_45),
.B1(n_35),
.B2(n_48),
.Y(n_252)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_223),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_254),
.B(n_256),
.Y(n_318)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_262),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_234),
.A2(n_183),
.B1(n_167),
.B2(n_197),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_258),
.A2(n_260),
.B(n_277),
.Y(n_308)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_215),
.A2(n_161),
.B(n_157),
.Y(n_260)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_261),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_162),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_263),
.B(n_214),
.C(n_251),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_279),
.Y(n_295)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_186),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_272),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_230),
.A2(n_202),
.B1(n_156),
.B2(n_177),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_285),
.B1(n_220),
.B2(n_231),
.Y(n_296)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_218),
.Y(n_271)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_184),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_197),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_275),
.Y(n_324)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_281),
.B1(n_283),
.B2(n_289),
.Y(n_293)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_233),
.B(n_167),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_235),
.B(n_176),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_225),
.B(n_211),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_222),
.A2(n_174),
.B1(n_178),
.B2(n_47),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_287),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_204),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_159),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_211),
.A2(n_204),
.B(n_184),
.C(n_170),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_290),
.A2(n_247),
.B(n_219),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_227),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_234),
.B1(n_222),
.B2(n_238),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_299),
.A2(n_300),
.B1(n_307),
.B2(n_312),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_267),
.A2(n_222),
.B1(n_238),
.B2(n_246),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_264),
.A2(n_228),
.B1(n_237),
.B2(n_215),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_303),
.A2(n_309),
.B1(n_311),
.B2(n_313),
.Y(n_333)
);

AO22x1_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_215),
.B1(n_217),
.B2(n_221),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_265),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_215),
.B1(n_221),
.B2(n_240),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_268),
.A2(n_242),
.B1(n_244),
.B2(n_221),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_310),
.A2(n_319),
.B(n_2),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_279),
.A2(n_241),
.B1(n_240),
.B2(n_249),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_260),
.A2(n_241),
.B1(n_248),
.B2(n_239),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_248),
.B1(n_236),
.B2(n_214),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_314),
.B(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_172),
.B(n_158),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_260),
.A2(n_126),
.B1(n_159),
.B2(n_59),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_321),
.A2(n_258),
.B1(n_265),
.B2(n_290),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_263),
.B(n_124),
.C(n_75),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_2),
.Y(n_353)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_318),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_330),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_331),
.A2(n_334),
.B1(n_346),
.B2(n_316),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_338),
.C(n_350),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_299),
.A2(n_265),
.B1(n_272),
.B2(n_262),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_335),
.B(n_337),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_322),
.Y(n_336)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_277),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_269),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_295),
.A2(n_291),
.B1(n_284),
.B2(n_266),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

A2O1A1O1Ixp25_ASAP7_75t_L g341 ( 
.A1(n_302),
.A2(n_271),
.B(n_270),
.C(n_274),
.D(n_276),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_341),
.B(n_349),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_322),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_295),
.Y(n_362)
);

BUFx12_ASAP7_75t_L g343 ( 
.A(n_327),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_343),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_302),
.A2(n_286),
.B(n_280),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_300),
.A2(n_289),
.B1(n_253),
.B2(n_255),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_347),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_303),
.A2(n_273),
.B1(n_261),
.B2(n_259),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_348),
.A2(n_351),
.B(n_355),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_273),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_273),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_295),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_292),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_292),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_354),
.B(n_357),
.Y(n_366)
);

INVx13_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_356),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_3),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_321),
.A2(n_4),
.B(n_5),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_310),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_328),
.A2(n_293),
.B1(n_296),
.B2(n_307),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_360),
.A2(n_382),
.B1(n_386),
.B2(n_331),
.Y(n_403)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_367),
.A2(n_370),
.B1(n_372),
.B2(n_335),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_298),
.C(n_308),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_379),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_357),
.B(n_319),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_369),
.B(n_371),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_338),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_311),
.B1(n_316),
.B2(n_306),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_325),
.Y(n_375)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_375),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_336),
.B(n_323),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_376),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_333),
.A2(n_312),
.B1(n_306),
.B2(n_323),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_333),
.A2(n_301),
.B1(n_297),
.B2(n_294),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_350),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_404),
.C(n_408),
.Y(n_420)
);

XOR2x1_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_329),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_395),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_341),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_391),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_393),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_334),
.C(n_328),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_396),
.C(n_401),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_347),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_345),
.C(n_353),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_397),
.A2(n_373),
.B1(n_385),
.B2(n_361),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_304),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_398),
.B(n_380),
.Y(n_425)
);

OAI21xp33_ASAP7_75t_SL g400 ( 
.A1(n_363),
.A2(n_355),
.B(n_345),
.Y(n_400)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_339),
.Y(n_401)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_348),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_382),
.A2(n_346),
.B1(n_352),
.B2(n_351),
.Y(n_405)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_373),
.B1(n_372),
.B2(n_359),
.Y(n_407)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_407),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_361),
.B(n_301),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_363),
.C(n_360),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_414),
.B(n_415),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_402),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_391),
.A2(n_362),
.B(n_359),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_404),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_366),
.Y(n_423)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_425),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_399),
.B(n_366),
.Y(n_426)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_410),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_427),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_428),
.A2(n_375),
.B1(n_377),
.B2(n_365),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_389),
.C(n_401),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_433),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_418),
.A2(n_373),
.B1(n_406),
.B2(n_387),
.Y(n_433)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_434),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_418),
.A2(n_424),
.B1(n_428),
.B2(n_413),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_437),
.Y(n_449)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_416),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_412),
.A2(n_400),
.B1(n_365),
.B2(n_376),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_419),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_388),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_441),
.C(n_420),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_396),
.C(n_408),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_422),
.A2(n_390),
.B1(n_393),
.B2(n_369),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_443),
.A2(n_421),
.B(n_417),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_444),
.A2(n_419),
.B1(n_429),
.B2(n_304),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_445),
.A2(n_440),
.B(n_358),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_451),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_444),
.A2(n_417),
.B1(n_427),
.B2(n_420),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_441),
.Y(n_463)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_450),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_416),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_436),
.A2(n_377),
.B(n_429),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_454),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_453),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_294),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_430),
.A2(n_431),
.B1(n_434),
.B2(n_437),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_455),
.A2(n_438),
.B1(n_430),
.B2(n_443),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_320),
.C(n_317),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_320),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_455),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_466),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_459),
.A2(n_468),
.B1(n_467),
.B2(n_465),
.Y(n_475)
);

BUFx24_ASAP7_75t_SL g462 ( 
.A(n_457),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_456),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_448),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_464),
.A2(n_445),
.B(n_447),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_449),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_SL g469 ( 
.A(n_463),
.B(n_446),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_470),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_471),
.B(n_472),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_453),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_475),
.Y(n_479)
);

AOI322xp5_ASAP7_75t_L g477 ( 
.A1(n_472),
.A2(n_460),
.A3(n_356),
.B1(n_464),
.B2(n_343),
.C1(n_9),
.C2(n_10),
.Y(n_477)
);

AOI21x1_ASAP7_75t_SL g480 ( 
.A1(n_477),
.A2(n_474),
.B(n_356),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_480),
.B(n_481),
.C(n_479),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_343),
.Y(n_481)
);

AOI21xp33_ASAP7_75t_L g484 ( 
.A1(n_482),
.A2(n_483),
.B(n_4),
.Y(n_484)
);

AOI322xp5_ASAP7_75t_L g483 ( 
.A1(n_480),
.A2(n_476),
.A3(n_343),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_483)
);

AOI322xp5_ASAP7_75t_L g485 ( 
.A1(n_484),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_10),
.C1(n_11),
.C2(n_13),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_485),
.A2(n_6),
.B1(n_14),
.B2(n_15),
.Y(n_486)
);

AO21x1_ASAP7_75t_L g487 ( 
.A1(n_486),
.A2(n_15),
.B(n_6),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_14),
.B(n_236),
.Y(n_488)
);


endmodule