module fake_jpeg_2785_n_129 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_5),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_11),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_45),
.C(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_23),
.B(n_27),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_48),
.Y(n_51)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_1),
.B1(n_7),
.B2(n_6),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_6),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_30),
.A2(n_13),
.B1(n_24),
.B2(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_13),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_43),
.B1(n_24),
.B2(n_31),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_69),
.B1(n_72),
.B2(n_52),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_27),
.B1(n_15),
.B2(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_15),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_38),
.B1(n_45),
.B2(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_69)
);

NOR2x1_ASAP7_75t_R g74 ( 
.A(n_71),
.B(n_51),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_33),
.A2(n_46),
.B1(n_16),
.B2(n_40),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_84),
.B1(n_68),
.B2(n_57),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_70),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_76),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_88),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_89),
.B(n_87),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_67),
.B1(n_55),
.B2(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_92),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_76),
.C(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_104),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_111)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_97),
.B1(n_95),
.B2(n_99),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_100),
.B1(n_94),
.B2(n_98),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_77),
.B1(n_97),
.B2(n_99),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_96),
.B(n_100),
.C(n_74),
.D(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_102),
.B(n_77),
.Y(n_117)
);

BUFx12f_ASAP7_75t_SL g122 ( 
.A(n_117),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_115),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_114),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_117),
.B(n_119),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_113),
.C(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

OAI33xp33_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_125),
.A3(n_122),
.B1(n_113),
.B2(n_86),
.B3(n_82),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_122),
.Y(n_129)
);


endmodule