module fake_jpeg_26927_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_42),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_40),
.Y(n_47)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_24),
.B1(n_34),
.B2(n_21),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_41),
.B1(n_20),
.B2(n_17),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_18),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_40),
.C(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_62),
.B(n_65),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_64),
.B(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_42),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_93),
.B1(n_33),
.B2(n_26),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_70),
.Y(n_114)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_43),
.B(n_39),
.C(n_27),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_97),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_24),
.B1(n_35),
.B2(n_36),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_96),
.B1(n_40),
.B2(n_16),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_78),
.Y(n_122)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_21),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_80),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_40),
.C(n_18),
.Y(n_120)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_94),
.Y(n_118)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_36),
.B1(n_41),
.B2(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_49),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_33),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_38),
.B1(n_16),
.B2(n_23),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_R g97 ( 
.A(n_49),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_20),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_20),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_116),
.B1(n_64),
.B2(n_89),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_33),
.B(n_1),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_107),
.A2(n_32),
.B(n_26),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_38),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_40),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_89),
.B(n_26),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_30),
.B1(n_25),
.B2(n_22),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_17),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_32),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_127),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_88),
.C(n_73),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_32),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_76),
.B(n_87),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_137),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_67),
.B1(n_76),
.B2(n_70),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_131),
.A2(n_127),
.B1(n_103),
.B2(n_109),
.Y(n_168)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_134),
.A2(n_23),
.B1(n_16),
.B2(n_73),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_111),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_96),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_141),
.C(n_151),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_143),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_106),
.B(n_96),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_140),
.A2(n_149),
.B(n_23),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_91),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_148),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_69),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_155),
.B(n_23),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_75),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_69),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_84),
.B1(n_78),
.B2(n_82),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_159),
.B1(n_103),
.B2(n_102),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_107),
.A2(n_30),
.B(n_16),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_158),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_0),
.C(n_2),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_72),
.B1(n_94),
.B2(n_88),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_129),
.B(n_126),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_150),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_115),
.B1(n_129),
.B2(n_102),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_163),
.A2(n_166),
.B1(n_176),
.B2(n_179),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_115),
.B1(n_123),
.B2(n_119),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_164),
.A2(n_168),
.B1(n_173),
.B2(n_180),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_109),
.B(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_171),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_172),
.B(n_177),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_72),
.B1(n_104),
.B2(n_100),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_117),
.B1(n_105),
.B2(n_108),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_174),
.A2(n_185),
.B1(n_189),
.B2(n_136),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_134),
.A2(n_104),
.B1(n_101),
.B2(n_25),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_73),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_178),
.B(n_188),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_25),
.B1(n_22),
.B2(n_29),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_25),
.B1(n_22),
.B2(n_29),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_183),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_135),
.A2(n_22),
.B1(n_29),
.B2(n_23),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_29),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_145),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_155),
.C(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_197),
.B(n_198),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_177),
.B(n_176),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_147),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_141),
.C(n_137),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_190),
.C(n_171),
.Y(n_232)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_157),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_214),
.Y(n_226)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_192),
.B1(n_187),
.B2(n_186),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_151),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_196),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_213),
.B1(n_219),
.B2(n_166),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_191),
.A2(n_152),
.B1(n_148),
.B2(n_136),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_167),
.B(n_132),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_158),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_217),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_168),
.A2(n_171),
.B1(n_162),
.B2(n_163),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_132),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_10),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_174),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_223),
.B(n_212),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_182),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_232),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_233),
.B1(n_244),
.B2(n_218),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_184),
.C(n_164),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_231),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_177),
.B(n_187),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_234),
.A2(n_194),
.B(n_193),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_185),
.C(n_180),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_179),
.C(n_10),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_15),
.C(n_9),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_15),
.C(n_9),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_198),
.C(n_221),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_218),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_224),
.B(n_222),
.C(n_229),
.Y(n_273)
);

XNOR2x2_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_215),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_SL g272 ( 
.A(n_247),
.B(n_257),
.C(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_250),
.C(n_246),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_204),
.Y(n_251)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_252),
.B(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_219),
.B1(n_216),
.B2(n_213),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_194),
.B1(n_209),
.B2(n_205),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_262),
.B(n_263),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_228),
.Y(n_261)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_234),
.A2(n_193),
.B1(n_207),
.B2(n_4),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_226),
.C(n_227),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_226),
.C(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_268),
.C(n_274),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_239),
.C(n_223),
.Y(n_268)
);

BUFx12f_ASAP7_75t_SL g270 ( 
.A(n_247),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_258),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_256),
.B1(n_245),
.B2(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_229),
.C(n_243),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_246),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_11),
.C(n_13),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_279),
.C(n_250),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_5),
.C(n_7),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_11),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_268),
.C(n_267),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_255),
.B1(n_254),
.B2(n_5),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_292),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_7),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_2),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_297),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_291),
.A2(n_270),
.B(n_269),
.Y(n_297)
);

AOI211xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_277),
.B(n_279),
.C(n_266),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_290),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_285),
.B(n_276),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_308),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_288),
.C(n_281),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_287),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_281),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_308),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_316),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_313),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_314),
.C(n_304),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_312),
.B(n_303),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_306),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.C1(n_3),
.C2(n_2),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_12),
.Y(n_321)
);


endmodule