module real_aes_17146_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_0), .A2(n_190), .B1(n_506), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_0), .A2(n_56), .B1(n_399), .B2(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g621 ( .A(n_1), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_1), .A2(n_91), .B1(n_506), .B2(n_642), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_2), .A2(n_790), .B(n_791), .C(n_797), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_2), .B(n_467), .Y(n_809) );
INVx1_ASAP7_75t_L g1272 ( .A(n_3), .Y(n_1272) );
AOI221xp5_ASAP7_75t_L g1294 ( .A1(n_3), .A2(n_141), .B1(n_1020), .B2(n_1287), .C(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g721 ( .A(n_4), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g741 ( .A1(n_4), .A2(n_58), .B1(n_405), .B2(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_5), .A2(n_64), .B1(n_583), .B2(n_1000), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_5), .A2(n_46), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_6), .A2(n_202), .B1(n_506), .B2(n_710), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_6), .A2(n_232), .B1(n_399), .B2(n_470), .Y(n_773) );
INVx1_ASAP7_75t_L g857 ( .A(n_7), .Y(n_857) );
AO22x1_ASAP7_75t_L g893 ( .A1(n_7), .A2(n_139), .B1(n_331), .B2(n_359), .Y(n_893) );
INVx1_ASAP7_75t_L g259 ( .A(n_8), .Y(n_259) );
AND2x2_ASAP7_75t_L g298 ( .A(n_8), .B(n_208), .Y(n_298) );
AND2x2_ASAP7_75t_L g334 ( .A(n_8), .B(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_8), .B(n_269), .Y(n_891) );
INVx1_ASAP7_75t_L g867 ( .A(n_9), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_9), .A2(n_92), .B1(n_350), .B2(n_389), .Y(n_892) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_10), .B(n_1055), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_10), .B(n_98), .Y(n_1057) );
INVx2_ASAP7_75t_L g1061 ( .A(n_10), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_11), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_12), .A2(n_79), .B1(n_467), .B2(n_609), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_13), .A2(n_210), .B1(n_851), .B2(n_1256), .Y(n_1255) );
INVxp67_ASAP7_75t_SL g1305 ( .A(n_13), .Y(n_1305) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_14), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g491 ( .A(n_15), .Y(n_491) );
INVx1_ASAP7_75t_L g646 ( .A(n_16), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_17), .A2(n_63), .B1(n_623), .B2(n_624), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_17), .A2(n_243), .B1(n_500), .B2(n_501), .C(n_502), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_18), .A2(n_159), .B1(n_1056), .B2(n_1062), .Y(n_1094) );
INVx1_ASAP7_75t_L g340 ( .A(n_19), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_19), .A2(n_158), .B1(n_405), .B2(n_411), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_20), .A2(n_48), .B1(n_365), .B2(n_369), .C(n_375), .Y(n_364) );
INVx1_ASAP7_75t_L g443 ( .A(n_20), .Y(n_443) );
INVx1_ASAP7_75t_L g645 ( .A(n_21), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g798 ( .A1(n_22), .A2(n_514), .B(n_799), .C(n_801), .Y(n_798) );
INVx1_ASAP7_75t_L g833 ( .A(n_22), .Y(n_833) );
XNOR2xp5_ASAP7_75t_L g1318 ( .A(n_23), .B(n_1319), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_24), .A2(n_184), .B1(n_1052), .B2(n_1059), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_25), .A2(n_85), .B1(n_467), .B2(n_609), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_26), .A2(n_243), .B1(n_623), .B2(n_624), .Y(n_633) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_26), .A2(n_63), .B1(n_361), .B2(n_652), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g1371 ( .A1(n_27), .A2(n_235), .B1(n_1372), .B2(n_1376), .Y(n_1371) );
OAI22xp33_ASAP7_75t_L g1410 ( .A1(n_27), .A2(n_235), .B1(n_1411), .B2(n_1414), .Y(n_1410) );
NAND2xp5_ASAP7_75t_SL g952 ( .A(n_28), .B(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_28), .A2(n_150), .B1(n_472), .B2(n_976), .Y(n_975) );
XNOR2xp5_ASAP7_75t_L g746 ( .A(n_29), .B(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_30), .A2(n_150), .B1(n_331), .B2(n_505), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_30), .A2(n_221), .B1(n_422), .B2(n_472), .Y(n_970) );
INVx1_ASAP7_75t_L g704 ( .A(n_31), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g1081 ( .A1(n_32), .A2(n_191), .B1(n_1052), .B2(n_1062), .Y(n_1081) );
AOI22xp5_ASAP7_75t_L g1091 ( .A1(n_33), .A2(n_103), .B1(n_1052), .B2(n_1059), .Y(n_1091) );
XOR2x2_ASAP7_75t_L g531 ( .A(n_34), .B(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_35), .A2(n_155), .B1(n_506), .B2(n_716), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g775 ( .A1(n_35), .A2(n_118), .B1(n_414), .B2(n_735), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g1093 ( .A1(n_36), .A2(n_84), .B1(n_1052), .B2(n_1059), .Y(n_1093) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_37), .A2(n_500), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g684 ( .A(n_37), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_38), .A2(n_57), .B1(n_505), .B2(n_665), .Y(n_792) );
AOI22xp33_ASAP7_75t_SL g812 ( .A1(n_38), .A2(n_240), .B1(n_623), .B2(n_624), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_39), .A2(n_127), .B1(n_480), .B2(n_1006), .Y(n_1005) );
INVxp67_ASAP7_75t_SL g1038 ( .A(n_39), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g1258 ( .A1(n_40), .A2(n_108), .B1(n_1003), .B2(n_1259), .C(n_1260), .Y(n_1258) );
INVx1_ASAP7_75t_L g1289 ( .A(n_40), .Y(n_1289) );
INVx1_ASAP7_75t_L g287 ( .A(n_41), .Y(n_287) );
INVx1_ASAP7_75t_L g321 ( .A(n_41), .Y(n_321) );
INVxp67_ASAP7_75t_SL g277 ( .A(n_42), .Y(n_277) );
AND4x1_ASAP7_75t_L g452 ( .A(n_42), .B(n_279), .C(n_327), .D(n_396), .Y(n_452) );
INVx1_ASAP7_75t_L g607 ( .A(n_43), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_44), .A2(n_185), .B1(n_522), .B2(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g685 ( .A(n_44), .Y(n_685) );
INVx1_ASAP7_75t_L g936 ( .A(n_45), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_46), .A2(n_135), .B1(n_583), .B2(n_1003), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g1269 ( .A1(n_47), .A2(n_81), .B1(n_583), .B2(n_1270), .C(n_1271), .Y(n_1269) );
INVx1_ASAP7_75t_L g1298 ( .A(n_47), .Y(n_1298) );
INVx1_ASAP7_75t_L g447 ( .A(n_48), .Y(n_447) );
INVx1_ASAP7_75t_L g253 ( .A(n_49), .Y(n_253) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_50), .A2(n_212), .B1(n_502), .B2(n_547), .C(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_50), .A2(n_242), .B1(n_399), .B2(n_623), .Y(n_686) );
INVx2_ASAP7_75t_L g293 ( .A(n_51), .Y(n_293) );
INVx1_ASAP7_75t_L g925 ( .A(n_52), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_53), .A2(n_73), .B1(n_1059), .B2(n_1066), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g538 ( .A1(n_54), .A2(n_114), .B1(n_356), .B2(n_388), .C(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g592 ( .A(n_54), .Y(n_592) );
INVx1_ASAP7_75t_L g1010 ( .A(n_55), .Y(n_1010) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_56), .A2(n_182), .B1(n_501), .B2(n_502), .C(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g816 ( .A1(n_57), .A2(n_88), .B1(n_623), .B2(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g718 ( .A(n_58), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_59), .A2(n_124), .B1(n_522), .B2(n_541), .Y(n_545) );
INVx1_ASAP7_75t_L g574 ( .A(n_59), .Y(n_574) );
INVx1_ASAP7_75t_L g978 ( .A(n_60), .Y(n_978) );
INVx1_ASAP7_75t_L g1273 ( .A(n_61), .Y(n_1273) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_62), .A2(n_167), .B1(n_470), .B2(n_472), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_62), .A2(n_214), .B1(n_361), .B2(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g1033 ( .A(n_64), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_65), .A2(n_123), .B1(n_1052), .B2(n_1059), .Y(n_1075) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_66), .A2(n_547), .B(n_676), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_66), .A2(n_160), .B1(n_734), .B2(n_735), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_67), .A2(n_193), .B1(n_304), .B2(n_315), .Y(n_303) );
OAI211xp5_ASAP7_75t_L g328 ( .A1(n_67), .A2(n_329), .B(n_336), .C(n_346), .Y(n_328) );
OAI211xp5_ASAP7_75t_L g702 ( .A1(n_68), .A2(n_365), .B(n_703), .C(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g729 ( .A(n_68), .Y(n_729) );
OAI222xp33_ASAP7_75t_L g877 ( .A1(n_69), .A2(n_192), .B1(n_878), .B2(n_880), .C1(n_882), .C2(n_884), .Y(n_877) );
INVx1_ASAP7_75t_L g897 ( .A(n_69), .Y(n_897) );
INVx1_ASAP7_75t_L g992 ( .A(n_70), .Y(n_992) );
OAI222xp33_ASAP7_75t_L g1026 ( .A1(n_70), .A2(n_120), .B1(n_369), .B2(n_536), .C1(n_1027), .C2(n_1034), .Y(n_1026) );
OAI22xp5_ASAP7_75t_SL g945 ( .A1(n_71), .A2(n_95), .B1(n_946), .B2(n_947), .Y(n_945) );
OAI21xp33_ASAP7_75t_L g960 ( .A1(n_71), .A2(n_742), .B(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g550 ( .A(n_72), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g1331 ( .A(n_74), .Y(n_1331) );
INVx1_ASAP7_75t_L g751 ( .A(n_75), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g1079 ( .A1(n_76), .A2(n_122), .B1(n_1052), .B2(n_1059), .Y(n_1079) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_77), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_78), .A2(n_237), .B1(n_359), .B2(n_361), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_78), .A2(n_106), .B1(n_425), .B2(n_428), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g758 ( .A1(n_79), .A2(n_497), .B(n_759), .C(n_762), .Y(n_758) );
AOI22xp5_ASAP7_75t_SL g1078 ( .A1(n_80), .A2(n_233), .B1(n_1062), .B2(n_1066), .Y(n_1078) );
AOI221xp5_ASAP7_75t_L g1286 ( .A1(n_81), .A2(n_179), .B1(n_1020), .B2(n_1287), .C(n_1288), .Y(n_1286) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_82), .Y(n_255) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_82), .B(n_253), .Y(n_1053) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_83), .A2(n_248), .B1(n_474), .B2(n_477), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g518 ( .A1(n_83), .A2(n_390), .B(n_519), .Y(n_518) );
OAI211xp5_ASAP7_75t_SL g711 ( .A1(n_85), .A2(n_329), .B(n_712), .C(n_717), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_86), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_87), .Y(n_671) );
AOI221xp5_ASAP7_75t_SL g795 ( .A1(n_88), .A2(n_240), .B1(n_350), .B2(n_354), .C(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_89), .A2(n_231), .B1(n_493), .B2(n_494), .Y(n_492) );
INVx1_ASAP7_75t_L g508 ( .A(n_89), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_90), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_91), .Y(n_632) );
INVx1_ASAP7_75t_L g863 ( .A(n_92), .Y(n_863) );
OAI211xp5_ASAP7_75t_L g939 ( .A1(n_93), .A2(n_940), .B(n_941), .C(n_942), .Y(n_939) );
INVxp33_ASAP7_75t_SL g962 ( .A(n_93), .Y(n_962) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_94), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_94), .A2(n_195), .B1(n_438), .B2(n_440), .Y(n_437) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_95), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_96), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g986 ( .A(n_97), .Y(n_986) );
INVx1_ASAP7_75t_L g1055 ( .A(n_98), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_98), .B(n_1061), .Y(n_1063) );
AOI22xp33_ASAP7_75t_SL g1090 ( .A1(n_99), .A2(n_105), .B1(n_1056), .B2(n_1062), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_100), .A2(n_241), .B1(n_1052), .B2(n_1056), .Y(n_1051) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_101), .Y(n_302) );
INVx1_ASAP7_75t_L g555 ( .A(n_102), .Y(n_555) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_104), .A2(n_149), .B1(n_1264), .B2(n_1267), .Y(n_1263) );
INVxp67_ASAP7_75t_SL g1307 ( .A(n_104), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_106), .A2(n_201), .B1(n_388), .B2(n_389), .C(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g616 ( .A(n_107), .Y(n_616) );
AOI21xp33_ASAP7_75t_L g650 ( .A1(n_107), .A2(n_390), .B(n_500), .Y(n_650) );
INVx1_ASAP7_75t_L g1296 ( .A(n_108), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_109), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g325 ( .A(n_109), .Y(n_325) );
INVx1_ASAP7_75t_L g436 ( .A(n_109), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g1343 ( .A(n_110), .Y(n_1343) );
AOI21xp33_ASAP7_75t_L g754 ( .A1(n_111), .A2(n_755), .B(n_756), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_111), .A2(n_155), .B1(n_734), .B2(n_735), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g1067 ( .A1(n_112), .A2(n_213), .B1(n_1052), .B2(n_1059), .Y(n_1067) );
OAI22xp33_ASAP7_75t_L g1381 ( .A1(n_113), .A2(n_161), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
OAI22xp33_ASAP7_75t_L g1389 ( .A1(n_113), .A2(n_161), .B1(n_1390), .B2(n_1393), .Y(n_1389) );
INVx1_ASAP7_75t_L g575 ( .A(n_114), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_115), .A2(n_134), .B1(n_707), .B2(n_799), .Y(n_808) );
INVx1_ASAP7_75t_L g820 ( .A(n_115), .Y(n_820) );
INVx1_ASAP7_75t_L g873 ( .A(n_116), .Y(n_873) );
NAND2xp33_ASAP7_75t_SL g915 ( .A(n_116), .B(n_350), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_117), .B(n_281), .Y(n_598) );
INVxp67_ASAP7_75t_SL g753 ( .A(n_118), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_119), .A2(n_209), .B1(n_315), .B2(n_609), .Y(n_608) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_119), .A2(n_497), .B(n_639), .C(n_644), .Y(n_638) );
INVx1_ASAP7_75t_L g990 ( .A(n_120), .Y(n_990) );
INVx1_ASAP7_75t_L g766 ( .A(n_121), .Y(n_766) );
INVx1_ASAP7_75t_L g587 ( .A(n_124), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g1332 ( .A(n_125), .Y(n_1332) );
OAI211xp5_ASAP7_75t_SL g1359 ( .A1(n_126), .A2(n_1354), .B(n_1360), .C(n_1363), .Y(n_1359) );
INVx1_ASAP7_75t_L g1409 ( .A(n_126), .Y(n_1409) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_127), .A2(n_236), .B1(n_356), .B2(n_1017), .C(n_1020), .Y(n_1016) );
OAI221xp5_ASAP7_75t_L g1254 ( .A1(n_128), .A2(n_180), .B1(n_875), .B2(n_882), .C(n_884), .Y(n_1254) );
OAI21xp33_ASAP7_75t_L g1282 ( .A1(n_128), .A2(n_905), .B(n_916), .Y(n_1282) );
INVx1_ASAP7_75t_L g764 ( .A(n_129), .Y(n_764) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_129), .A2(n_165), .B1(n_493), .B2(n_742), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g1339 ( .A(n_130), .Y(n_1339) );
INVx1_ASAP7_75t_L g668 ( .A(n_131), .Y(n_668) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_132), .Y(n_465) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_132), .A2(n_497), .B(n_498), .C(n_507), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_133), .A2(n_227), .B1(n_474), .B2(n_477), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_133), .A2(n_248), .B1(n_504), .B2(n_506), .Y(n_503) );
INVx1_ASAP7_75t_L g831 ( .A(n_134), .Y(n_831) );
INVx1_ASAP7_75t_L g1029 ( .A(n_135), .Y(n_1029) );
CKINVDCx16_ASAP7_75t_R g879 ( .A(n_136), .Y(n_879) );
NAND5xp2_ASAP7_75t_L g787 ( .A(n_137), .B(n_788), .C(n_810), .D(n_821), .E(n_828), .Y(n_787) );
INVx1_ASAP7_75t_L g837 ( .A(n_137), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g1073 ( .A1(n_137), .A2(n_223), .B1(n_1062), .B2(n_1074), .Y(n_1073) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_138), .A2(n_242), .B1(n_331), .B2(n_652), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_138), .A2(n_212), .B1(n_623), .B2(n_691), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_139), .A2(n_439), .B(n_579), .Y(n_874) );
INVx1_ASAP7_75t_L g919 ( .A(n_140), .Y(n_919) );
INVx1_ASAP7_75t_L g1261 ( .A(n_141), .Y(n_1261) );
INVx1_ASAP7_75t_L g667 ( .A(n_142), .Y(n_667) );
INVx1_ASAP7_75t_L g460 ( .A(n_143), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_143), .A2(n_145), .B1(n_370), .B2(n_511), .C(n_512), .Y(n_510) );
BUFx3_ASAP7_75t_L g286 ( .A(n_144), .Y(n_286) );
INVx1_ASAP7_75t_L g463 ( .A(n_145), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g1342 ( .A(n_146), .Y(n_1342) );
INVx1_ASAP7_75t_L g1253 ( .A(n_147), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_148), .A2(n_214), .B1(n_472), .B2(n_480), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g499 ( .A1(n_148), .A2(n_167), .B1(n_500), .B2(n_501), .C(n_502), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_149), .A2(n_180), .B1(n_896), .B2(n_1284), .Y(n_1283) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_151), .A2(n_232), .B1(n_356), .B2(n_501), .C(n_539), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_151), .A2(n_202), .B1(n_480), .B2(n_737), .Y(n_776) );
INVx1_ASAP7_75t_L g561 ( .A(n_152), .Y(n_561) );
OAI21xp33_ASAP7_75t_L g1008 ( .A1(n_153), .A2(n_304), .B(n_1009), .Y(n_1008) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_154), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_156), .A2(n_189), .B1(n_359), .B2(n_665), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_156), .A2(n_183), .B1(n_735), .B2(n_815), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g1367 ( .A(n_157), .Y(n_1367) );
INVx1_ASAP7_75t_L g337 ( .A(n_158), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_160), .A2(n_224), .B1(n_506), .B2(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g1011 ( .A(n_162), .Y(n_1011) );
CKINVDCx5p33_ASAP7_75t_R g1328 ( .A(n_163), .Y(n_1328) );
INVx1_ASAP7_75t_L g848 ( .A(n_164), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_164), .B(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g763 ( .A(n_165), .Y(n_763) );
INVx1_ASAP7_75t_L g995 ( .A(n_166), .Y(n_995) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_168), .A2(n_216), .B1(n_370), .B2(n_511), .C(n_670), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_168), .A2(n_216), .B1(n_462), .B2(n_635), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g1065 ( .A1(n_169), .A2(n_246), .B1(n_1062), .B2(n_1066), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_170), .A2(n_173), .B1(n_1056), .B2(n_1062), .Y(n_1108) );
AOI21xp33_ASAP7_75t_L g956 ( .A1(n_171), .A2(n_500), .B(n_756), .Y(n_956) );
INVx1_ASAP7_75t_L g967 ( .A(n_171), .Y(n_967) );
INVx1_ASAP7_75t_L g1368 ( .A(n_172), .Y(n_1368) );
OAI211xp5_ASAP7_75t_L g1396 ( .A1(n_172), .A2(n_1397), .B(n_1399), .C(n_1401), .Y(n_1396) );
OAI211xp5_ASAP7_75t_L g535 ( .A1(n_174), .A2(n_536), .B(n_537), .C(n_542), .Y(n_535) );
INVx1_ASAP7_75t_L g595 ( .A(n_174), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_175), .A2(n_228), .B1(n_501), .B2(n_547), .C(n_549), .Y(n_546) );
INVx1_ASAP7_75t_L g564 ( .A(n_175), .Y(n_564) );
INVx1_ASAP7_75t_L g827 ( .A(n_176), .Y(n_827) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_177), .Y(n_379) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_177), .A2(n_200), .B1(n_422), .B2(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g559 ( .A(n_178), .Y(n_559) );
OAI332xp33_ASAP7_75t_SL g562 ( .A1(n_178), .A2(n_405), .A3(n_563), .B1(n_569), .B2(n_572), .B3(n_578), .C1(n_580), .C2(n_586), .Y(n_562) );
INVx1_ASAP7_75t_L g1262 ( .A(n_179), .Y(n_1262) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_181), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_182), .A2(n_190), .B1(n_732), .B2(n_737), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_183), .A2(n_219), .B1(n_350), .B2(n_389), .C(n_756), .Y(n_793) );
XNOR2x1_ASAP7_75t_L g1248 ( .A(n_184), .B(n_1249), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_184), .A2(n_1315), .B1(n_1317), .B2(n_1421), .Y(n_1314) );
INVx1_ASAP7_75t_L g689 ( .A(n_185), .Y(n_689) );
XOR2x2_ASAP7_75t_L g931 ( .A(n_186), .B(n_932), .Y(n_931) );
AOI22xp33_ASAP7_75t_SL g950 ( .A1(n_187), .A2(n_229), .B1(n_331), .B2(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g969 ( .A(n_187), .Y(n_969) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_188), .Y(n_706) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_188), .A2(n_224), .B1(n_414), .B2(n_740), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_189), .A2(n_219), .B1(n_583), .B2(n_735), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_191), .B(n_456), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_191), .A2(n_487), .B1(n_488), .B2(n_525), .Y(n_486) );
INVx1_ASAP7_75t_L g527 ( .A(n_191), .Y(n_527) );
NOR2xp33_ASAP7_75t_R g904 ( .A(n_192), .B(n_905), .Y(n_904) );
OA22x2_ASAP7_75t_L g699 ( .A1(n_194), .A2(n_700), .B1(n_744), .B2(n_745), .Y(n_699) );
CKINVDCx16_ASAP7_75t_R g744 ( .A(n_194), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_195), .A2(n_200), .B1(n_348), .B2(n_352), .C(n_356), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g1326 ( .A(n_196), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_197), .A2(n_215), .B1(n_522), .B2(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g584 ( .A(n_197), .Y(n_584) );
INVx1_ASAP7_75t_L g842 ( .A(n_198), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_199), .A2(n_244), .B1(n_315), .B2(n_609), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_201), .A2(n_237), .B1(n_425), .B2(n_428), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_203), .A2(n_236), .B1(n_470), .B2(n_691), .Y(n_998) );
INVxp67_ASAP7_75t_SL g1035 ( .A(n_203), .Y(n_1035) );
INVx1_ASAP7_75t_L g694 ( .A(n_204), .Y(n_694) );
INVx1_ASAP7_75t_L g554 ( .A(n_205), .Y(n_554) );
OAI211xp5_ASAP7_75t_L g749 ( .A1(n_206), .A2(n_365), .B(n_750), .C(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g771 ( .A(n_206), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_207), .Y(n_944) );
BUFx3_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
INVx1_ASAP7_75t_L g335 ( .A(n_208), .Y(n_335) );
INVxp67_ASAP7_75t_SL g1277 ( .A(n_210), .Y(n_1277) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_211), .Y(n_802) );
INVx1_ASAP7_75t_L g566 ( .A(n_215), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g1336 ( .A(n_217), .Y(n_1336) );
INVx1_ASAP7_75t_L g291 ( .A(n_218), .Y(n_291) );
INVx1_ASAP7_75t_L g296 ( .A(n_218), .Y(n_296) );
INVx2_ASAP7_75t_L g395 ( .A(n_218), .Y(n_395) );
INVx1_ASAP7_75t_L g859 ( .A(n_220), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_220), .A2(n_247), .B1(n_359), .B2(n_665), .Y(n_914) );
NAND2xp5_ASAP7_75t_SL g949 ( .A(n_221), .B(n_500), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_222), .A2(n_226), .B1(n_1059), .B2(n_1062), .Y(n_1058) );
INVx1_ASAP7_75t_L g723 ( .A(n_225), .Y(n_723) );
INVx1_ASAP7_75t_L g513 ( .A(n_227), .Y(n_513) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_228), .Y(n_581) );
INVxp67_ASAP7_75t_SL g974 ( .A(n_229), .Y(n_974) );
OAI22xp33_ASAP7_75t_SL g634 ( .A1(n_230), .A2(n_238), .B1(n_462), .B2(n_635), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_230), .A2(n_238), .B1(n_365), .B2(n_370), .C(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g509 ( .A(n_231), .Y(n_509) );
XNOR2xp5_ASAP7_75t_L g604 ( .A(n_233), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g1041 ( .A(n_234), .Y(n_1041) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_239), .Y(n_943) );
OAI211xp5_ASAP7_75t_L g660 ( .A1(n_244), .A2(n_497), .B(n_661), .C(n_666), .Y(n_660) );
INVx1_ASAP7_75t_L g955 ( .A(n_245), .Y(n_955) );
INVx1_ASAP7_75t_L g869 ( .A(n_247), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_1044), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx1_ASAP7_75t_L g1313 ( .A(n_251), .Y(n_1313) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_252), .B(n_255), .Y(n_1316) );
INVx1_ASAP7_75t_L g1425 ( .A(n_252), .Y(n_1425) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1427 ( .A(n_255), .B(n_1425), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_258), .B(n_1313), .Y(n_1312) );
AND2x4_ASAP7_75t_L g1386 ( .A(n_258), .B(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g357 ( .A(n_259), .B(n_269), .Y(n_357) );
AND2x4_ASAP7_75t_L g391 ( .A(n_259), .B(n_268), .Y(n_391) );
AND2x4_ASAP7_75t_SL g1311 ( .A(n_260), .B(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1382 ( .A(n_260), .Y(n_1382) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
INVxp67_ASAP7_75t_L g1291 ( .A(n_262), .Y(n_1291) );
BUFx4f_ASAP7_75t_L g1297 ( .A(n_262), .Y(n_1297) );
OR2x6_ASAP7_75t_L g1374 ( .A(n_262), .B(n_1375), .Y(n_1374) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g378 ( .A(n_263), .Y(n_378) );
BUFx4f_ASAP7_75t_L g800 ( .A(n_263), .Y(n_800) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g300 ( .A(n_265), .Y(n_300) );
INVx1_ASAP7_75t_L g308 ( .A(n_265), .Y(n_308) );
INVx2_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
AND2x2_ASAP7_75t_L g344 ( .A(n_265), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g351 ( .A(n_265), .B(n_266), .Y(n_351) );
NAND2x1_ASAP7_75t_L g517 ( .A(n_265), .B(n_266), .Y(n_517) );
INVx1_ASAP7_75t_L g301 ( .A(n_266), .Y(n_301) );
AND2x2_ASAP7_75t_L g332 ( .A(n_266), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g345 ( .A(n_266), .Y(n_345) );
BUFx2_ASAP7_75t_L g373 ( .A(n_266), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_266), .B(n_333), .Y(n_385) );
OR2x2_ASAP7_75t_L g913 ( .A(n_266), .B(n_300), .Y(n_913) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g1362 ( .A(n_268), .Y(n_1362) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g1366 ( .A(n_269), .Y(n_1366) );
AND2x4_ASAP7_75t_L g1370 ( .A(n_269), .B(n_307), .Y(n_1370) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_780), .B2(n_781), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_600), .B2(n_779), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_529), .B1(n_530), .B2(n_599), .Y(n_274) );
INVx2_ASAP7_75t_L g599 ( .A(n_275), .Y(n_599) );
OAI22x1_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_453), .B1(n_454), .B2(n_528), .Y(n_275) );
INVx2_ASAP7_75t_L g528 ( .A(n_276), .Y(n_528) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B(n_452), .Y(n_276) );
NAND3xp33_ASAP7_75t_SL g278 ( .A(n_279), .B(n_327), .C(n_396), .Y(n_278) );
AOI21xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_302), .B(n_303), .Y(n_279) );
NAND2xp33_ASAP7_75t_L g484 ( .A(n_280), .B(n_485), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_280), .A2(n_607), .B(n_608), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_280), .A2(n_694), .B(n_695), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_280), .A2(n_723), .B(n_724), .Y(n_722) );
AOI21xp33_ASAP7_75t_L g765 ( .A1(n_280), .A2(n_766), .B(n_767), .Y(n_765) );
AOI211x1_ASAP7_75t_L g985 ( .A1(n_280), .A2(n_986), .B(n_987), .C(n_1008), .Y(n_985) );
INVx8_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_294), .Y(n_281) );
INVx1_ASAP7_75t_L g832 ( .A(n_282), .Y(n_832) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_288), .Y(n_282) );
INVx1_ASAP7_75t_L g568 ( .A(n_283), .Y(n_568) );
BUFx3_ASAP7_75t_L g585 ( .A(n_283), .Y(n_585) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_284), .Y(n_631) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g620 ( .A(n_285), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_286), .Y(n_314) );
INVx2_ASAP7_75t_L g318 ( .A(n_286), .Y(n_318) );
AND2x4_ASAP7_75t_L g400 ( .A(n_286), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g408 ( .A(n_286), .B(n_320), .Y(n_408) );
INVx1_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
INVx2_ASAP7_75t_L g401 ( .A(n_287), .Y(n_401) );
OR2x2_ASAP7_75t_L g310 ( .A(n_288), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g410 ( .A(n_288), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_288), .Y(n_413) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
OR2x2_ASAP7_75t_L g570 ( .A(n_289), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_SL g909 ( .A(n_289), .B(n_357), .Y(n_909) );
INVx1_ASAP7_75t_L g1301 ( .A(n_289), .Y(n_1301) );
HB1xp67_ASAP7_75t_L g1420 ( .A(n_289), .Y(n_1420) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g853 ( .A(n_292), .Y(n_853) );
INVx1_ASAP7_75t_L g1266 ( .A(n_292), .Y(n_1266) );
INVx3_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
BUFx3_ASAP7_75t_L g419 ( .A(n_293), .Y(n_419) );
NAND2xp33_ASAP7_75t_SL g571 ( .A(n_293), .B(n_325), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_294), .B(n_927), .Y(n_926) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x4_ASAP7_75t_L g402 ( .A(n_295), .B(n_322), .Y(n_402) );
INVx1_ASAP7_75t_L g1303 ( .A(n_295), .Y(n_1303) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g435 ( .A(n_296), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_296), .B(n_334), .Y(n_906) );
INVx1_ASAP7_75t_L g1304 ( .A(n_297), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_298), .B(n_307), .Y(n_306) );
AND2x6_ASAP7_75t_L g363 ( .A(n_298), .B(n_350), .Y(n_363) );
INVx1_ASAP7_75t_L g374 ( .A(n_298), .Y(n_374) );
AND2x2_ASAP7_75t_L g551 ( .A(n_298), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_298), .B(n_395), .Y(n_901) );
AND2x2_ASAP7_75t_L g339 ( .A(n_299), .B(n_334), .Y(n_339) );
INVx3_ASAP7_75t_L g360 ( .A(n_299), .Y(n_360) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_299), .Y(n_505) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_300), .Y(n_804) );
INVx2_ASAP7_75t_L g490 ( .A(n_304), .Y(n_490) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_310), .Y(n_304) );
AND2x4_ASAP7_75t_L g609 ( .A(n_305), .B(n_310), .Y(n_609) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
OR2x2_ASAP7_75t_L g896 ( .A(n_306), .B(n_309), .Y(n_896) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_L g326 ( .A(n_309), .Y(n_326) );
INVx1_ASAP7_75t_L g825 ( .A(n_309), .Y(n_825) );
INVx1_ASAP7_75t_L g1387 ( .A(n_309), .Y(n_1387) );
INVx2_ASAP7_75t_L g829 ( .A(n_310), .Y(n_829) );
INVx4_ASAP7_75t_L g577 ( .A(n_311), .Y(n_577) );
INVx3_ASAP7_75t_L g872 ( .A(n_311), .Y(n_872) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_L g591 ( .A(n_312), .Y(n_591) );
BUFx3_ASAP7_75t_L g1338 ( .A(n_312), .Y(n_1338) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
BUFx2_ASAP7_75t_L g1408 ( .A(n_313), .Y(n_1408) );
AND2x4_ASAP7_75t_L g429 ( .A(n_314), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g446 ( .A(n_314), .Y(n_446) );
BUFx2_ASAP7_75t_L g1405 ( .A(n_314), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_315), .B(n_921), .Y(n_920) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_326), .Y(n_315) );
OR2x6_ASAP7_75t_L g467 ( .A(n_316), .B(n_326), .Y(n_467) );
INVx2_ASAP7_75t_L g1252 ( .A(n_316), .Y(n_1252) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_317), .B(n_322), .Y(n_316) );
BUFx3_ASAP7_75t_L g422 ( .A(n_317), .Y(n_422) );
BUFx3_ASAP7_75t_L g439 ( .A(n_317), .Y(n_439) );
INVx8_ASAP7_75t_L g481 ( .A(n_317), .Y(n_481) );
HB1xp67_ASAP7_75t_L g976 ( .A(n_317), .Y(n_976) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_317), .B(n_1266), .Y(n_1265) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x4_ASAP7_75t_L g415 ( .A(n_318), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVxp67_ASAP7_75t_L g416 ( .A(n_321), .Y(n_416) );
INVx1_ASAP7_75t_L g876 ( .A(n_322), .Y(n_876) );
AND2x6_ASAP7_75t_L g883 ( .A(n_322), .B(n_445), .Y(n_883) );
AND2x2_ASAP7_75t_L g885 ( .A(n_322), .B(n_451), .Y(n_885) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND3x1_ASAP7_75t_L g434 ( .A(n_323), .B(n_435), .C(n_436), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g579 ( .A(n_323), .B(n_436), .Y(n_579) );
OR2x4_ASAP7_75t_L g1392 ( .A(n_323), .B(n_408), .Y(n_1392) );
INVx1_ASAP7_75t_L g1395 ( .A(n_323), .Y(n_1395) );
AND2x4_ASAP7_75t_L g1400 ( .A(n_323), .B(n_400), .Y(n_1400) );
OR2x6_ASAP7_75t_L g1415 ( .A(n_323), .B(n_620), .Y(n_1415) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND3x4_ASAP7_75t_L g418 ( .A(n_325), .B(n_419), .C(n_420), .Y(n_418) );
AND2x2_ASAP7_75t_L g864 ( .A(n_325), .B(n_419), .Y(n_864) );
HB1xp67_ASAP7_75t_L g1418 ( .A(n_325), .Y(n_1418) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_364), .B(n_392), .Y(n_327) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_SL g497 ( .A(n_330), .Y(n_497) );
NAND2xp5_ASAP7_75t_R g1025 ( .A(n_330), .B(n_995), .Y(n_1025) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_334), .Y(n_330) );
BUFx2_ASAP7_75t_L g541 ( .A(n_331), .Y(n_541) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g362 ( .A(n_332), .Y(n_362) );
BUFx3_ASAP7_75t_L g506 ( .A(n_332), .Y(n_506) );
BUFx3_ASAP7_75t_L g665 ( .A(n_332), .Y(n_665) );
AND2x4_ASAP7_75t_L g342 ( .A(n_334), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_SL g368 ( .A(n_334), .B(n_350), .Y(n_368) );
AND2x2_ASAP7_75t_L g556 ( .A(n_334), .B(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g807 ( .A(n_334), .Y(n_807) );
AND2x2_ASAP7_75t_L g826 ( .A(n_334), .B(n_343), .Y(n_826) );
HB1xp67_ASAP7_75t_L g1375 ( .A(n_335), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B1(n_340), .B2(n_341), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_338), .A2(n_342), .B1(n_508), .B2(n_509), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_338), .B(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_338), .A2(n_342), .B1(n_645), .B2(n_646), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_338), .A2(n_341), .B1(n_763), .B2(n_764), .Y(n_762) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_339), .A2(n_342), .B1(n_667), .B2(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g720 ( .A(n_339), .Y(n_720) );
AND2x4_ASAP7_75t_L g847 ( .A(n_339), .B(n_825), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_341), .A2(n_718), .B1(n_719), .B2(n_721), .Y(n_717) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_342), .A2(n_554), .B1(n_555), .B2(n_556), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_342), .A2(n_719), .B1(n_1010), .B2(n_1011), .Y(n_1014) );
INVx1_ASAP7_75t_L g548 ( .A(n_343), .Y(n_548) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_343), .Y(n_755) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g355 ( .A(n_344), .Y(n_355) );
BUFx3_ASAP7_75t_L g500 ( .A(n_344), .Y(n_500) );
AND2x4_ASAP7_75t_L g1384 ( .A(n_344), .B(n_1375), .Y(n_1384) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_358), .B(n_363), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_350), .Y(n_501) );
BUFx3_ASAP7_75t_L g663 ( .A(n_350), .Y(n_663) );
BUFx3_ASAP7_75t_L g953 ( .A(n_350), .Y(n_953) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_350), .B(n_1362), .Y(n_1361) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g1019 ( .A(n_351), .Y(n_1019) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g389 ( .A(n_355), .Y(n_389) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx4_ASAP7_75t_L g502 ( .A(n_357), .Y(n_502) );
INVx4_ASAP7_75t_L g796 ( .A(n_357), .Y(n_796) );
NAND4xp25_ASAP7_75t_L g948 ( .A(n_357), .B(n_949), .C(n_950), .D(n_952), .Y(n_948) );
AND2x4_ASAP7_75t_L g1299 ( .A(n_357), .B(n_1300), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_357), .B(n_1300), .Y(n_1357) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g522 ( .A(n_360), .Y(n_522) );
INVx2_ASAP7_75t_SL g652 ( .A(n_360), .Y(n_652) );
INVx1_ASAP7_75t_L g710 ( .A(n_360), .Y(n_710) );
INVx1_ASAP7_75t_L g951 ( .A(n_360), .Y(n_951) );
INVx2_ASAP7_75t_L g1022 ( .A(n_360), .Y(n_1022) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx3_ASAP7_75t_L g557 ( .A(n_362), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_363), .A2(n_499), .B(n_503), .Y(n_498) );
INVx1_ASAP7_75t_L g542 ( .A(n_363), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_363), .A2(n_640), .B(n_641), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_363), .A2(n_662), .B(n_664), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_363), .A2(n_713), .B(n_715), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_363), .A2(n_760), .B(n_761), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g1015 ( .A1(n_363), .A2(n_1016), .B(n_1021), .Y(n_1015) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g511 ( .A(n_366), .Y(n_511) );
INVx1_ASAP7_75t_L g536 ( .A(n_366), .Y(n_536) );
INVx4_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g937 ( .A(n_368), .Y(n_937) );
BUFx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g552 ( .A(n_373), .Y(n_552) );
INVx1_ASAP7_75t_L g903 ( .A(n_373), .Y(n_903) );
AND2x4_ASAP7_75t_L g1365 ( .A(n_373), .B(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g806 ( .A(n_374), .Y(n_806) );
OAI221xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_380), .B2(n_386), .C(n_387), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g1353 ( .A1(n_376), .A2(n_1332), .B1(n_1339), .B2(n_1354), .Y(n_1353) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx4_ASAP7_75t_L g947 ( .A(n_383), .Y(n_947) );
BUFx6f_ASAP7_75t_L g1040 ( .A(n_383), .Y(n_1040) );
INVx8_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_L g1292 ( .A(n_384), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1380 ( .A(n_384), .B(n_1366), .Y(n_1380) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g549 ( .A(n_391), .Y(n_549) );
INVx1_ASAP7_75t_L g676 ( .A(n_391), .Y(n_676) );
INVx3_ASAP7_75t_L g756 ( .A(n_391), .Y(n_756) );
OAI221xp5_ASAP7_75t_L g1027 ( .A1(n_391), .A2(n_1028), .B1(n_1029), .B2(n_1030), .C(n_1033), .Y(n_1027) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g524 ( .A(n_393), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_393), .B(n_928), .Y(n_927) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x6_ASAP7_75t_L g578 ( .A(n_394), .B(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g890 ( .A(n_394), .B(n_891), .Y(n_890) );
BUFx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
AND4x1_ASAP7_75t_L g396 ( .A(n_397), .B(n_403), .C(n_417), .D(n_442), .Y(n_396) );
AND5x1_ASAP7_75t_L g932 ( .A(n_397), .B(n_933), .C(n_963), .D(n_977), .E(n_981), .Y(n_932) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx3_ASAP7_75t_L g483 ( .A(n_398), .Y(n_483) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_398), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g680 ( .A(n_398), .B(n_681), .C(n_692), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_398), .B(n_726), .C(n_741), .Y(n_725) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_398), .A2(n_636), .B1(n_728), .B2(n_802), .C(n_820), .Y(n_819) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
INVx2_ASAP7_75t_L g441 ( .A(n_400), .Y(n_441) );
BUFx3_ASAP7_75t_L g472 ( .A(n_400), .Y(n_472) );
BUFx2_ASAP7_75t_L g624 ( .A(n_400), .Y(n_624) );
BUFx2_ASAP7_75t_L g737 ( .A(n_400), .Y(n_737) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_400), .B(n_1266), .Y(n_1268) );
INVx1_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
AND2x2_ASAP7_75t_L g444 ( .A(n_402), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g448 ( .A(n_402), .B(n_449), .Y(n_448) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_402), .B(n_445), .Y(n_462) );
AND2x4_ASAP7_75t_SL g636 ( .A(n_402), .B(n_449), .Y(n_636) );
AND2x4_ASAP7_75t_SL g728 ( .A(n_402), .B(n_445), .Y(n_728) );
AND2x2_ASAP7_75t_L g991 ( .A(n_402), .B(n_445), .Y(n_991) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_405), .B(n_980), .Y(n_979) );
OR2x6_ASAP7_75t_L g405 ( .A(n_406), .B(n_409), .Y(n_405) );
OR2x2_ASAP7_75t_L g493 ( .A(n_406), .B(n_409), .Y(n_493) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx3_ASAP7_75t_L g573 ( .A(n_408), .Y(n_573) );
BUFx3_ASAP7_75t_L g588 ( .A(n_408), .Y(n_588) );
BUFx4f_ASAP7_75t_L g856 ( .A(n_408), .Y(n_856) );
OR2x4_ASAP7_75t_L g1413 ( .A(n_408), .B(n_1395), .Y(n_1413) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g743 ( .A(n_410), .B(n_734), .Y(n_743) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g494 ( .A(n_412), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_412), .B(n_554), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_412), .A2(n_645), .B1(n_646), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_412), .A2(n_654), .B1(n_667), .B2(n_668), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_412), .A2(n_654), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
AND2x4_ASAP7_75t_L g654 ( .A(n_413), .B(n_655), .Y(n_654) );
AND2x4_ASAP7_75t_L g830 ( .A(n_413), .B(n_655), .Y(n_830) );
INVx3_ASAP7_75t_L g565 ( .A(n_414), .Y(n_565) );
INVx2_ASAP7_75t_SL g683 ( .A(n_414), .Y(n_683) );
BUFx8_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_415), .Y(n_427) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_415), .Y(n_476) );
INVx2_ASAP7_75t_L g615 ( .A(n_415), .Y(n_615) );
AOI33xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .A3(n_424), .B1(n_431), .B2(n_432), .B3(n_437), .Y(n_417) );
AOI33xp33_ASAP7_75t_L g468 ( .A1(n_418), .A2(n_469), .A3(n_473), .B1(n_478), .B2(n_479), .B3(n_482), .Y(n_468) );
AOI33xp33_ASAP7_75t_L g730 ( .A1(n_418), .A2(n_731), .A3(n_733), .B1(n_736), .B2(n_738), .B3(n_739), .Y(n_730) );
AOI33xp33_ASAP7_75t_L g772 ( .A1(n_418), .A2(n_738), .A3(n_773), .B1(n_774), .B2(n_775), .B3(n_776), .Y(n_772) );
AOI33xp33_ASAP7_75t_L g811 ( .A1(n_418), .A2(n_812), .A3(n_813), .B1(n_814), .B2(n_816), .B3(n_818), .Y(n_811) );
BUFx3_ASAP7_75t_L g997 ( .A(n_418), .Y(n_997) );
INVx3_ASAP7_75t_L g1404 ( .A(n_419), .Y(n_1404) );
INVx1_ASAP7_75t_L g679 ( .A(n_420), .Y(n_679) );
OAI31xp33_ASAP7_75t_L g849 ( .A1(n_420), .A2(n_850), .A3(n_854), .B(n_877), .Y(n_849) );
INVx2_ASAP7_75t_SL g471 ( .A(n_422), .Y(n_471) );
BUFx3_ASAP7_75t_L g732 ( .A(n_422), .Y(n_732) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_426), .A2(n_868), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_427), .Y(n_583) );
INVx2_ASAP7_75t_L g628 ( .A(n_427), .Y(n_628) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_427), .Y(n_815) );
AND2x4_ASAP7_75t_L g1394 ( .A(n_427), .B(n_1395), .Y(n_1394) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g477 ( .A(n_429), .Y(n_477) );
BUFx12f_ASAP7_75t_L g735 ( .A(n_429), .Y(n_735) );
BUFx3_ASAP7_75t_L g740 ( .A(n_429), .Y(n_740) );
AND2x4_ASAP7_75t_L g928 ( .A(n_429), .B(n_853), .Y(n_928) );
INVx5_ASAP7_75t_L g1001 ( .A(n_429), .Y(n_1001) );
INVx1_ASAP7_75t_L g451 ( .A(n_430), .Y(n_451) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g482 ( .A(n_433), .Y(n_482) );
BUFx2_ASAP7_75t_L g1004 ( .A(n_433), .Y(n_1004) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g626 ( .A(n_434), .Y(n_626) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g691 ( .A(n_441), .Y(n_691) );
INVx2_ASAP7_75t_L g817 ( .A(n_441), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_447), .B2(n_448), .Y(n_442) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_448), .A2(n_460), .B1(n_461), .B2(n_463), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_448), .A2(n_461), .B1(n_550), .B2(n_595), .Y(n_594) );
AOI221x1_ASAP7_75t_L g963 ( .A1(n_448), .A2(n_461), .B1(n_936), .B2(n_943), .C(n_964), .Y(n_963) );
AO22x1_ASAP7_75t_L g989 ( .A1(n_448), .A2(n_990), .B1(n_991), .B2(n_992), .Y(n_989) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g454 ( .A(n_455), .B(n_486), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_484), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_SL g525 ( .A(n_458), .B(n_526), .Y(n_525) );
NAND4xp25_ASAP7_75t_SL g458 ( .A(n_459), .B(n_464), .C(n_468), .D(n_483), .Y(n_458) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_466), .B(n_555), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_466), .B(n_982), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_466), .B(n_995), .Y(n_994) );
INVx5_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_SL g1259 ( .A(n_470), .Y(n_1259) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
INVx3_ASAP7_75t_L g862 ( .A(n_476), .Y(n_862) );
INVx2_ASAP7_75t_SL g866 ( .A(n_476), .Y(n_866) );
INVx5_ASAP7_75t_L g973 ( .A(n_476), .Y(n_973) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx8_ASAP7_75t_L g623 ( .A(n_481), .Y(n_623) );
INVx2_ASAP7_75t_L g655 ( .A(n_481), .Y(n_655) );
INVx1_ASAP7_75t_L g1340 ( .A(n_482), .Y(n_1340) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_483), .B(n_594), .C(n_596), .D(n_597), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g993 ( .A(n_483), .B(n_994), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_484), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_495), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_492), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_490), .A2(n_561), .B(n_562), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_510), .B(n_523), .Y(n_495) );
INVx1_ASAP7_75t_L g520 ( .A(n_500), .Y(n_520) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_500), .Y(n_714) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g643 ( .A(n_505), .Y(n_643) );
INVx1_ASAP7_75t_SL g1024 ( .A(n_506), .Y(n_1024) );
OAI211xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_518), .C(n_521), .Y(n_512) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g649 ( .A(n_515), .Y(n_649) );
INVx2_ASAP7_75t_L g941 ( .A(n_515), .Y(n_941) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx4f_ASAP7_75t_L g707 ( .A(n_516), .Y(n_707) );
OR2x6_ASAP7_75t_L g916 ( .A(n_516), .B(n_917), .Y(n_916) );
BUFx4f_ASAP7_75t_L g1028 ( .A(n_516), .Y(n_1028) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g674 ( .A(n_517), .Y(n_674) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g539 ( .A(n_520), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_523), .A2(n_535), .B(n_543), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_523), .A2(n_638), .B(n_647), .Y(n_637) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_523), .A2(n_702), .B(n_711), .Y(n_701) );
OAI21xp5_ASAP7_75t_SL g748 ( .A1(n_523), .A2(n_749), .B(n_758), .Y(n_748) );
OAI21xp5_ASAP7_75t_L g1012 ( .A1(n_523), .A2(n_1013), .B(n_1026), .Y(n_1012) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g1275 ( .A(n_524), .Y(n_1275) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_593), .C(n_598), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_560), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_553), .C(n_558), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_550), .B2(n_551), .Y(n_544) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_551), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_551), .B(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_552), .A2(n_802), .B1(n_803), .B2(n_805), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_552), .A2(n_803), .B1(n_943), .B2(n_944), .Y(n_942) );
INVx2_ASAP7_75t_L g790 ( .A(n_556), .Y(n_790) );
AND2x4_ASAP7_75t_L g922 ( .A(n_557), .B(n_923), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_566), .B2(n_567), .Y(n_563) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI22xp5_ASAP7_75t_SL g681 ( .A1(n_569), .A2(n_682), .B1(n_687), .B2(n_688), .Y(n_681) );
BUFx8_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx4f_ASAP7_75t_L g613 ( .A(n_570), .Y(n_613) );
BUFx2_ASAP7_75t_L g965 ( .A(n_570), .Y(n_965) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_575), .B2(n_576), .Y(n_572) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g738 ( .A(n_578), .Y(n_738) );
INVx1_ASAP7_75t_L g818 ( .A(n_578), .Y(n_818) );
INVx3_ASAP7_75t_L g1274 ( .A(n_579), .Y(n_1274) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B1(n_584), .B2(n_585), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g972 ( .A1(n_585), .A2(n_955), .B1(n_973), .B2(n_974), .C(n_975), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_589), .B2(n_592), .Y(n_586) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_588), .A2(n_871), .B1(n_1272), .B2(n_1273), .C(n_1274), .Y(n_1271) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g860 ( .A1(n_591), .A2(n_861), .B1(n_862), .B2(n_863), .C(n_864), .Y(n_860) );
OR2x6_ASAP7_75t_L g875 ( .A(n_591), .B(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g779 ( .A(n_600), .Y(n_779) );
AOI22x1_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_698), .B2(n_778), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AO22x2_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_656), .B1(n_657), .B2(n_697), .Y(n_603) );
INVx1_ASAP7_75t_L g697 ( .A(n_604), .Y(n_697) );
AND4x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_610), .C(n_637), .D(n_653), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .C(n_634), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_611), .B(n_769), .C(n_777), .Y(n_768) );
OAI22xp5_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_614), .B1(n_625), .B2(n_627), .Y(n_612) );
BUFx3_ASAP7_75t_L g1324 ( .A(n_613), .Y(n_1324) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B1(n_617), .B2(n_621), .C(n_622), .Y(n_614) );
INVx3_ASAP7_75t_L g734 ( .A(n_615), .Y(n_734) );
OR2x6_ASAP7_75t_SL g851 ( .A(n_615), .B(n_852), .Y(n_851) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_617), .A2(n_683), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_682) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_626), .Y(n_687) );
INVx2_ASAP7_75t_L g971 ( .A(n_626), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_630), .B2(n_632), .C(n_633), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g648 ( .A1(n_629), .A2(n_649), .B(n_650), .C(n_651), .Y(n_648) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_630), .A2(n_671), .B1(n_683), .B2(n_689), .C(n_690), .Y(n_688) );
CKINVDCx8_ASAP7_75t_R g630 ( .A(n_631), .Y(n_630) );
INVx3_ASAP7_75t_L g858 ( .A(n_631), .Y(n_858) );
INVx3_ASAP7_75t_L g868 ( .A(n_631), .Y(n_868) );
INVx3_ASAP7_75t_L g968 ( .A(n_631), .Y(n_968) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_636), .A2(n_704), .B1(n_728), .B2(n_729), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_636), .A2(n_728), .B1(n_751), .B2(n_771), .Y(n_770) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g716 ( .A(n_643), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_655), .A2(n_817), .B1(n_846), .B2(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND4x1_ASAP7_75t_L g658 ( .A(n_659), .B(n_680), .C(n_693), .D(n_696), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_669), .B(n_678), .Y(n_659) );
OAI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_675), .C(n_677), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g954 ( .A1(n_672), .A2(n_955), .B(n_956), .C(n_957), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g1351 ( .A1(n_672), .A2(n_946), .B1(n_1331), .B2(n_1336), .Y(n_1351) );
INVx5_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g905 ( .A(n_674), .B(n_906), .Y(n_905) );
BUFx2_ASAP7_75t_SL g1354 ( .A(n_674), .Y(n_1354) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI21x1_ASAP7_75t_L g788 ( .A1(n_679), .A2(n_789), .B(n_809), .Y(n_788) );
BUFx2_ASAP7_75t_L g959 ( .A(n_679), .Y(n_959) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_683), .A2(n_864), .B1(n_871), .B2(n_1261), .C(n_1262), .Y(n_1260) );
INVx1_ASAP7_75t_L g778 ( .A(n_698), .Y(n_778) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_746), .Y(n_698) );
INVx1_ASAP7_75t_L g745 ( .A(n_700), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_722), .C(n_725), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B(n_708), .C(n_709), .Y(n_705) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_707), .A2(n_753), .B(n_754), .C(n_757), .Y(n_752) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .Y(n_726) );
BUFx2_ASAP7_75t_L g1003 ( .A(n_735), .Y(n_1003) );
INVx1_ASAP7_75t_L g1007 ( .A(n_737), .Y(n_1007) );
NAND2x1_ASAP7_75t_L g822 ( .A(n_742), .B(n_823), .Y(n_822) );
INVx2_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_765), .C(n_768), .Y(n_747) );
BUFx3_ASAP7_75t_L g1020 ( .A(n_755), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AO22x2_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_983), .B1(n_1042), .B2(n_1043), .Y(n_783) );
INVx1_ASAP7_75t_L g1042 ( .A(n_784), .Y(n_1042) );
XNOR2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_931), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_841), .B1(n_929), .B2(n_930), .Y(n_785) );
INVx1_ASAP7_75t_L g930 ( .A(n_786), .Y(n_930) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_834), .C(n_838), .Y(n_786) );
INVx1_ASAP7_75t_L g835 ( .A(n_788), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_797) );
INVx2_ASAP7_75t_SL g1348 ( .A(n_799), .Y(n_1348) );
INVx3_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx4_ASAP7_75t_L g940 ( .A(n_800), .Y(n_940) );
BUFx6f_ASAP7_75t_L g1037 ( .A(n_800), .Y(n_1037) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AOI222xp33_ASAP7_75t_L g828 ( .A1(n_805), .A2(n_829), .B1(n_830), .B2(n_831), .C1(n_832), .C2(n_833), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_806), .A2(n_807), .B1(n_939), .B2(n_945), .Y(n_938) );
INVx1_ASAP7_75t_L g836 ( .A(n_810), .Y(n_836) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_819), .Y(n_810) );
INVx1_ASAP7_75t_L g840 ( .A(n_821), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_827), .Y(n_821) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_824), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_845) );
INVx1_ASAP7_75t_L g1279 ( .A(n_824), .Y(n_1279) );
AND2x4_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
INVx1_ASAP7_75t_L g839 ( .A(n_828), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_829), .A2(n_832), .B1(n_944), .B2(n_962), .Y(n_961) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_836), .B(n_837), .Y(n_834) );
OAI21xp33_ASAP7_75t_L g838 ( .A1(n_837), .A2(n_839), .B(n_840), .Y(n_838) );
INVx1_ASAP7_75t_L g929 ( .A(n_841), .Y(n_929) );
XNOR2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_844), .B(n_886), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_849), .Y(n_844) );
INVx3_ASAP7_75t_L g980 ( .A(n_847), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_847), .B(n_1307), .Y(n_1306) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_853), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_860), .B1(n_865), .B2(n_870), .C(n_875), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_855) );
HB1xp67_ASAP7_75t_L g1327 ( .A(n_856), .Y(n_1327) );
OAI22xp33_ASAP7_75t_L g1341 ( .A1(n_858), .A2(n_1327), .B1(n_1342), .B2(n_1343), .Y(n_1341) );
OAI211xp5_ASAP7_75t_L g910 ( .A1(n_861), .A2(n_911), .B(n_914), .C(n_915), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_867), .B1(n_868), .B2(n_869), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g966 ( .A1(n_866), .A2(n_967), .B1(n_968), .B2(n_969), .C(n_970), .Y(n_966) );
OAI21xp5_ASAP7_75t_SL g870 ( .A1(n_871), .A2(n_873), .B(n_874), .Y(n_870) );
INVx3_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g1329 ( .A(n_872), .Y(n_1329) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_879), .A2(n_895), .B1(n_897), .B2(n_898), .Y(n_894) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx4_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx2_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NAND3xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_918), .C(n_924), .Y(n_886) );
NOR3xp33_ASAP7_75t_SL g887 ( .A(n_888), .B(n_904), .C(n_907), .Y(n_887) );
OAI21xp5_ASAP7_75t_SL g888 ( .A1(n_889), .A2(n_893), .B(n_894), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_892), .Y(n_889) );
HB1xp67_ASAP7_75t_L g1293 ( .A(n_890), .Y(n_1293) );
INVx4_ASAP7_75t_L g1345 ( .A(n_890), .Y(n_1345) );
INVx1_ASAP7_75t_SL g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_SL g898 ( .A(n_899), .Y(n_898) );
HB1xp67_ASAP7_75t_L g1284 ( .A(n_899), .Y(n_1284) );
NAND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_902), .Y(n_899) );
INVx1_ASAP7_75t_L g917 ( .A(n_900), .Y(n_917) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx2_ASAP7_75t_SL g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g923 ( .A(n_906), .Y(n_923) );
OAI21xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_910), .B(n_916), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
BUFx2_ASAP7_75t_L g946 ( .A(n_913), .Y(n_946) );
BUFx2_ASAP7_75t_L g1032 ( .A(n_913), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .Y(n_918) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AOI211xp5_ASAP7_75t_L g1281 ( .A1(n_922), .A2(n_1253), .B(n_1282), .C(n_1283), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_925), .B(n_926), .Y(n_924) );
INVx3_ASAP7_75t_L g1256 ( .A(n_928), .Y(n_1256) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_958), .B(n_960), .Y(n_933) );
NAND4xp25_ASAP7_75t_L g934 ( .A(n_935), .B(n_938), .C(n_948), .D(n_954), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_946), .A2(n_1328), .B1(n_1343), .B2(n_1349), .Y(n_1352) );
INVx2_ASAP7_75t_L g1350 ( .A(n_947), .Y(n_1350) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
OAI22xp5_ASAP7_75t_SL g964 ( .A1(n_965), .A2(n_966), .B1(n_971), .B2(n_972), .Y(n_964) );
INVx8_ASAP7_75t_L g1335 ( .A(n_973), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
INVx2_ASAP7_75t_L g1043 ( .A(n_983), .Y(n_1043) );
XOR2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_1041), .Y(n_983) );
NAND2xp5_ASAP7_75t_SL g984 ( .A(n_985), .B(n_1012), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_988), .B(n_996), .Y(n_987) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_993), .Y(n_988) );
AOI33xp33_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .A3(n_999), .B1(n_1002), .B2(n_1004), .B3(n_1005), .Y(n_996) );
INVx2_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx2_ASAP7_75t_R g1270 ( .A(n_1001), .Y(n_1270) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
NAND3xp33_ASAP7_75t_SL g1013 ( .A(n_1014), .B(n_1015), .C(n_1025), .Y(n_1013) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1018), .Y(n_1287) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_SL g1023 ( .A(n_1024), .Y(n_1023) );
INVx2_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx4_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1036), .B1(n_1038), .B2(n_1039), .Y(n_1034) );
INVx2_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx5_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
OAI221xp5_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1244), .B1(n_1247), .B2(n_1308), .C(n_1314), .Y(n_1044) );
NOR2xp33_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1199), .Y(n_1045) );
NAND3xp33_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1138), .C(n_1168), .Y(n_1046) );
AOI211xp5_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1068), .B(n_1101), .C(n_1118), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1048), .B(n_1142), .Y(n_1141) );
AOI322xp5_ASAP7_75t_L g1150 ( .A1(n_1048), .A2(n_1076), .A3(n_1099), .B1(n_1103), .B2(n_1146), .C1(n_1151), .C2(n_1154), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1064), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1049), .B(n_1180), .Y(n_1179) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1049), .B(n_1181), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1049), .B(n_1092), .Y(n_1236) );
INVx3_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1050), .B(n_1106), .Y(n_1105) );
INVx3_ASAP7_75t_L g1117 ( .A(n_1050), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1050), .B(n_1064), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1050), .B(n_1167), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1050), .B(n_1142), .Y(n_1185) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_1050), .B(n_1147), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1050), .B(n_1126), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1050), .B(n_1064), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1050), .B(n_1240), .Y(n_1239) );
AND2x4_ASAP7_75t_SL g1050 ( .A(n_1051), .B(n_1058), .Y(n_1050) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1052), .Y(n_1246) );
AND2x6_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1054), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1053), .B(n_1057), .Y(n_1056) );
AND2x4_ASAP7_75t_L g1059 ( .A(n_1053), .B(n_1060), .Y(n_1059) );
AND2x6_ASAP7_75t_L g1062 ( .A(n_1053), .B(n_1063), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1053), .B(n_1057), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1053), .B(n_1057), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g1424 ( .A(n_1054), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1055), .B(n_1061), .Y(n_1060) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1064), .B(n_1098), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1064), .B(n_1089), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1064), .B(n_1089), .Y(n_1181) );
OAI221xp5_ASAP7_75t_SL g1205 ( .A1(n_1064), .A2(n_1069), .B1(n_1206), .B2(n_1207), .C(n_1208), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1067), .Y(n_1064) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_1065), .B(n_1067), .Y(n_1104) );
A2O1A1Ixp33_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1083), .B(n_1087), .C(n_1095), .Y(n_1068) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1069), .B(n_1111), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1069), .B(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1070), .B(n_1099), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1076), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1071), .B(n_1084), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1071), .B(n_1121), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1071), .B(n_1152), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1071), .B(n_1176), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1071), .B(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1071), .B(n_1113), .Y(n_1233) );
CKINVDCx5p33_ASAP7_75t_R g1071 ( .A(n_1072), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1072), .B(n_1076), .Y(n_1100) );
NOR2xp33_ASAP7_75t_L g1123 ( .A(n_1072), .B(n_1092), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1148 ( .A(n_1072), .B(n_1080), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1072), .B(n_1113), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1072), .B(n_1092), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1072), .B(n_1176), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1075), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1073), .B(n_1075), .Y(n_1158) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1076), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1076), .B(n_1222), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1080), .Y(n_1076) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1077), .Y(n_1086) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1077), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1079), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1080), .B(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1080), .Y(n_1122) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1080), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1080), .B(n_1086), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
NOR2xp33_ASAP7_75t_L g1224 ( .A(n_1083), .B(n_1225), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1084), .B(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1085), .B(n_1132), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1086), .B(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1086), .Y(n_1176) );
INVxp33_ASAP7_75t_SL g1174 ( .A(n_1087), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1092), .Y(n_1087) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1088), .Y(n_1133) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1088), .Y(n_1202) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1089), .Y(n_1098) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1089), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1091), .Y(n_1089) );
INVx3_ASAP7_75t_L g1099 ( .A(n_1092), .Y(n_1099) );
INVx2_ASAP7_75t_L g1111 ( .A(n_1092), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1092), .B(n_1098), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1209 ( .A(n_1092), .B(n_1183), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1094), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1100), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1172 ( .A(n_1097), .B(n_1173), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1099), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1098), .B(n_1104), .Y(n_1103) );
NAND3xp33_ASAP7_75t_L g1127 ( .A(n_1099), .B(n_1106), .C(n_1112), .Y(n_1127) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1099), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1154 ( .A(n_1099), .B(n_1155), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1099), .B(n_1189), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1099), .B(n_1175), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1100), .B(n_1115), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1100), .B(n_1143), .Y(n_1149) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1100), .Y(n_1186) );
OAI21xp5_ASAP7_75t_L g1232 ( .A1(n_1100), .A2(n_1233), .B(n_1234), .Y(n_1232) );
OAI21xp33_ASAP7_75t_L g1101 ( .A1(n_1102), .A2(n_1112), .B(n_1114), .Y(n_1101) );
NAND3xp33_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1105), .C(n_1110), .Y(n_1102) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1103), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_1104), .A2(n_1172), .B1(n_1174), .B2(n_1175), .Y(n_1171) );
OAI211xp5_ASAP7_75t_L g1190 ( .A1(n_1104), .A2(n_1191), .B(n_1193), .C(n_1197), .Y(n_1190) );
INVx2_ASAP7_75t_L g1240 ( .A(n_1104), .Y(n_1240) );
OAI21xp33_ASAP7_75t_L g1200 ( .A1(n_1105), .A2(n_1201), .B(n_1205), .Y(n_1200) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1107), .Y(n_1116) );
OAI31xp33_ASAP7_75t_SL g1168 ( .A1(n_1107), .A2(n_1169), .A3(n_1178), .B(n_1190), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1109), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1110), .B(n_1140), .Y(n_1139) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NAND2xp5_ASAP7_75t_SL g1192 ( .A(n_1111), .B(n_1152), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1111), .B(n_1180), .Y(n_1231) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1115), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1117), .Y(n_1115) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1116), .Y(n_1135) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1117), .Y(n_1177) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1124), .B1(n_1125), .B2(n_1127), .C(n_1128), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1123), .Y(n_1120) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1121), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1121), .B(n_1158), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1123), .B(n_1152), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1206 ( .A(n_1123), .B(n_1137), .Y(n_1206) );
INVx2_ASAP7_75t_SL g1167 ( .A(n_1124), .Y(n_1167) );
OAI322xp33_ASAP7_75t_L g1156 ( .A1(n_1125), .A2(n_1157), .A3(n_1159), .B1(n_1160), .B2(n_1161), .C1(n_1163), .C2(n_1165), .Y(n_1156) );
CKINVDCx14_ASAP7_75t_R g1125 ( .A(n_1126), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1126), .B(n_1132), .Y(n_1195) );
NAND4xp25_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1131), .C(n_1134), .D(n_1136), .Y(n_1128) );
OAI21xp5_ASAP7_75t_L g1187 ( .A1(n_1129), .A2(n_1188), .B(n_1189), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1129), .B(n_1204), .Y(n_1226) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1133), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1132), .B(n_1148), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1132), .B(n_1167), .Y(n_1213) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1132), .B(n_1242), .Y(n_1241) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_1134), .A2(n_1139), .B1(n_1141), .B2(n_1144), .C(n_1156), .Y(n_1138) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
AOI221xp5_ASAP7_75t_L g1208 ( .A1(n_1136), .A2(n_1146), .B1(n_1152), .B2(n_1167), .C(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
OAI21xp33_ASAP7_75t_L g1145 ( .A1(n_1141), .A2(n_1146), .B(n_1148), .Y(n_1145) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1142), .Y(n_1207) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
NAND3xp33_ASAP7_75t_SL g1144 ( .A(n_1145), .B(n_1149), .C(n_1150), .Y(n_1144) );
CKINVDCx14_ASAP7_75t_R g1146 ( .A(n_1147), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1151), .B(n_1198), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1152), .B(n_1158), .Y(n_1164) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1155), .Y(n_1196) );
OAI21xp33_ASAP7_75t_L g1229 ( .A1(n_1155), .A2(n_1230), .B(n_1232), .Y(n_1229) );
OAI321xp33_ASAP7_75t_L g1178 ( .A1(n_1158), .A2(n_1179), .A3(n_1182), .B1(n_1184), .B2(n_1186), .C(n_1187), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1158), .B(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
CKINVDCx5p33_ASAP7_75t_R g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
AOI21xp33_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1171), .B(n_1177), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1173), .B(n_1183), .Y(n_1182) );
AOI211xp5_ASAP7_75t_L g1227 ( .A1(n_1180), .A2(n_1228), .B(n_1229), .C(n_1237), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_1180), .B(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1237 ( .A1(n_1184), .A2(n_1238), .B1(n_1241), .B2(n_1243), .Y(n_1237) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1189), .Y(n_1212) );
OAI21xp5_ASAP7_75t_L g1193 ( .A1(n_1194), .A2(n_1195), .B(n_1196), .Y(n_1193) );
NAND4xp25_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1210), .C(n_1223), .D(n_1227), .Y(n_1199) );
NOR2xp33_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1203), .Y(n_1201) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1207), .B(n_1221), .Y(n_1220) );
AOI211xp5_ASAP7_75t_L g1210 ( .A1(n_1211), .A2(n_1213), .B(n_1214), .C(n_1219), .Y(n_1210) );
AOI21xp33_ASAP7_75t_SL g1214 ( .A1(n_1215), .A2(n_1217), .B(n_1218), .Y(n_1214) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1215), .Y(n_1228) );
NOR2xp33_ASAP7_75t_L g1219 ( .A(n_1218), .B(n_1220), .Y(n_1219) );
NOR2xp33_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1226), .Y(n_1223) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
CKINVDCx20_ASAP7_75t_R g1244 ( .A(n_1245), .Y(n_1244) );
CKINVDCx20_ASAP7_75t_R g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1280), .Y(n_1249) );
A2O1A1Ixp33_ASAP7_75t_SL g1250 ( .A1(n_1251), .A2(n_1257), .B(n_1275), .C(n_1276), .Y(n_1250) );
AOI211xp5_ASAP7_75t_L g1251 ( .A1(n_1252), .A2(n_1253), .B(n_1254), .C(n_1255), .Y(n_1251) );
NOR3xp33_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1263), .C(n_1269), .Y(n_1257) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
OAI22xp33_ASAP7_75t_L g1288 ( .A1(n_1273), .A2(n_1289), .B1(n_1290), .B2(n_1292), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
NAND3xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1285), .C(n_1306), .Y(n_1280) );
AOI222xp33_ASAP7_75t_L g1285 ( .A1(n_1286), .A2(n_1293), .B1(n_1294), .B2(n_1299), .C1(n_1302), .C2(n_1305), .Y(n_1285) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
OAI22xp5_ASAP7_75t_L g1295 ( .A1(n_1292), .A2(n_1296), .B1(n_1297), .B2(n_1298), .Y(n_1295) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1304), .Y(n_1302) );
CKINVDCx20_ASAP7_75t_R g1308 ( .A(n_1309), .Y(n_1308) );
CKINVDCx20_ASAP7_75t_R g1309 ( .A(n_1310), .Y(n_1309) );
INVx3_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
HB1xp67_ASAP7_75t_SL g1315 ( .A(n_1316), .Y(n_1315) );
INVxp33_ASAP7_75t_SL g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
HB1xp67_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
NAND3xp33_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1358), .C(n_1388), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1344), .Y(n_1322) );
OAI33xp33_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1325), .A3(n_1330), .B1(n_1333), .B2(n_1340), .B3(n_1341), .Y(n_1323) );
OAI22xp33_ASAP7_75t_L g1325 ( .A1(n_1326), .A2(n_1327), .B1(n_1328), .B2(n_1329), .Y(n_1325) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_1326), .A2(n_1342), .B1(n_1347), .B2(n_1349), .Y(n_1346) );
OAI22xp5_ASAP7_75t_L g1333 ( .A1(n_1334), .A2(n_1336), .B1(n_1337), .B2(n_1339), .Y(n_1333) );
INVx2_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx2_ASAP7_75t_L g1398 ( .A(n_1338), .Y(n_1398) );
OAI33xp33_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1346), .A3(n_1351), .B1(n_1352), .B2(n_1353), .B3(n_1355), .Y(n_1344) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx2_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
OAI31xp33_ASAP7_75t_SL g1358 ( .A1(n_1359), .A2(n_1371), .A3(n_1381), .B(n_1385), .Y(n_1358) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1367), .B1(n_1368), .B2(n_1369), .Y(n_1363) );
BUFx3_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1401 ( .A1(n_1367), .A2(n_1402), .B1(n_1406), .B2(n_1409), .Y(n_1401) );
BUFx3_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx2_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx2_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx3_ASAP7_75t_SL g1383 ( .A(n_1384), .Y(n_1383) );
BUFx3_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
OAI31xp33_ASAP7_75t_SL g1388 ( .A1(n_1389), .A2(n_1396), .A3(n_1410), .B(n_1416), .Y(n_1388) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
INVx2_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
CKINVDCx8_ASAP7_75t_R g1399 ( .A(n_1400), .Y(n_1399) );
BUFx3_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1405), .Y(n_1403) );
AND2x4_ASAP7_75t_L g1407 ( .A(n_1404), .B(n_1408), .Y(n_1407) );
BUFx6f_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx2_ASAP7_75t_SL g1412 ( .A(n_1413), .Y(n_1412) );
BUFx3_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1419), .Y(n_1416) );
INVx1_ASAP7_75t_SL g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx2_ASAP7_75t_SL g1421 ( .A(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
OAI21xp5_ASAP7_75t_L g1423 ( .A1(n_1424), .A2(n_1425), .B(n_1426), .Y(n_1423) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
endmodule