module fake_jpeg_19468_n_105 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_20),
.B1(n_15),
.B2(n_18),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_20),
.B1(n_15),
.B2(n_18),
.Y(n_41)
);

OR2x4_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_11),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_12),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_17),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_45),
.B(n_14),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_34),
.B1(n_10),
.B2(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_11),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_15),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_27),
.C(n_31),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_18),
.B1(n_19),
.B2(n_13),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_34),
.B1(n_13),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_34),
.B1(n_13),
.B2(n_31),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_52),
.B1(n_54),
.B2(n_53),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_60),
.B1(n_48),
.B2(n_41),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_31),
.B1(n_22),
.B2(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_64),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_40),
.B(n_45),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_69),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_1),
.B(n_2),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_49),
.B1(n_52),
.B2(n_58),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_50),
.C(n_57),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_80),
.C(n_62),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_71),
.B1(n_69),
.B2(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_9),
.Y(n_87)
);

OAI322xp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_14),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_1),
.C2(n_7),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_85),
.C(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_63),
.B(n_70),
.C(n_68),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_68),
.B1(n_4),
.B2(n_6),
.Y(n_84)
);

OAI221xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_77),
.C(n_80),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_1),
.B(n_4),
.Y(n_85)
);

OAI211xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_73),
.C(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_86),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_92),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_79),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_90),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_100),
.B(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_78),
.B1(n_76),
.B2(n_74),
.Y(n_102)
);

AOI221xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_99),
.B1(n_74),
.B2(n_76),
.C(n_9),
.Y(n_105)
);


endmodule