module fake_jpeg_11416_n_501 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_501);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_501;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_23),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_64),
.B(n_93),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_92),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_23),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_91),
.Y(n_154)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_29),
.B(n_3),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_94),
.B(n_98),
.Y(n_150)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_46),
.B1(n_39),
.B2(n_42),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_26),
.B(n_29),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_27),
.B1(n_18),
.B2(n_26),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_104),
.A2(n_122),
.B1(n_136),
.B2(n_31),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_115),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_20),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_59),
.A2(n_78),
.B1(n_75),
.B2(n_79),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_116),
.A2(n_118),
.B1(n_54),
.B2(n_91),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_54),
.A2(n_42),
.B1(n_46),
.B2(n_39),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_27),
.B1(n_18),
.B2(n_39),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_20),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_123),
.B(n_139),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_53),
.A2(n_27),
.B1(n_18),
.B2(n_46),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_148),
.B1(n_82),
.B2(n_84),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_55),
.A2(n_27),
.B1(n_44),
.B2(n_46),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_57),
.B(n_32),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_58),
.A2(n_63),
.B1(n_70),
.B2(n_80),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_69),
.C(n_90),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_168),
.C(n_118),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_85),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_170),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_49),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_158),
.A2(n_184),
.B(n_195),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_159),
.A2(n_173),
.B1(n_155),
.B2(n_183),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_113),
.A2(n_86),
.B1(n_93),
.B2(n_73),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g243 ( 
.A1(n_166),
.A2(n_36),
.B1(n_49),
.B2(n_48),
.Y(n_243)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_85),
.C(n_21),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_32),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_181),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_177),
.A2(n_184),
.B1(n_195),
.B2(n_196),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_28),
.B1(n_30),
.B2(n_45),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_130),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_190),
.Y(n_228)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_191),
.Y(n_230)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_194),
.Y(n_231)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_144),
.A2(n_28),
.B1(n_30),
.B2(n_45),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_146),
.A2(n_116),
.B1(n_126),
.B2(n_147),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_197),
.Y(n_212)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_200),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_119),
.B(n_28),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_199),
.B(n_208),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_122),
.A2(n_91),
.B1(n_30),
.B2(n_45),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_21),
.B1(n_31),
.B2(n_34),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_203),
.Y(n_245)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_204),
.Y(n_247)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_206),
.Y(n_214)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_149),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_137),
.B(n_49),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_255),
.C(n_206),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_117),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_216),
.B(n_236),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_220),
.A2(n_226),
.B1(n_241),
.B2(n_253),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_173),
.A2(n_117),
.B1(n_141),
.B2(n_129),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_168),
.B(n_137),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_158),
.A2(n_120),
.B(n_127),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_237),
.A2(n_34),
.B(n_188),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_238),
.A2(n_250),
.B1(n_5),
.B2(n_6),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_21),
.B(n_31),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_237),
.B(n_234),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_177),
.A2(n_141),
.B1(n_129),
.B2(n_127),
.Y(n_241)
);

AO22x2_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_14),
.B1(n_9),
.B2(n_10),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_166),
.A2(n_48),
.B1(n_41),
.B2(n_36),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_203),
.A2(n_48),
.B1(n_41),
.B2(n_36),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_169),
.B(n_97),
.C(n_41),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_219),
.B(n_192),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_256),
.B(n_261),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_191),
.B1(n_200),
.B2(n_157),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_257),
.A2(n_278),
.B1(n_296),
.B2(n_210),
.Y(n_307)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_209),
.A2(n_204),
.B1(n_186),
.B2(n_165),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_260),
.A2(n_265),
.B1(n_268),
.B2(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_269),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_202),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_264),
.B(n_281),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_196),
.B1(n_174),
.B2(n_178),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_266),
.A2(n_271),
.B(n_235),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_274),
.C(n_288),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_236),
.A2(n_179),
.B1(n_198),
.B2(n_143),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_275),
.Y(n_316)
);

OAI32xp33_ASAP7_75t_L g273 ( 
.A1(n_227),
.A2(n_167),
.A3(n_34),
.B1(n_207),
.B2(n_143),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_276),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_175),
.C(n_4),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_211),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_227),
.B(n_3),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_217),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_291),
.B1(n_295),
.B2(n_218),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_226),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_283),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_280),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_215),
.B(n_6),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_217),
.B(n_7),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_282),
.B(n_285),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_212),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_212),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_253),
.B1(n_248),
.B2(n_242),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_217),
.B(n_10),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_292),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_239),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_213),
.B(n_11),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_14),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_252),
.C(n_240),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_243),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_221),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_298),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_245),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_L g299 ( 
.A1(n_213),
.A2(n_12),
.B(n_13),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_SL g332 ( 
.A1(n_299),
.A2(n_229),
.B(n_246),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_300),
.B(n_304),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_263),
.A2(n_230),
.B1(n_247),
.B2(n_243),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_303),
.A2(n_315),
.B(n_319),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_292),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_307),
.A2(n_332),
.B1(n_334),
.B2(n_268),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_264),
.B(n_232),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_309),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_262),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_272),
.A2(n_243),
.B1(n_247),
.B2(n_218),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_313),
.A2(n_288),
.B1(n_298),
.B2(n_280),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_281),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_314),
.B(n_323),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_271),
.A2(n_233),
.B(n_252),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_223),
.C(n_235),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_322),
.C(n_324),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_286),
.B(n_223),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_321),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_249),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_279),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_249),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_328),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_260),
.A2(n_248),
.B1(n_254),
.B2(n_242),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_326),
.A2(n_296),
.B1(n_295),
.B2(n_256),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_259),
.B(n_240),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_244),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_270),
.C(n_289),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_258),
.A2(n_254),
.B(n_229),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_331),
.A2(n_291),
.B(n_272),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_265),
.A2(n_222),
.B1(n_210),
.B2(n_246),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_261),
.B(n_222),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_338),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_316),
.Y(n_339)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_303),
.A2(n_317),
.B(n_313),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_344),
.A2(n_350),
.B(n_354),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_337),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_311),
.Y(n_347)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_333),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_309),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_321),
.B(n_305),
.Y(n_351)
);

A2O1A1O1Ixp25_ASAP7_75t_L g354 ( 
.A1(n_319),
.A2(n_274),
.B(n_282),
.C(n_266),
.D(n_273),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_306),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_305),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_358),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_304),
.B(n_269),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_359),
.A2(n_312),
.B1(n_314),
.B2(n_325),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_360),
.A2(n_320),
.B(n_317),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_329),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_361),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_369),
.C(n_371),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_285),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_363),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_336),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_365),
.A2(n_312),
.B1(n_300),
.B2(n_323),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_322),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_367),
.Y(n_381)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_368),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_318),
.B(n_277),
.C(n_284),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_333),
.B(n_287),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_327),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_308),
.B(n_285),
.C(n_324),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_349),
.B(n_308),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_377),
.B(n_390),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_310),
.C(n_315),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_383),
.C(n_386),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_382),
.A2(n_393),
.B(n_360),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_335),
.C(n_330),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_343),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_387),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_358),
.Y(n_387)
);

NOR3xp33_ASAP7_75t_SL g388 ( 
.A(n_346),
.B(n_301),
.C(n_327),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_388),
.B(n_351),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_301),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_353),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_354),
.A2(n_320),
.B(n_336),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_331),
.C(n_326),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_399),
.C(n_369),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_396),
.A2(n_344),
.B1(n_348),
.B2(n_340),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_398),
.A2(n_340),
.B1(n_345),
.B2(n_363),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_367),
.B(n_338),
.C(n_285),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_408),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_379),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_416),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_357),
.Y(n_405)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_406),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_407),
.A2(n_350),
.B(n_373),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_353),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_398),
.A2(n_352),
.B1(n_359),
.B2(n_347),
.Y(n_409)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_410),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_352),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_423),
.Y(n_442)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_412),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_421),
.C(n_391),
.Y(n_440)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_414),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_376),
.B(n_361),
.CI(n_366),
.CON(n_416),
.SN(n_416)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_374),
.B1(n_344),
.B2(n_396),
.Y(n_427)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_420),
.Y(n_437)
);

FAx1_ASAP7_75t_SL g420 ( 
.A(n_376),
.B(n_341),
.CI(n_370),
.CON(n_420),
.SN(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_378),
.C(n_392),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_397),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_405),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_344),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_390),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_395),
.Y(n_435)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_427),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_407),
.A2(n_373),
.B(n_382),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_432),
.A2(n_414),
.B(n_397),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_433),
.A2(n_385),
.B(n_372),
.Y(n_453)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_434),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_436),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_393),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_399),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_439),
.B(n_440),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_391),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_413),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_438),
.A2(n_417),
.B1(n_406),
.B2(n_415),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_444),
.A2(n_457),
.B1(n_429),
.B2(n_427),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_425),
.A2(n_416),
.B(n_420),
.Y(n_445)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_445),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_434),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_448),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

BUFx5_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_450),
.B(n_454),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_452),
.A2(n_453),
.B(n_432),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_437),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_455),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_456),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_403),
.B1(n_385),
.B2(n_372),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_435),
.C(n_421),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_461),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_402),
.C(n_411),
.Y(n_461)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_463),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_465),
.B(n_453),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_451),
.A2(n_431),
.B1(n_430),
.B2(n_436),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_467),
.A2(n_381),
.B1(n_400),
.B2(n_433),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_402),
.C(n_443),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_468),
.B(n_469),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_408),
.C(n_442),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_444),
.A2(n_356),
.B1(n_339),
.B2(n_342),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_470),
.B(n_472),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_442),
.C(n_426),
.Y(n_472)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_475),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_450),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_478),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_459),
.B(n_458),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_426),
.C(n_439),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_479),
.B(n_461),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_471),
.A2(n_400),
.B1(n_457),
.B2(n_445),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_467),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_482),
.B(n_466),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_486),
.B(n_488),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

NOR2x1_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_460),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_474),
.A2(n_468),
.B(n_472),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_489),
.A2(n_476),
.B1(n_469),
.B2(n_479),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_490),
.B(n_483),
.C(n_418),
.Y(n_495)
);

OAI21xp33_ASAP7_75t_L g493 ( 
.A1(n_485),
.A2(n_480),
.B(n_481),
.Y(n_493)
);

O2A1O1Ixp33_ASAP7_75t_SL g494 ( 
.A1(n_493),
.A2(n_489),
.B(n_487),
.C(n_475),
.Y(n_494)
);

AO21x2_ASAP7_75t_L g497 ( 
.A1(n_494),
.A2(n_416),
.B(n_343),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_491),
.B(n_492),
.Y(n_496)
);

OAI321xp33_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_497),
.A3(n_356),
.B1(n_441),
.B2(n_368),
.C(n_355),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_498),
.B(n_389),
.C(n_365),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_420),
.B(n_418),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_285),
.Y(n_501)
);


endmodule