module fake_netlist_1_10053_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NOR2xp33_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
BUFx6f_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
NOR2xp33_ASAP7_75t_SL g6 ( .A(n_4), .B(n_0), .Y(n_6) );
BUFx2_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_5), .B(n_4), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_6), .Y(n_9) );
NOR2x1_ASAP7_75t_L g10 ( .A(n_9), .B(n_8), .Y(n_10) );
NAND3xp33_ASAP7_75t_SL g11 ( .A(n_9), .B(n_6), .C(n_8), .Y(n_11) );
NAND3xp33_ASAP7_75t_SL g12 ( .A(n_11), .B(n_0), .C(n_1), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_10), .B1(n_4), .B2(n_2), .Y(n_13) );
endmodule