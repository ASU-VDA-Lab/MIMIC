module fake_jpeg_14605_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_15),
.B(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_26),
.C(n_24),
.Y(n_43)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_21),
.C(n_15),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_55),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_17),
.B1(n_26),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_26),
.B1(n_35),
.B2(n_28),
.Y(n_84)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_41),
.B1(n_17),
.B2(n_37),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_79),
.B1(n_85),
.B2(n_63),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_36),
.B(n_20),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_19),
.C(n_25),
.Y(n_100)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_83),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_78),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_35),
.B1(n_37),
.B2(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_39),
.B1(n_16),
.B2(n_20),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_38),
.C(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_97),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_60),
.B1(n_55),
.B2(n_34),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_101),
.B1(n_107),
.B2(n_83),
.Y(n_125)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_43),
.B(n_34),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_24),
.C(n_38),
.Y(n_112)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_102),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_45),
.B1(n_54),
.B2(n_44),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_18),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_77),
.Y(n_120)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_54),
.B1(n_44),
.B2(n_47),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_33),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_112),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_103),
.Y(n_109)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_86),
.B(n_93),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_116),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_67),
.C(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_70),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_80),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_104),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_126),
.B(n_101),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_25),
.B(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_133),
.A2(n_150),
.B1(n_114),
.B2(n_110),
.Y(n_167)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_117),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_98),
.B1(n_101),
.B2(n_107),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_107),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_151),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_81),
.B(n_70),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_125),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_31),
.B(n_29),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_113),
.C(n_127),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_158),
.C(n_166),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_108),
.C(n_112),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_119),
.B1(n_109),
.B2(n_116),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_165),
.B1(n_169),
.B2(n_130),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_124),
.B(n_120),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_140),
.B1(n_143),
.B2(n_149),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_168),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_114),
.B1(n_110),
.B2(n_66),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_126),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_137),
.B(n_135),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_72),
.C(n_47),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_169)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_140),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_159),
.B(n_134),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_188),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_160),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_184),
.C(n_189),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_139),
.B1(n_147),
.B2(n_145),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_183),
.B1(n_171),
.B2(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_61),
.B(n_4),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_151),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_185),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_130),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_187),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_137),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_135),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_158),
.C(n_163),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_192),
.C(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_167),
.C(n_162),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_135),
.C(n_72),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_197),
.B1(n_31),
.B2(n_29),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_24),
.C(n_27),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_204),
.C(n_31),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_24),
.C(n_27),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_188),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_213),
.C(n_214),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_177),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_3),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_33),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_33),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_29),
.C(n_5),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_4),
.C(n_5),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_193),
.B1(n_192),
.B2(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_193),
.B(n_5),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_4),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_214),
.B(n_205),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_227),
.B(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_216),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_206),
.B1(n_210),
.B2(n_10),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_224),
.B1(n_225),
.B2(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_236),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_228),
.A2(n_219),
.B1(n_9),
.B2(n_10),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_235),
.A2(n_230),
.B1(n_13),
.B2(n_14),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_8),
.C(n_9),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_8),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

AOI21x1_ASAP7_75t_SL g239 ( 
.A1(n_234),
.A2(n_226),
.B(n_13),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_240),
.C(n_239),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_244),
.B(n_236),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_242),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_14),
.Y(n_247)
);


endmodule