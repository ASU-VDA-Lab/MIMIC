module real_jpeg_5022_n_15 (n_108, n_8, n_0, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_100, n_106, n_11, n_14, n_7, n_3, n_5, n_4, n_102, n_105, n_109, n_101, n_1, n_13, n_103, n_15);

input n_108;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_100;
input n_106;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_102;
input n_105;
input n_109;
input n_101;
input n_1;
input n_13;
input n_103;

output n_15;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_2),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_2),
.B(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_5),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_5),
.B(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_8),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_8),
.B(n_43),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_9),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_11),
.B(n_68),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_13),
.B(n_32),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_14),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_14),
.B(n_90),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_25),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_23),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B(n_97),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_88),
.B(n_94),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_81),
.B(n_87),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_76),
.B(n_80),
.Y(n_39)
);

AO221x1_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_51),
.B1(n_73),
.B2(n_74),
.C(n_75),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_54),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_78),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_72),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_55),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_67),
.B(n_71),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_66),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_100),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_101),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_102),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_103),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_104),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_105),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_106),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_107),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_108),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_109),
.Y(n_91)
);


endmodule