module real_aes_2329_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_759, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_760, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_759;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_760;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_358;
wire n_214;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g185 ( .A(n_0), .B(n_159), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_1), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_2), .B(n_143), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_3), .B(n_161), .Y(n_488) );
INVx1_ASAP7_75t_L g150 ( .A(n_4), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_5), .B(n_143), .Y(n_212) );
NAND2xp33_ASAP7_75t_SL g255 ( .A(n_6), .B(n_149), .Y(n_255) );
XNOR2xp5_ASAP7_75t_L g750 ( .A(n_7), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g247 ( .A(n_8), .Y(n_247) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_9), .Y(n_114) );
AND2x2_ASAP7_75t_L g210 ( .A(n_10), .B(n_167), .Y(n_210) );
AND2x2_ASAP7_75t_L g490 ( .A(n_11), .B(n_163), .Y(n_490) );
AND2x2_ASAP7_75t_L g500 ( .A(n_12), .B(n_253), .Y(n_500) );
INVx2_ASAP7_75t_L g165 ( .A(n_13), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_14), .B(n_161), .Y(n_540) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_15), .Y(n_115) );
AOI221x1_ASAP7_75t_L g250 ( .A1(n_16), .A2(n_152), .B1(n_251), .B2(n_253), .C(n_254), .Y(n_250) );
AOI22xp5_ASAP7_75t_SL g751 ( .A1(n_17), .A2(n_76), .B1(n_752), .B2(n_753), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_17), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_18), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_19), .B(n_143), .Y(n_545) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_20), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g127 ( .A(n_20), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_21), .A2(n_92), .B1(n_143), .B2(n_196), .Y(n_504) );
AOI221xp5_ASAP7_75t_SL g174 ( .A1(n_22), .A2(n_40), .B1(n_143), .B2(n_152), .C(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_23), .A2(n_152), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_24), .B(n_159), .Y(n_215) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_25), .A2(n_91), .B(n_165), .Y(n_164) );
OR2x2_ASAP7_75t_L g168 ( .A(n_25), .B(n_91), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_26), .B(n_161), .Y(n_160) );
INVxp67_ASAP7_75t_L g249 ( .A(n_27), .Y(n_249) );
AND2x2_ASAP7_75t_L g236 ( .A(n_28), .B(n_173), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_29), .A2(n_152), .B(n_184), .Y(n_183) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_30), .A2(n_253), .B(n_536), .Y(n_535) );
INVxp33_ASAP7_75t_L g756 ( .A(n_31), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_32), .B(n_161), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_33), .A2(n_73), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_33), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_34), .A2(n_152), .B(n_486), .Y(n_485) );
XOR2xp5_ASAP7_75t_L g749 ( .A(n_35), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_36), .B(n_161), .Y(n_560) );
AND2x2_ASAP7_75t_L g149 ( .A(n_37), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g153 ( .A(n_37), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g204 ( .A(n_37), .Y(n_204) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_38), .B(n_113), .C(n_115), .Y(n_112) );
OR2x6_ASAP7_75t_L g125 ( .A(n_38), .B(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_39), .A2(n_81), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_39), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_41), .B(n_143), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_42), .A2(n_84), .B1(n_152), .B2(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_43), .B(n_161), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_44), .B(n_143), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_45), .B(n_159), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_46), .A2(n_152), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g188 ( .A(n_47), .B(n_173), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_48), .B(n_159), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_49), .B(n_173), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_50), .B(n_143), .Y(n_537) );
INVx1_ASAP7_75t_L g146 ( .A(n_51), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_51), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_52), .B(n_161), .Y(n_498) );
AND2x2_ASAP7_75t_L g527 ( .A(n_53), .B(n_173), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_54), .B(n_143), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_55), .B(n_159), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_56), .B(n_159), .Y(n_559) );
AND2x2_ASAP7_75t_L g227 ( .A(n_57), .B(n_173), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_58), .B(n_143), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_59), .B(n_161), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_60), .B(n_143), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_61), .A2(n_152), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_62), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_63), .B(n_159), .Y(n_224) );
AND2x2_ASAP7_75t_L g551 ( .A(n_64), .B(n_167), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_65), .B(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_66), .A2(n_152), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_67), .B(n_161), .Y(n_216) );
AND2x2_ASAP7_75t_SL g207 ( .A(n_68), .B(n_163), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_69), .B(n_159), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_70), .B(n_159), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_71), .A2(n_94), .B1(n_152), .B2(n_202), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_72), .B(n_161), .Y(n_548) );
INVx1_ASAP7_75t_L g450 ( .A(n_73), .Y(n_450) );
INVx1_ASAP7_75t_L g148 ( .A(n_74), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_74), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_75), .B(n_159), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_76), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_77), .A2(n_152), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_78), .A2(n_152), .B(n_478), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_79), .A2(n_152), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g562 ( .A(n_80), .B(n_167), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_81), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_81), .B(n_173), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_82), .A2(n_86), .B1(n_143), .B2(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_83), .B(n_143), .Y(n_225) );
INVx1_ASAP7_75t_L g111 ( .A(n_85), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_87), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_88), .B(n_159), .Y(n_177) );
AND2x2_ASAP7_75t_L g481 ( .A(n_89), .B(n_163), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_90), .A2(n_152), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_93), .B(n_161), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_95), .A2(n_152), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_96), .B(n_161), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_97), .B(n_143), .Y(n_187) );
INVxp67_ASAP7_75t_L g252 ( .A(n_98), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_99), .B(n_161), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_100), .A2(n_152), .B(n_157), .Y(n_151) );
BUFx2_ASAP7_75t_L g550 ( .A(n_101), .Y(n_550) );
BUFx2_ASAP7_75t_SL g119 ( .A(n_102), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_102), .B(n_120), .C(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_103), .B(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_116), .B(n_755), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx3_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g757 ( .A(n_108), .Y(n_757) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_112), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_111), .B(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_115), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g461 ( .A(n_115), .B(n_125), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_115), .A2(n_135), .B1(n_464), .B2(n_465), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g464 ( .A(n_115), .Y(n_464) );
OA22x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_128), .B1(n_456), .B2(n_462), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
CKINVDCx8_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx2_ASAP7_75t_L g455 ( .A(n_123), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_124), .A2(n_463), .B(n_749), .C(n_754), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
AOI21xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_452), .B(n_454), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_133), .Y(n_129) );
INVx1_ASAP7_75t_L g453 ( .A(n_130), .Y(n_453) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp33_ASAP7_75t_SL g452 ( .A(n_134), .B(n_453), .Y(n_452) );
XNOR2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_449), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_341), .Y(n_135) );
NOR3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_269), .C(n_319), .Y(n_136) );
OAI211xp5_ASAP7_75t_SL g137 ( .A1(n_138), .A2(n_189), .B(n_237), .C(n_258), .Y(n_137) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_169), .Y(n_138) );
AND2x2_ASAP7_75t_L g268 ( .A(n_139), .B(n_170), .Y(n_268) );
INVx1_ASAP7_75t_L g399 ( .A(n_139), .Y(n_399) );
NOR2x1p5_ASAP7_75t_L g431 ( .A(n_139), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g242 ( .A(n_140), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g290 ( .A(n_140), .Y(n_290) );
OR2x2_ASAP7_75t_L g294 ( .A(n_140), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_140), .B(n_172), .Y(n_306) );
OR2x2_ASAP7_75t_L g328 ( .A(n_140), .B(n_172), .Y(n_328) );
AND2x4_ASAP7_75t_L g334 ( .A(n_140), .B(n_298), .Y(n_334) );
OR2x2_ASAP7_75t_L g351 ( .A(n_140), .B(n_244), .Y(n_351) );
INVx1_ASAP7_75t_L g386 ( .A(n_140), .Y(n_386) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_140), .Y(n_408) );
OR2x2_ASAP7_75t_L g422 ( .A(n_140), .B(n_355), .Y(n_422) );
AND2x4_ASAP7_75t_SL g426 ( .A(n_140), .B(n_244), .Y(n_426) );
OR2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_166), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_151), .B(n_163), .Y(n_141) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g256 ( .A(n_144), .Y(n_256) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
AND2x6_ASAP7_75t_L g159 ( .A(n_145), .B(n_154), .Y(n_159) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g161 ( .A(n_147), .B(n_156), .Y(n_161) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
AND2x2_ASAP7_75t_L g155 ( .A(n_150), .B(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_150), .Y(n_199) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
BUFx3_ASAP7_75t_L g200 ( .A(n_153), .Y(n_200) );
INVx2_ASAP7_75t_L g206 ( .A(n_154), .Y(n_206) );
AND2x4_ASAP7_75t_L g202 ( .A(n_155), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g198 ( .A(n_156), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_160), .B(n_162), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_159), .B(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_162), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_162), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_162), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_162), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_162), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_162), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_162), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_162), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_162), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_162), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_162), .A2(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_162), .A2(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_SL g193 ( .A(n_163), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_163), .A2(n_545), .B(n_546), .Y(n_544) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_165), .B(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g217 ( .A(n_165), .B(n_168), .Y(n_217) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_167), .Y(n_173) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g378 ( .A(n_170), .B(n_334), .Y(n_378) );
AND2x2_ASAP7_75t_L g425 ( .A(n_170), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_179), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g241 ( .A(n_172), .Y(n_241) );
AND2x2_ASAP7_75t_L g288 ( .A(n_172), .B(n_179), .Y(n_288) );
INVx2_ASAP7_75t_L g295 ( .A(n_172), .Y(n_295) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_172), .Y(n_416) );
BUFx3_ASAP7_75t_L g432 ( .A(n_172), .Y(n_432) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_178), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_173), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_173), .A2(n_476), .B(n_477), .Y(n_475) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_173), .A2(n_504), .B(n_505), .Y(n_503) );
INVx2_ASAP7_75t_L g257 ( .A(n_179), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_179), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g355 ( .A(n_179), .B(n_295), .Y(n_355) );
INVx1_ASAP7_75t_L g373 ( .A(n_179), .Y(n_373) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_179), .Y(n_389) );
INVx1_ASAP7_75t_L g411 ( .A(n_179), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_179), .B(n_290), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_179), .B(n_244), .Y(n_448) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21x1_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_188), .Y(n_180) );
INVx4_ASAP7_75t_L g253 ( .A(n_181), .Y(n_253) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_181), .A2(n_494), .B(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
INVx1_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_208), .Y(n_190) );
AND2x4_ASAP7_75t_L g262 ( .A(n_191), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g273 ( .A(n_191), .Y(n_273) );
AND2x2_ASAP7_75t_L g278 ( .A(n_191), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g313 ( .A(n_191), .B(n_218), .Y(n_313) );
AND2x2_ASAP7_75t_L g323 ( .A(n_191), .B(n_219), .Y(n_323) );
OR2x2_ASAP7_75t_L g403 ( .A(n_191), .B(n_318), .Y(n_403) );
OAI322xp33_ASAP7_75t_L g433 ( .A1(n_191), .A2(n_346), .A3(n_385), .B1(n_418), .B2(n_434), .C1(n_435), .C2(n_436), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_191), .B(n_416), .Y(n_434) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g267 ( .A(n_192), .Y(n_267) );
AOI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_207), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_201), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_196), .A2(n_202), .B1(n_246), .B2(n_248), .Y(n_245) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_200), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2x1p5_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_208), .A2(n_380), .B1(n_384), .B2(n_387), .Y(n_379) );
AOI211xp5_ASAP7_75t_L g439 ( .A1(n_208), .A2(n_440), .B(n_441), .C(n_444), .Y(n_439) );
AND2x4_ASAP7_75t_SL g208 ( .A(n_209), .B(n_218), .Y(n_208) );
AND2x4_ASAP7_75t_L g261 ( .A(n_209), .B(n_229), .Y(n_261) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
INVx5_ASAP7_75t_L g277 ( .A(n_209), .Y(n_277) );
INVx2_ASAP7_75t_L g286 ( .A(n_209), .Y(n_286) );
AND2x2_ASAP7_75t_L g309 ( .A(n_209), .B(n_219), .Y(n_309) );
AND2x2_ASAP7_75t_L g338 ( .A(n_209), .B(n_228), .Y(n_338) );
OR2x2_ASAP7_75t_L g347 ( .A(n_209), .B(n_267), .Y(n_347) );
OR2x2_ASAP7_75t_L g362 ( .A(n_209), .B(n_276), .Y(n_362) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_217), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_217), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_217), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_217), .B(n_252), .Y(n_251) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_217), .B(n_255), .C(n_256), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_217), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_217), .A2(n_537), .B(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_218), .B(n_238), .Y(n_237) );
INVx3_ASAP7_75t_SL g346 ( .A(n_218), .Y(n_346) );
AND2x2_ASAP7_75t_L g369 ( .A(n_218), .B(n_277), .Y(n_369) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
INVx2_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
AND2x2_ASAP7_75t_L g266 ( .A(n_219), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g280 ( .A(n_219), .B(n_229), .Y(n_280) );
INVx1_ASAP7_75t_L g284 ( .A(n_219), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_219), .B(n_229), .Y(n_318) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_219), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_219), .B(n_277), .Y(n_393) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_226), .B(n_227), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_225), .Y(n_220) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_226), .A2(n_230), .B(n_236), .Y(n_229) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_226), .A2(n_230), .B(n_236), .Y(n_276) );
AOI21x1_ASAP7_75t_L g483 ( .A1(n_226), .A2(n_484), .B(n_490), .Y(n_483) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_229), .Y(n_299) );
AND2x2_ASAP7_75t_L g383 ( .A(n_229), .B(n_267), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_242), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_239), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x6_ASAP7_75t_SL g447 ( .A(n_240), .B(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_241), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_241), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g395 ( .A(n_241), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_242), .A2(n_304), .B1(n_307), .B2(n_314), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_243), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_243), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_243), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_SL g394 ( .A(n_243), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_257), .Y(n_243) );
AND2x2_ASAP7_75t_L g289 ( .A(n_244), .B(n_290), .Y(n_289) );
INVx3_ASAP7_75t_L g298 ( .A(n_244), .Y(n_298) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_244), .A2(n_305), .B1(n_357), .B2(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g364 ( .A(n_244), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_244), .B(n_358), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_244), .B(n_288), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_244), .B(n_295), .Y(n_437) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
INVx3_ASAP7_75t_L g555 ( .A(n_253), .Y(n_555) );
OAI21xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_264), .B(n_268), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
NAND4xp25_ASAP7_75t_SL g307 ( .A(n_260), .B(n_308), .C(n_310), .D(n_312), .Y(n_307) );
INVx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_261), .B(n_368), .Y(n_397) );
AND2x2_ASAP7_75t_L g424 ( .A(n_261), .B(n_262), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_261), .B(n_284), .Y(n_435) );
INVx1_ASAP7_75t_L g300 ( .A(n_262), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_262), .A2(n_325), .B1(n_336), .B2(n_339), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_262), .B(n_275), .C(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_262), .B(n_277), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_262), .B(n_285), .Y(n_428) );
AND2x2_ASAP7_75t_L g360 ( .A(n_263), .B(n_267), .Y(n_360) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_263), .Y(n_421) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g316 ( .A(n_265), .Y(n_316) );
INVx1_ASAP7_75t_L g406 ( .A(n_266), .Y(n_406) );
AND2x2_ASAP7_75t_L g413 ( .A(n_266), .B(n_277), .Y(n_413) );
BUFx2_ASAP7_75t_L g368 ( .A(n_267), .Y(n_368) );
NAND3xp33_ASAP7_75t_SL g269 ( .A(n_270), .B(n_291), .C(n_303), .Y(n_269) );
OAI31xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_278), .A3(n_281), .B(n_287), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_271), .A2(n_325), .B1(n_329), .B2(n_330), .Y(n_324) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
OR2x2_ASAP7_75t_L g310 ( .A(n_273), .B(n_311), .Y(n_310) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_273), .B(n_337), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g405 ( .A1(n_274), .A2(n_376), .B(n_406), .C(n_407), .Y(n_405) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_275), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_276), .B(n_284), .Y(n_311) );
AND2x2_ASAP7_75t_L g329 ( .A(n_276), .B(n_309), .Y(n_329) );
AND2x2_ASAP7_75t_L g446 ( .A(n_279), .B(n_368), .Y(n_446) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g302 ( .A(n_280), .B(n_286), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_285), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g377 ( .A(n_285), .B(n_360), .Y(n_377) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_286), .B(n_360), .Y(n_366) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g358 ( .A(n_288), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_289), .B(n_389), .Y(n_388) );
AOI32xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_299), .A3(n_300), .B1(n_301), .B2(n_759), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_292), .A2(n_377), .B1(n_413), .B2(n_414), .C(n_417), .Y(n_412) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g305 ( .A(n_297), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g410 ( .A(n_298), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_299), .B(n_321), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_301), .A2(n_344), .B1(n_348), .B2(n_352), .C(n_356), .Y(n_343) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI211xp5_ASAP7_75t_L g319 ( .A1(n_306), .A2(n_320), .B(n_324), .C(n_335), .Y(n_319) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI322xp33_ASAP7_75t_L g417 ( .A1(n_312), .A2(n_322), .A3(n_371), .B1(n_418), .B2(n_419), .C1(n_420), .C2(n_422), .Y(n_417) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI21xp33_ASAP7_75t_L g444 ( .A1(n_315), .A2(n_445), .B(n_447), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_321), .A2(n_402), .B(n_404), .C(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g443 ( .A(n_328), .B(n_409), .Y(n_443) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVxp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_334), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g418 ( .A(n_334), .Y(n_418) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI31xp33_ASAP7_75t_L g374 ( .A1(n_338), .A2(n_375), .A3(n_377), .B(n_378), .Y(n_374) );
NOR2x1_ASAP7_75t_L g341 ( .A(n_342), .B(n_400), .Y(n_341) );
NAND5xp2_ASAP7_75t_L g342 ( .A(n_343), .B(n_363), .C(n_374), .D(n_379), .E(n_390), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AOI21xp33_ASAP7_75t_L g441 ( .A1(n_346), .A2(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g414 ( .A(n_350), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B(n_367), .C(n_370), .Y(n_363) );
INVxp33_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
OR2x2_ASAP7_75t_L g392 ( .A(n_368), .B(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_371), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g442 ( .A(n_383), .Y(n_442) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_394), .B(n_396), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_392), .A2(n_397), .B(n_398), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_401), .B(n_412), .C(n_423), .D(n_439), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_410), .B(n_431), .Y(n_430) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g440 ( .A(n_422), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_427), .B2(n_429), .C(n_433), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_463), .B(n_749), .Y(n_754) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_662), .Y(n_465) );
NOR4xp75_ASAP7_75t_L g466 ( .A(n_467), .B(n_585), .C(n_610), .D(n_637), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_522), .B(n_563), .Y(n_467) );
NOR4xp25_ASAP7_75t_L g468 ( .A(n_469), .B(n_506), .C(n_513), .D(n_517), .Y(n_468) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_491), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_473), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_473), .B(n_510), .Y(n_656) );
AND2x2_ASAP7_75t_L g681 ( .A(n_473), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g706 ( .A(n_473), .B(n_501), .Y(n_706) );
AND2x2_ASAP7_75t_L g747 ( .A(n_473), .B(n_515), .Y(n_747) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_SL g519 ( .A(n_474), .B(n_512), .Y(n_519) );
AND2x2_ASAP7_75t_L g521 ( .A(n_474), .B(n_493), .Y(n_521) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_474), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g582 ( .A(n_474), .Y(n_582) );
AND2x2_ASAP7_75t_L g588 ( .A(n_474), .B(n_515), .Y(n_588) );
BUFx2_ASAP7_75t_L g601 ( .A(n_474), .Y(n_601) );
AND2x4_ASAP7_75t_L g632 ( .A(n_474), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g679 ( .A(n_474), .B(n_680), .Y(n_679) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_481), .Y(n_474) );
INVx1_ASAP7_75t_L g673 ( .A(n_482), .Y(n_673) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx3_ASAP7_75t_L g512 ( .A(n_483), .Y(n_512) );
AND2x2_ASAP7_75t_L g515 ( .A(n_483), .B(n_493), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_489), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_491), .B(n_691), .Y(n_744) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
OR2x2_ASAP7_75t_L g581 ( .A(n_492), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
INVx2_ASAP7_75t_L g511 ( .A(n_493), .Y(n_511) );
INVx2_ASAP7_75t_L g572 ( .A(n_493), .Y(n_572) );
AND2x2_ASAP7_75t_L g682 ( .A(n_493), .B(n_512), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_499), .Y(n_494) );
INVx2_ASAP7_75t_L g570 ( .A(n_501), .Y(n_570) );
BUFx3_ASAP7_75t_L g587 ( .A(n_501), .Y(n_587) );
AND2x2_ASAP7_75t_L g614 ( .A(n_501), .B(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
AND2x4_ASAP7_75t_L g508 ( .A(n_502), .B(n_503), .Y(n_508) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx2_ASAP7_75t_L g516 ( .A(n_507), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_507), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g685 ( .A(n_507), .B(n_625), .Y(n_685) );
AND2x2_ASAP7_75t_L g709 ( .A(n_507), .B(n_519), .Y(n_709) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g605 ( .A(n_508), .B(n_511), .Y(n_605) );
AND2x2_ASAP7_75t_L g687 ( .A(n_508), .B(n_680), .Y(n_687) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_SL g730 ( .A(n_510), .Y(n_730) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g615 ( .A(n_511), .Y(n_615) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_512), .Y(n_619) );
INVx2_ASAP7_75t_L g627 ( .A(n_512), .Y(n_627) );
INVx1_ASAP7_75t_L g633 ( .A(n_512), .Y(n_633) );
AOI222xp33_ASAP7_75t_SL g563 ( .A1(n_513), .A2(n_564), .B1(n_568), .B2(n_573), .C1(n_580), .C2(n_583), .Y(n_563) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g640 ( .A(n_515), .Y(n_640) );
BUFx2_ASAP7_75t_L g669 ( .A(n_515), .Y(n_669) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_516), .A2(n_664), .B(n_668), .C(n_676), .Y(n_663) );
OR2x2_ASAP7_75t_L g734 ( .A(n_516), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g742 ( .A(n_516), .B(n_647), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_520), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_SL g699 ( .A(n_519), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g717 ( .A(n_519), .B(n_605), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_519), .B(n_697), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_520), .B(n_587), .Y(n_725) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g647 ( .A(n_521), .B(n_619), .Y(n_647) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_542), .Y(n_523) );
INVx1_ASAP7_75t_L g741 ( .A(n_524), .Y(n_741) );
NOR2xp67_ASAP7_75t_L g524 ( .A(n_525), .B(n_534), .Y(n_524) );
AND2x2_ASAP7_75t_L g584 ( .A(n_525), .B(n_543), .Y(n_584) );
INVx1_ASAP7_75t_L g661 ( .A(n_525), .Y(n_661) );
OR2x2_ASAP7_75t_L g720 ( .A(n_525), .B(n_543), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_525), .B(n_592), .Y(n_726) );
INVx4_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g567 ( .A(n_526), .Y(n_567) );
OR2x2_ASAP7_75t_L g599 ( .A(n_526), .B(n_553), .Y(n_599) );
AND2x2_ASAP7_75t_L g608 ( .A(n_526), .B(n_535), .Y(n_608) );
NAND2x1_ASAP7_75t_L g636 ( .A(n_526), .B(n_543), .Y(n_636) );
AND2x2_ASAP7_75t_L g683 ( .A(n_526), .B(n_578), .Y(n_683) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g566 ( .A(n_535), .Y(n_566) );
INVx1_ASAP7_75t_L g576 ( .A(n_535), .Y(n_576) );
AND2x2_ASAP7_75t_L g592 ( .A(n_535), .B(n_579), .Y(n_592) );
INVx2_ASAP7_75t_L g597 ( .A(n_535), .Y(n_597) );
OR2x2_ASAP7_75t_L g693 ( .A(n_535), .B(n_543), .Y(n_693) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_552), .Y(n_542) );
NOR2x1_ASAP7_75t_SL g578 ( .A(n_543), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g596 ( .A(n_543), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g609 ( .A(n_543), .B(n_553), .Y(n_609) );
BUFx2_ASAP7_75t_L g628 ( .A(n_543), .Y(n_628) );
INVx2_ASAP7_75t_SL g655 ( .A(n_543), .Y(n_655) );
OR2x6_ASAP7_75t_L g543 ( .A(n_544), .B(n_551), .Y(n_543) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g565 ( .A(n_553), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g711 ( .A(n_553), .B(n_653), .Y(n_711) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B(n_562), .Y(n_554) );
AO21x1_ASAP7_75t_SL g579 ( .A1(n_555), .A2(n_556), .B(n_562), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .Y(n_556) );
AOI211xp5_ASAP7_75t_L g727 ( .A1(n_564), .A2(n_588), .B(n_728), .C(n_732), .Y(n_727) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_565), .B(n_643), .Y(n_678) );
BUFx2_ASAP7_75t_L g642 ( .A(n_566), .Y(n_642) );
OR2x2_ASAP7_75t_L g590 ( .A(n_567), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g675 ( .A(n_567), .B(n_609), .Y(n_675) );
AND2x2_ASAP7_75t_L g696 ( .A(n_567), .B(n_652), .Y(n_696) );
INVx2_ASAP7_75t_L g703 ( .A(n_567), .Y(n_703) );
OAI21xp5_ASAP7_75t_SL g708 ( .A1(n_568), .A2(n_709), .B(n_710), .Y(n_708) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_L g650 ( .A(n_569), .B(n_632), .Y(n_650) );
OR2x2_ASAP7_75t_L g729 ( .A(n_569), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_570), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_572), .Y(n_603) );
AND2x2_ASAP7_75t_L g680 ( .A(n_572), .B(n_627), .Y(n_680) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
AND2x2_ASAP7_75t_L g665 ( .A(n_575), .B(n_666), .Y(n_665) );
AND2x4_ASAP7_75t_SL g674 ( .A(n_575), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_575), .B(n_584), .Y(n_707) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g583 ( .A(n_576), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g702 ( .A(n_577), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g652 ( .A(n_578), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g622 ( .A(n_579), .B(n_597), .Y(n_622) );
OAI31xp33_ASAP7_75t_L g629 ( .A1(n_580), .A2(n_630), .A3(n_632), .B(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_582), .B(n_605), .Y(n_631) );
AO21x1_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_589), .B(n_593), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g641 ( .A(n_587), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g746 ( .A(n_587), .Y(n_746) );
INVx2_ASAP7_75t_SL g731 ( .A(n_588), .Y(n_731) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g635 ( .A(n_591), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g719 ( .A(n_591), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_592), .B(n_655), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_600), .B1(n_604), .B2(n_606), .Y(n_593) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_594), .A2(n_713), .B(n_714), .Y(n_712) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_L g653 ( .A(n_597), .Y(n_653) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g667 ( .A(n_599), .B(n_628), .Y(n_667) );
OR2x2_ASAP7_75t_L g692 ( .A(n_599), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_601), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_601), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g691 ( .A(n_601), .Y(n_691) );
INVx2_ASAP7_75t_L g620 ( .A(n_602), .Y(n_620) );
INVx1_ASAP7_75t_L g700 ( .A(n_603), .Y(n_700) );
AND2x2_ASAP7_75t_L g623 ( .A(n_605), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g697 ( .A(n_605), .Y(n_697) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_611), .B(n_629), .Y(n_610) );
OAI321xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_616), .A3(n_621), .B1(n_622), .B2(n_623), .C(n_628), .Y(n_611) );
AOI322xp5_ASAP7_75t_L g737 ( .A1(n_612), .A2(n_643), .A3(n_738), .B1(n_740), .B2(n_742), .C1(n_743), .C2(n_748), .Y(n_737) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g690 ( .A(n_615), .Y(n_690) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_617), .B(n_697), .Y(n_714) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g722 ( .A(n_620), .Y(n_722) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp33_ASAP7_75t_SL g654 ( .A(n_622), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g721 ( .A1(n_625), .A2(n_631), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g643 ( .A(n_636), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_657), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_643), .B1(n_644), .B2(n_645), .C(n_648), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_640), .Y(n_659) );
AND2x2_ASAP7_75t_L g644 ( .A(n_642), .B(n_643), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp33_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_651), .B1(n_654), .B2(n_656), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g660 ( .A(n_652), .B(n_661), .Y(n_660) );
OAI21xp33_ASAP7_75t_L g743 ( .A1(n_655), .A2(n_744), .B(n_745), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR3xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_694), .C(n_715), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_667), .A2(n_702), .B1(n_729), .B2(n_731), .Y(n_728) );
OAI21xp33_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_670), .B(n_674), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_669), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_675), .A2(n_717), .B1(n_718), .B2(n_721), .C(n_723), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B1(n_681), .B2(n_683), .C(n_684), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g713 ( .A(n_679), .Y(n_713) );
INVx1_ASAP7_75t_L g735 ( .A(n_680), .Y(n_735) );
INVx1_ASAP7_75t_SL g733 ( .A(n_681), .Y(n_733) );
AOI31xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .A3(n_688), .B(n_692), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_685), .A2(n_695), .B1(n_697), .B2(n_698), .C(n_760), .Y(n_694) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B(n_704), .C(n_712), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g710 ( .A(n_703), .B(n_711), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g704 ( .A1(n_705), .A2(n_707), .B(n_708), .Y(n_704) );
INVx1_ASAP7_75t_L g739 ( .A(n_711), .Y(n_739) );
BUFx2_ASAP7_75t_SL g748 ( .A(n_711), .Y(n_748) );
NAND3xp33_ASAP7_75t_SL g715 ( .A(n_716), .B(n_727), .C(n_737), .Y(n_715) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI21xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B(n_726), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B(n_736), .Y(n_732) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
endmodule