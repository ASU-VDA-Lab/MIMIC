module real_jpeg_26144_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_0),
.B(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_0),
.B(n_75),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_0),
.B(n_57),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_0),
.B(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_0),
.B(n_29),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_0),
.B(n_25),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_0),
.B(n_54),
.Y(n_266)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_2),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_3),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_3),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_3),
.B(n_17),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_3),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_3),
.B(n_75),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_3),
.B(n_57),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_3),
.B(n_33),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_4),
.B(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_103),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_4),
.B(n_75),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_4),
.B(n_29),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_4),
.B(n_25),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_7),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_7),
.B(n_103),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_7),
.B(n_75),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_7),
.B(n_33),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_7),
.B(n_29),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_10),
.B(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_10),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_10),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_10),
.B(n_57),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_10),
.B(n_33),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_10),
.B(n_29),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_10),
.B(n_25),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_10),
.B(n_36),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_12),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_12),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_12),
.B(n_75),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_12),
.B(n_57),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_12),
.B(n_33),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_12),
.B(n_29),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_12),
.B(n_54),
.Y(n_337)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_14),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_14),
.B(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_14),
.B(n_75),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_14),
.B(n_57),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_14),
.B(n_33),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_29),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_14),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_14),
.B(n_54),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_33),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_15),
.B(n_103),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_15),
.B(n_75),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_15),
.B(n_57),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_16),
.B(n_57),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_16),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_16),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_16),
.B(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_16),
.B(n_29),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_16),
.B(n_25),
.Y(n_182)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_17),
.Y(n_124)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_17),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_59),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.C(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_52),
.C(n_55),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_49),
.B1(n_55),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_33),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_39),
.B(n_118),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_43),
.B(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_43),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_44),
.B(n_124),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_44),
.B(n_246),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_51),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_53),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_72),
.C(n_74),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_55),
.A2(n_74),
.B1(n_79),
.B2(n_324),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_56),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_56),
.B(n_73),
.Y(n_257)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.C(n_81),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_60),
.B(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_71),
.C(n_77),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_61),
.B(n_368),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_62),
.B(n_81),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_64),
.CI(n_65),
.CON(n_62),
.SN(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.C(n_69),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_66),
.B(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_71),
.B(n_77),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_72),
.B(n_349),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_74),
.A2(n_295),
.B1(n_296),
.B2(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_74),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_SL g353 ( 
.A(n_74),
.B(n_295),
.C(n_322),
.Y(n_353)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_372),
.C(n_373),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_363),
.C(n_364),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_341),
.C(n_342),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_317),
.C(n_318),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_285),
.C(n_286),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_251),
.C(n_252),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_216),
.C(n_217),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_186),
.C(n_187),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_165),
.C(n_166),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_147),
.C(n_148),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_125),
.C(n_126),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.C(n_115),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_106),
.B2(n_107),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_108),
.C(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_105),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_103),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.C(n_120),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_124),
.B(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_138),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.C(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_132),
.Y(n_137)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_146),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_151),
.C(n_156),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_154),
.C(n_155),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_164),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_180),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_181),
.C(n_185),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_175),
.C(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_174),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_176),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.CI(n_179),
.CON(n_176),
.SN(n_176)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_178),
.C(n_179),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.CI(n_184),
.CON(n_181),
.SN(n_181)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_202),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_191),
.C(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_198),
.C(n_201),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_193),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.CI(n_196),
.CON(n_193),
.SN(n_193)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_195),
.C(n_196),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_209),
.C(n_214),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_209),
.B1(n_214),
.B2(n_215),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_205),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_207),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_208),
.B(n_241),
.C(n_242),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_209),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_237),
.B2(n_250),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_238),
.C(n_239),
.Y(n_251)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_222),
.C(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_226),
.C(n_229),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_228),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_234),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_249),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_247),
.C(n_249),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_283),
.B2(n_284),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_274),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_274),
.C(n_283),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_263),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_264),
.C(n_265),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_257),
.B(n_259),
.C(n_261),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_273),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_266),
.Y(n_273)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_270),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_269),
.B(n_292),
.C(n_295),
.Y(n_339)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_277),
.C(n_278),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_281),
.C(n_282),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_289),
.C(n_316),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_303),
.B2(n_316),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_291),
.B(n_298),
.C(n_299),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_299),
.Y(n_378)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.CI(n_302),
.CON(n_299),
.SN(n_299)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_301),
.C(n_302),
.Y(n_326)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_315),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_311),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_312),
.A2(n_313),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_338),
.C(n_339),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_340),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_331),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_331),
.C(n_340),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_326),
.C(n_327),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_327),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.CI(n_330),
.CON(n_327),
.SN(n_327)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_329),
.C(n_330),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_334),
.C(n_335),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_337),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_345),
.C(n_355),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_354),
.B2(n_355),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_352),
.C(n_353),
.Y(n_366)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_358),
.C(n_361),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_365),
.A2(n_369),
.B1(n_370),
.B2(n_371),
.Y(n_364)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_365),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_367),
.C(n_371),
.Y(n_372)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_369),
.Y(n_371)
);


endmodule