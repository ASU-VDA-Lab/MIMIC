module real_jpeg_26886_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_0),
.B(n_210),
.Y(n_215)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_0),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_2),
.A2(n_31),
.B1(n_56),
.B2(n_57),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_4),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_4),
.A2(n_35),
.B1(n_37),
.B2(n_53),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_53),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_28),
.B1(n_35),
.B2(n_37),
.Y(n_85)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_8),
.A2(n_35),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_8),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_8),
.B(n_51),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_8),
.A2(n_51),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_92),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_8),
.A2(n_10),
.B(n_35),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_8),
.A2(n_23),
.B(n_40),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_8),
.B(n_71),
.Y(n_205)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_137),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_136),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_110),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_16),
.B(n_110),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_76),
.C(n_87),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_17),
.B(n_76),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_46),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_18),
.B(n_48),
.C(n_64),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_32),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_19),
.B(n_32),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_27),
.B(n_29),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_20),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_21),
.A2(n_25),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_21),
.B(n_79),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_21),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_22),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_25),
.B(n_79),
.Y(n_78)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_27),
.A2(n_80),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_29),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_29),
.B(n_209),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_41),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_33),
.A2(n_85),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_33),
.B(n_192),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_34),
.B(n_44),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_35),
.A2(n_37),
.B1(n_70),
.B2(n_72),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_35),
.A2(n_39),
.B(n_43),
.C(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_38),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_38),
.B(n_42),
.Y(n_191)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_41),
.B(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_42),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_43),
.A2(n_57),
.B(n_174),
.C(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_43),
.B(n_84),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_43),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_44),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_44),
.B(n_182),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_64),
.B2(n_65),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_60),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_49),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_54),
.B(n_55),
.C(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_55),
.Y(n_63)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_54)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_59),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_68),
.B(n_69),
.C(n_71),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_57),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_62),
.B(n_120),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_73),
.B(n_74),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_67),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_67),
.B(n_125),
.Y(n_151)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_71),
.B(n_101),
.Y(n_150)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_72),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_78),
.B(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_81),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_84),
.A2(n_132),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_86),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_87),
.A2(n_88),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_97),
.C(n_102),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_89),
.A2(n_90),
.B1(n_97),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_100),
.B(n_124),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_102),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_108),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_135),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_128),
.B2(n_129),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_150),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_130),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_133),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_130),
.B(n_173),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_167),
.B(n_244),
.C(n_249),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_155),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_139),
.B(n_155),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_152),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_141),
.B(n_142),
.C(n_152),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_148),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_156),
.A2(n_157),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.C(n_165),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_243),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_236),
.B(n_242),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_194),
.B(n_235),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_183),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_171),
.B(n_183),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.C(n_179),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_190),
.C(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_230),
.B(n_234),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_211),
.B(n_229),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_200),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_218),
.B(n_228),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_216),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_222),
.B(n_227),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);


endmodule