module fake_aes_9245_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_12), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_5), .B(n_6), .Y(n_16) );
AND2x6_ASAP7_75t_L g17 ( .A(n_10), .B(n_1), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_1), .Y(n_18) );
AOI22xp5_ASAP7_75t_L g19 ( .A1(n_14), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_15), .B(n_0), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
OAI211xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .B(n_18), .C(n_13), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_21), .Y(n_23) );
AOI222xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_21), .B1(n_17), .B2(n_15), .C1(n_16), .C2(n_2), .Y(n_24) );
OAI21xp33_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_17), .B(n_4), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g26 ( .A(n_24), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_26), .Y(n_27) );
NOR3xp33_ASAP7_75t_SL g28 ( .A(n_25), .B(n_17), .C(n_3), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
AOI322xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_28), .A3(n_15), .B1(n_17), .B2(n_8), .C1(n_9), .C2(n_7), .Y(n_30) );
endmodule