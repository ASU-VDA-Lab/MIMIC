module fake_ariane_322_n_785 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_785);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_785;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_571;
wire n_414;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_484;
wire n_411;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_42),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_35),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_125),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_77),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_83),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_51),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_30),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_43),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_61),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_52),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_91),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_31),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_71),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_6),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_122),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_60),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_126),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_121),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_128),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_56),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_5),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_59),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_64),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_41),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_79),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_24),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_11),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_6),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_92),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_80),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_66),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_11),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_26),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_0),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_85),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_73),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_75),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_3),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_142),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_33),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_100),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_48),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_113),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_156),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_0),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

BUFx8_ASAP7_75t_SL g228 ( 
.A(n_165),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_176),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_176),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_176),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_153),
.B(n_1),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_160),
.B(n_162),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_1),
.Y(n_235)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_171),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_172),
.B(n_2),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

BUFx8_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_187),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_151),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_191),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_190),
.B(n_2),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_186),
.B1(n_167),
.B2(n_177),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_211),
.A2(n_178),
.B1(n_193),
.B2(n_195),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_208),
.A2(n_205),
.B1(n_194),
.B2(n_192),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_208),
.B(n_201),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_210),
.B(n_157),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_158),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_161),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

AO22x2_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_203),
.B1(n_202),
.B2(n_200),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_210),
.A2(n_247),
.B1(n_217),
.B2(n_239),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_199),
.B1(n_198),
.B2(n_196),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_209),
.A2(n_185),
.B1(n_183),
.B2(n_180),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_209),
.Y(n_269)
);

AOI22x1_ASAP7_75t_SL g270 ( 
.A1(n_247),
.A2(n_228),
.B1(n_246),
.B2(n_216),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_234),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_174),
.B1(n_170),
.B2(n_168),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_232),
.A2(n_164),
.B1(n_7),
.B2(n_8),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_4),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g276 ( 
.A(n_235),
.B(n_7),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_216),
.B(n_8),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g280 ( 
.A1(n_246),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_222),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_245),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_237),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_207),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_23),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_237),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_237),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_207),
.B(n_19),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_207),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_245),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_241),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_241),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_241),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_243),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_243),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_252),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_269),
.B(n_238),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_270),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_257),
.B(n_243),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_252),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_255),
.B(n_214),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_243),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_253),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_268),
.B(n_243),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_261),
.B(n_214),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_288),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_262),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_277),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_276),
.B(n_220),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_220),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_283),
.B(n_245),
.Y(n_340)
);

NAND2x1_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_225),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_263),
.B(n_245),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_285),
.B(n_245),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_284),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_284),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_244),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_287),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_296),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_287),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_293),
.B(n_225),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_297),
.B(n_244),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_293),
.Y(n_357)
);

XNOR2x2_ASAP7_75t_L g358 ( 
.A(n_260),
.B(n_297),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_260),
.B(n_226),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_280),
.B(n_244),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_271),
.B(n_226),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_254),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_327),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_328),
.A2(n_240),
.B(n_244),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_34),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_238),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_238),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_215),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_326),
.B(n_238),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_323),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_317),
.B(n_238),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_299),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_314),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_330),
.B(n_244),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_305),
.B(n_244),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_238),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_323),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g389 ( 
.A(n_306),
.B(n_240),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_362),
.A2(n_240),
.B(n_224),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_240),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_315),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_215),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_321),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_324),
.B(n_305),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_306),
.B(n_240),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_215),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_303),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_348),
.A2(n_224),
.B(n_227),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_215),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_347),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_349),
.B(n_351),
.Y(n_405)
);

AND2x2_ASAP7_75t_SL g406 ( 
.A(n_354),
.B(n_215),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_316),
.B(n_218),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_325),
.B(n_218),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_330),
.B(n_227),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_352),
.B(n_218),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_329),
.B(n_218),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_329),
.B(n_218),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_355),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_361),
.B(n_219),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_361),
.B(n_219),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_319),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_343),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_300),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_344),
.B(n_219),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_309),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_308),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_344),
.B(n_219),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_301),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_304),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_307),
.B(n_219),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_364),
.B(n_221),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_354),
.B(n_320),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_405),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_345),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_379),
.B(n_313),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_402),
.B(n_350),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_345),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_356),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_356),
.Y(n_444)
);

OR2x6_ASAP7_75t_L g445 ( 
.A(n_370),
.B(n_358),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_365),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_312),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_369),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_405),
.B(n_302),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_405),
.B(n_370),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_331),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_365),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_402),
.B(n_333),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_405),
.B(n_302),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_365),
.Y(n_460)
);

AO21x2_ASAP7_75t_L g461 ( 
.A1(n_389),
.A2(n_340),
.B(n_231),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_392),
.B(n_310),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_392),
.B(n_221),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_221),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_406),
.B(n_367),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_367),
.B(n_227),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_382),
.B(n_378),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_371),
.Y(n_468)
);

CKINVDCx8_ASAP7_75t_R g469 ( 
.A(n_426),
.Y(n_469)
);

CKINVDCx6p67_ASAP7_75t_R g470 ( 
.A(n_398),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_375),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_406),
.B(n_367),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_424),
.B(n_433),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_426),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_418),
.B(n_221),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_378),
.B(n_36),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_418),
.B(n_231),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_374),
.B(n_221),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_375),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_419),
.B(n_223),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_387),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_381),
.B(n_227),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_419),
.B(n_223),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_374),
.B(n_223),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_401),
.B(n_223),
.Y(n_487)
);

NAND2x1p5_ASAP7_75t_L g488 ( 
.A(n_374),
.B(n_227),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_430),
.B(n_223),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_401),
.B(n_230),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_384),
.B(n_230),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_413),
.Y(n_492)
);

INVx5_ASAP7_75t_SL g493 ( 
.A(n_470),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_444),
.B(n_412),
.Y(n_494)
);

BUFx2_ASAP7_75t_SL g495 ( 
.A(n_469),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

NAND2x1p5_ASAP7_75t_L g497 ( 
.A(n_434),
.B(n_416),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_438),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_438),
.Y(n_499)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_437),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_437),
.Y(n_501)
);

BUFx2_ASAP7_75t_SL g502 ( 
.A(n_474),
.Y(n_502)
);

BUFx12f_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

BUFx4f_ASAP7_75t_SL g504 ( 
.A(n_440),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_438),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g506 ( 
.A(n_443),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_450),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_434),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_447),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_453),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_467),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_439),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_444),
.B(n_384),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_445),
.A2(n_413),
.B1(n_388),
.B2(n_399),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_436),
.Y(n_517)
);

CKINVDCx8_ASAP7_75t_R g518 ( 
.A(n_445),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_447),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_434),
.B(n_416),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_479),
.B(n_376),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_447),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_467),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_441),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_456),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

BUFx5_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_473),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_473),
.Y(n_530)
);

BUFx12f_ASAP7_75t_L g531 ( 
.A(n_458),
.Y(n_531)
);

INVx8_ASAP7_75t_L g532 ( 
.A(n_478),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_446),
.B(n_421),
.Y(n_533)
);

INVx3_ASAP7_75t_SL g534 ( 
.A(n_478),
.Y(n_534)
);

INVx3_ASAP7_75t_SL g535 ( 
.A(n_478),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_451),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_455),
.A2(n_429),
.B1(n_421),
.B2(n_383),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_458),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_473),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_483),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_486),
.Y(n_542)
);

CKINVDCx6p67_ASAP7_75t_R g543 ( 
.A(n_495),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_514),
.Y(n_544)
);

INVx8_ASAP7_75t_L g545 ( 
.A(n_532),
.Y(n_545)
);

BUFx12f_ASAP7_75t_L g546 ( 
.A(n_503),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_507),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_514),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_496),
.B(n_457),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_526),
.B(n_471),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_508),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_524),
.A2(n_435),
.B1(n_442),
.B2(n_492),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_509),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_494),
.A2(n_455),
.B(n_442),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_524),
.A2(n_435),
.B1(n_484),
.B2(n_399),
.Y(n_555)
);

CKINVDCx11_ASAP7_75t_R g556 ( 
.A(n_503),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_516),
.A2(n_476),
.B1(n_472),
.B2(n_465),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_531),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_498),
.Y(n_559)
);

BUFx12f_ASAP7_75t_L g560 ( 
.A(n_500),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_518),
.A2(n_472),
.B1(n_465),
.B2(n_459),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_516),
.A2(n_468),
.B1(n_393),
.B2(n_449),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_493),
.Y(n_563)
);

BUFx4f_ASAP7_75t_SL g564 ( 
.A(n_531),
.Y(n_564)
);

INVx6_ASAP7_75t_L g565 ( 
.A(n_532),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_515),
.A2(n_430),
.B1(n_457),
.B2(n_460),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_502),
.Y(n_567)
);

BUFx12f_ASAP7_75t_L g568 ( 
.A(n_500),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_525),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_513),
.B(n_463),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_518),
.A2(n_459),
.B1(n_454),
.B2(n_449),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_512),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_501),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_504),
.A2(n_460),
.B1(n_454),
.B2(n_422),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_506),
.A2(n_393),
.B1(n_491),
.B2(n_422),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_506),
.A2(n_428),
.B1(n_376),
.B2(n_420),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_527),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_523),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_521),
.A2(n_428),
.B1(n_420),
.B2(n_403),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_505),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_504),
.A2(n_403),
.B1(n_389),
.B2(n_429),
.Y(n_582)
);

CKINVDCx11_ASAP7_75t_R g583 ( 
.A(n_517),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_525),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_557),
.A2(n_528),
.B1(n_538),
.B2(n_523),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_555),
.A2(n_538),
.B1(n_539),
.B2(n_529),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_567),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_576),
.A2(n_528),
.B1(n_536),
.B2(n_372),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_576),
.A2(n_528),
.B1(n_536),
.B2(n_407),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_550),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_555),
.A2(n_528),
.B1(n_407),
.B2(n_394),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_547),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_529),
.Y(n_593)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_552),
.B(n_539),
.C(n_411),
.Y(n_594)
);

BUFx5_ASAP7_75t_L g595 ( 
.A(n_581),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_579),
.A2(n_537),
.B1(n_535),
.B2(n_534),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_561),
.A2(n_528),
.B1(n_407),
.B2(n_394),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_571),
.A2(n_530),
.B(n_533),
.Y(n_598)
);

OAI21xp33_ASAP7_75t_L g599 ( 
.A1(n_554),
.A2(n_415),
.B(n_414),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_552),
.A2(n_528),
.B1(n_407),
.B2(n_394),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_570),
.B(n_578),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_575),
.A2(n_407),
.B1(n_394),
.B2(n_373),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_579),
.A2(n_535),
.B1(n_534),
.B2(n_493),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_575),
.A2(n_394),
.B1(n_373),
.B2(n_421),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_553),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_L g606 ( 
.A1(n_564),
.A2(n_532),
.B1(n_496),
.B2(n_542),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_562),
.A2(n_429),
.B1(n_542),
.B2(n_482),
.Y(n_607)
);

INVx3_ASAP7_75t_SL g608 ( 
.A(n_543),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_572),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_562),
.A2(n_482),
.B1(n_493),
.B2(n_396),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_583),
.A2(n_425),
.B1(n_477),
.B2(n_464),
.Y(n_611)
);

AND2x2_ASAP7_75t_SL g612 ( 
.A(n_577),
.B(n_496),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_560),
.A2(n_425),
.B1(n_464),
.B2(n_522),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_544),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_573),
.B(n_489),
.C(n_505),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_564),
.A2(n_560),
.B1(n_546),
.B2(n_568),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_580),
.B(n_498),
.Y(n_617)
);

INVx3_ASAP7_75t_SL g618 ( 
.A(n_563),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_566),
.A2(n_540),
.B1(n_533),
.B2(n_486),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_574),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_584),
.A2(n_425),
.B1(n_522),
.B2(n_499),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_546),
.A2(n_425),
.B1(n_511),
.B2(n_499),
.Y(n_622)
);

OAI21xp33_ASAP7_75t_L g623 ( 
.A1(n_582),
.A2(n_431),
.B(n_432),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_578),
.B(n_511),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_556),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_544),
.Y(n_626)
);

OAI21xp33_ASAP7_75t_L g627 ( 
.A1(n_559),
.A2(n_423),
.B(n_427),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_558),
.A2(n_510),
.B1(n_540),
.B2(n_519),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_559),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_548),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_548),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_558),
.A2(n_486),
.B1(n_510),
.B2(n_520),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_569),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_565),
.A2(n_497),
.B1(n_520),
.B2(n_409),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_565),
.A2(n_497),
.B1(n_505),
.B2(n_519),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_592),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_601),
.B(n_581),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_620),
.A2(n_565),
.B1(n_549),
.B2(n_545),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_594),
.A2(n_569),
.B1(n_545),
.B2(n_397),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_620),
.A2(n_596),
.B1(n_586),
.B2(n_603),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_605),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_588),
.A2(n_425),
.B1(n_461),
.B2(n_408),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_610),
.A2(n_461),
.B1(n_490),
.B2(n_487),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_615),
.A2(n_490),
.B1(n_487),
.B2(n_466),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_585),
.A2(n_545),
.B1(n_485),
.B2(n_475),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_590),
.B(n_505),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_602),
.A2(n_605),
.B1(n_604),
.B2(n_609),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_614),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_617),
.B(n_549),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_616),
.A2(n_410),
.B1(n_404),
.B2(n_377),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_626),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_597),
.A2(n_410),
.B1(n_404),
.B2(n_377),
.Y(n_652)
);

OAI21xp33_ASAP7_75t_SL g653 ( 
.A1(n_612),
.A2(n_485),
.B(n_480),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_SL g654 ( 
.A(n_608),
.B(n_385),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_598),
.A2(n_480),
.B1(n_475),
.B2(n_366),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_611),
.A2(n_400),
.B1(n_391),
.B2(n_390),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_589),
.A2(n_386),
.B1(n_385),
.B2(n_231),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_591),
.A2(n_386),
.B1(n_385),
.B2(n_409),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_629),
.B(n_37),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_593),
.B(n_230),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_SL g661 ( 
.A1(n_635),
.A2(n_231),
.B1(n_230),
.B2(n_488),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_628),
.A2(n_386),
.B1(n_409),
.B2(n_488),
.Y(n_662)
);

NAND4xp25_ASAP7_75t_L g663 ( 
.A(n_587),
.B(n_599),
.C(n_607),
.D(n_627),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_600),
.A2(n_229),
.B1(n_224),
.B2(n_40),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_630),
.A2(n_229),
.B1(n_224),
.B2(n_44),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_631),
.A2(n_229),
.B1(n_224),
.B2(n_45),
.Y(n_666)
);

OAI222xp33_ASAP7_75t_L g667 ( 
.A1(n_633),
.A2(n_229),
.B1(n_224),
.B2(n_46),
.C1(n_47),
.C2(n_49),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_619),
.A2(n_229),
.B1(n_39),
.B2(n_50),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_613),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_632),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_624),
.B(n_62),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_625),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_618),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_634),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_606),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_L g676 ( 
.A(n_663),
.B(n_623),
.C(n_608),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_641),
.B(n_618),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_636),
.B(n_595),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_640),
.A2(n_622),
.B(n_621),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_673),
.A2(n_595),
.B1(n_86),
.B2(n_87),
.Y(n_680)
);

OAI31xp33_ASAP7_75t_SL g681 ( 
.A1(n_638),
.A2(n_595),
.A3(n_88),
.B(n_89),
.Y(n_681)
);

OAI211xp5_ASAP7_75t_SL g682 ( 
.A1(n_660),
.A2(n_595),
.B(n_93),
.C(n_94),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_639),
.B(n_595),
.C(n_95),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_646),
.B(n_595),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_649),
.B(n_149),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_637),
.B(n_84),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_659),
.B(n_148),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_639),
.B(n_96),
.C(n_97),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_647),
.B(n_98),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_651),
.B(n_101),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_673),
.B(n_672),
.C(n_653),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_647),
.B(n_102),
.Y(n_692)
);

OAI21xp33_ASAP7_75t_L g693 ( 
.A1(n_672),
.A2(n_104),
.B(n_105),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_671),
.B(n_147),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_668),
.B(n_106),
.C(n_107),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_664),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_648),
.B(n_112),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_664),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_698)
);

OA211x2_ASAP7_75t_L g699 ( 
.A1(n_645),
.A2(n_119),
.B(n_120),
.C(n_123),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_655),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_643),
.B(n_124),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_675),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_702)
);

NAND3xp33_ASAP7_75t_L g703 ( 
.A(n_674),
.B(n_132),
.C(n_133),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_678),
.B(n_670),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_677),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_678),
.B(n_657),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_691),
.A2(n_654),
.B1(n_661),
.B2(n_650),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_684),
.B(n_657),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_700),
.B(n_642),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_700),
.Y(n_710)
);

OA211x2_ASAP7_75t_L g711 ( 
.A1(n_693),
.A2(n_683),
.B(n_679),
.C(n_692),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_690),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_686),
.B(n_662),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_676),
.B(n_667),
.C(n_652),
.Y(n_714)
);

NAND4xp75_ASAP7_75t_L g715 ( 
.A(n_699),
.B(n_669),
.C(n_666),
.D(n_665),
.Y(n_715)
);

OR3x1_ASAP7_75t_L g716 ( 
.A(n_682),
.B(n_644),
.C(n_658),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_686),
.B(n_656),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_687),
.B(n_135),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_689),
.B(n_137),
.C(n_139),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_685),
.B(n_681),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_690),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_708),
.B(n_697),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_710),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_721),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_705),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_708),
.B(n_697),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_706),
.B(n_680),
.Y(n_727)
);

INVx8_ASAP7_75t_L g728 ( 
.A(n_718),
.Y(n_728)
);

XNOR2x1_ASAP7_75t_L g729 ( 
.A(n_711),
.B(n_701),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_718),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_712),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_721),
.Y(n_732)
);

OAI31xp33_ASAP7_75t_L g733 ( 
.A1(n_720),
.A2(n_701),
.A3(n_688),
.B(n_695),
.Y(n_733)
);

XOR2x2_ASAP7_75t_L g734 ( 
.A(n_729),
.B(n_730),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_729),
.Y(n_735)
);

XOR2x2_ASAP7_75t_L g736 ( 
.A(n_722),
.B(n_715),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_725),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_727),
.B(n_717),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_734),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_736),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_737),
.Y(n_741)
);

INVx3_ASAP7_75t_SL g742 ( 
.A(n_735),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_738),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_741),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_743),
.Y(n_745)
);

OA22x2_ASAP7_75t_L g746 ( 
.A1(n_739),
.A2(n_738),
.B1(n_727),
.B2(n_726),
.Y(n_746)
);

OAI22x1_ASAP7_75t_L g747 ( 
.A1(n_744),
.A2(n_742),
.B1(n_740),
.B2(n_743),
.Y(n_747)
);

OAI322xp33_ASAP7_75t_L g748 ( 
.A1(n_746),
.A2(n_742),
.A3(n_731),
.B1(n_707),
.B2(n_741),
.C1(n_723),
.C2(n_733),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_747),
.A2(n_716),
.B1(n_745),
.B2(n_714),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_748),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_747),
.A2(n_716),
.B1(n_745),
.B2(n_709),
.Y(n_751)
);

NOR4xp25_ASAP7_75t_L g752 ( 
.A(n_750),
.B(n_719),
.C(n_696),
.D(n_698),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_749),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_751),
.A2(n_709),
.B1(n_728),
.B2(n_704),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_750),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_750),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_750),
.A2(n_728),
.B1(n_704),
.B2(n_694),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_751),
.B(n_728),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_753),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_755),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_756),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_752),
.B(n_757),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_758),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_754),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_761),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_762),
.A2(n_713),
.B1(n_704),
.B2(n_702),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_760),
.Y(n_767)
);

NOR2x1_ASAP7_75t_L g768 ( 
.A(n_760),
.B(n_703),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_765),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_767),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_768),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_766),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_767),
.Y(n_773)
);

INVxp67_ASAP7_75t_SL g774 ( 
.A(n_771),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_769),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_770),
.Y(n_776)
);

NAND4xp75_ASAP7_75t_L g777 ( 
.A(n_773),
.B(n_759),
.C(n_763),
.D(n_764),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_774),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_777),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_778),
.A2(n_776),
.B1(n_775),
.B2(n_772),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_780),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_781),
.A2(n_779),
.B(n_698),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_782),
.Y(n_783)
);

AOI221xp5_ASAP7_75t_L g784 ( 
.A1(n_783),
.A2(n_732),
.B1(n_724),
.B2(n_713),
.C(n_706),
.Y(n_784)
);

AOI211xp5_ASAP7_75t_L g785 ( 
.A1(n_784),
.A2(n_724),
.B(n_141),
.C(n_143),
.Y(n_785)
);


endmodule